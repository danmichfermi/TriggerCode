LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY code_450 IS
   PORT(
      --*************************************************
      -- V1495 Front Panel Ports (PORT A,B,C,G)
      --*************************************************
      A_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In A (32 x LVDS/ECL)
      B_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In B (32 x LVDS/ECL)
      D_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In D (32 x LVDS/ECL)
      E_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In E (32 x LVDS/ECL)
      F_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- OUT F (32 x LVDS/ECL)
      C_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- Out C (32 x LVDS)
      c1            : IN STD_LOGIC                            -- the PLL1 output
   );
END code_450 ;
ARCHITECTURE rtl OF code_450 IS
	signal A     : std_logic_vector(31 downto 0);
	signal B     : std_logic_vector(31 downto 0);
	signal C     : std_logic_vector(31 downto 0);
	signal D     : std_logic_vector(31 downto 0);
	signal E     : std_logic_vector(31 downto 0);
	signal F     : std_logic_vector(31 downto 0);
	signal G     : std_logic_vector(1 downto 0);
	signal output	: std_logic_vector(31 downto 0);
	signal cut : std_logic_vector(3 downto 0);
	signal results : std_logic_vector(3 downto 0);

component Adder_type
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
end component;
component  ADDM4K3S8RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S9RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S12RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S13RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S10RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S11RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S14RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S15RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S2RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S3RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S4RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S5RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S6RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S7RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S0RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S1RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

        signal cVar1S0S0P069P019P067P064: std_logic_vector(   0 downto 0);
        signal cVar1S1S0P069P019P067P064: std_logic_vector(   0 downto 0);
        signal cVar1S2S0P069P019P067P064: std_logic_vector(   0 downto 0);
        signal cVar1S3S0P069P019P067N064: std_logic_vector(   0 downto 0);
        signal cVar1S4S0P069P019P067N064: std_logic_vector(   0 downto 0);
        signal cVar1S5S0P069P019P067N064: std_logic_vector(   0 downto 0);
        signal cVar1S6S0P069P019P067N064: std_logic_vector(   0 downto 0);
        signal cVar1S7S0P069P019N067P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S0P069P019N067P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S0P069N019P036P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S0P069N019P036P017: std_logic_vector(   0 downto 0);
        signal cVar1S11S0P069N019P036P017: std_logic_vector(   0 downto 0);
        signal cVar1S12S0P069N019P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S13S0P069N019P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S14S0P069N019P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S15S0P069N019N036P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S0P069N019N036P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S0P069N019N036N018: std_logic_vector(   0 downto 0);
        signal cVar1S18S0N069P063P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S0N069P063P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S20S0N069P063P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S21S0N069P063P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S22S0N069P063P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S23S0N069P063P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S24S0N069P063P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S25S0N069P063P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S26S0N069P063N065P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S0N069P063N065P061: std_logic_vector(   0 downto 0);
        signal cVar1S28S0N069N063P061P059: std_logic_vector(   0 downto 0);
        signal cVar1S29S0N069N063P061P059: std_logic_vector(   0 downto 0);
        signal cVar1S30S0N069N063P061P059: std_logic_vector(   0 downto 0);
        signal cVar1S31S0N069N063P061P059: std_logic_vector(   0 downto 0);
        signal cVar1S32S0N069N063N061P055: std_logic_vector(   0 downto 0);
        signal cVar1S33S0N069N063N061P055: std_logic_vector(   0 downto 0);
        signal cVar1S34S0N069N063N061P055: std_logic_vector(   0 downto 0);
        signal cVar1S35S0N069N063N061P055: std_logic_vector(   0 downto 0);
        signal cVar1S36S0N069N063N061N055: std_logic_vector(   0 downto 0);
        signal cVar1S37S0N069N063N061N055: std_logic_vector(   0 downto 0);
        signal cVar1S0S1P052P050P010P068: std_logic_vector(   0 downto 0);
        signal cVar1S1S1P052P050P010P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S1P052P050P010P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S1P052P050P010P068: std_logic_vector(   0 downto 0);
        signal cVar1S4S1P052P050N010P069: std_logic_vector(   0 downto 0);
        signal cVar1S5S1P052P050N010P069: std_logic_vector(   0 downto 0);
        signal cVar1S6S1P052P050N010N069: std_logic_vector(   0 downto 0);
        signal cVar1S7S1P052P050N010N069: std_logic_vector(   0 downto 0);
        signal cVar1S8S1P052N050P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S1P052N050N029P028: std_logic_vector(   0 downto 0);
        signal cVar1S10S1P052N050N029N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S1N052P056P031P063: std_logic_vector(   0 downto 0);
        signal cVar1S12S1N052P056P031P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S1N052P056P031N063psss: std_logic_vector(   0 downto 0);
        signal cVar1S14S1N052P056N031P029: std_logic_vector(   0 downto 0);
        signal cVar1S15S1N052P056N031N029: std_logic_vector(   0 downto 0);
        signal cVar1S16S1N052P056N031N029: std_logic_vector(   0 downto 0);
        signal cVar1S17S1N052P056N031N029: std_logic_vector(   0 downto 0);
        signal cVar1S18S1N052P056N031N029: std_logic_vector(   0 downto 0);
        signal cVar1S19S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S21S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S22S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S23S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S25S1N052N056P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S26S1N052N056N060P046: std_logic_vector(   0 downto 0);
        signal cVar1S27S1N052N056N060P046: std_logic_vector(   0 downto 0);
        signal cVar1S28S1N052N056N060P046: std_logic_vector(   0 downto 0);
        signal cVar1S29S1N052N056N060N046: std_logic_vector(   0 downto 0);
        signal cVar1S30S1N052N056N060N046: std_logic_vector(   0 downto 0);
        signal cVar1S31S1N052N056N060N046: std_logic_vector(   0 downto 0);
        signal cVar1S0S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S1S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S2S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S3S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S4S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S5S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S6S2P068P067P066P035: std_logic_vector(   0 downto 0);
        signal cVar1S7S2P068P067N066P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S2P068P067N066P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S2P068P067N066N063: std_logic_vector(   0 downto 0);
        signal cVar1S10S2P068P067N066N063: std_logic_vector(   0 downto 0);
        signal cVar1S11S2P068P067P035P016: std_logic_vector(   0 downto 0);
        signal cVar1S12S2P068P067P035P016: std_logic_vector(   0 downto 0);
        signal cVar1S13S2P068P067P035P016: std_logic_vector(   0 downto 0);
        signal cVar1S14S2P068P067P035N016: std_logic_vector(   0 downto 0);
        signal cVar1S15S2P068P067P035N016: std_logic_vector(   0 downto 0);
        signal cVar1S16S2P068P067P035N016: std_logic_vector(   0 downto 0);
        signal cVar1S17S2P068P067P035P031nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S2P068P067P035N031: std_logic_vector(   0 downto 0);
        signal cVar1S19S2N068P063P062P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S2N068P063P062P065: std_logic_vector(   0 downto 0);
        signal cVar1S21S2N068P063P062P065: std_logic_vector(   0 downto 0);
        signal cVar1S22S2N068P063P062N065: std_logic_vector(   0 downto 0);
        signal cVar1S23S2N068P063P062N065: std_logic_vector(   0 downto 0);
        signal cVar1S24S2N068P063P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S25S2N068P063P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S26S2N068P063P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S27S2N068P063P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S28S2N068P063P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S29S2N068N063P051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S2N068N063P051N028: std_logic_vector(   0 downto 0);
        signal cVar1S31S2N068N063P051N028: std_logic_vector(   0 downto 0);
        signal cVar1S32S2N068N063P051N028: std_logic_vector(   0 downto 0);
        signal cVar1S33S2N068N063N051P067: std_logic_vector(   0 downto 0);
        signal cVar1S34S2N068N063N051P067: std_logic_vector(   0 downto 0);
        signal cVar1S35S2N068N063N051P067: std_logic_vector(   0 downto 0);
        signal cVar1S36S2N068N063N051P067: std_logic_vector(   0 downto 0);
        signal cVar1S37S2N068N063N051N067: std_logic_vector(   0 downto 0);
        signal cVar1S38S2N068N063N051N067: std_logic_vector(   0 downto 0);
        signal cVar1S39S2N068N063N051N067: std_logic_vector(   0 downto 0);
        signal cVar1S40S2N068N063N051N067: std_logic_vector(   0 downto 0);
        signal cVar1S0S3P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S3P043N022P007P015: std_logic_vector(   0 downto 0);
        signal cVar1S2S3P043N022P007P015: std_logic_vector(   0 downto 0);
        signal cVar1S3S3P043N022P007P015psss: std_logic_vector(   0 downto 0);
        signal cVar1S4S3P043N022N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S5S3P043N022N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S6S3P043N022N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S7S3N043P067P068P060: std_logic_vector(   0 downto 0);
        signal cVar1S8S3N043P067P068P060: std_logic_vector(   0 downto 0);
        signal cVar1S9S3N043P067P068P060: std_logic_vector(   0 downto 0);
        signal cVar1S10S3N043P067P068P060: std_logic_vector(   0 downto 0);
        signal cVar1S11S3N043P067P068P016: std_logic_vector(   0 downto 0);
        signal cVar1S12S3N043P067P068P016: std_logic_vector(   0 downto 0);
        signal cVar1S13S3N043P067P068N016: std_logic_vector(   0 downto 0);
        signal cVar1S14S3N043P067P068N016: std_logic_vector(   0 downto 0);
        signal cVar1S15S3N043P067P068N016: std_logic_vector(   0 downto 0);
        signal cVar1S16S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S17S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S18S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S19S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S20S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S21S3N043N067P034P062: std_logic_vector(   0 downto 0);
        signal cVar1S22S3N043N067N034P051: std_logic_vector(   0 downto 0);
        signal cVar1S23S3N043N067N034P051: std_logic_vector(   0 downto 0);
        signal cVar1S24S3N043N067N034P051: std_logic_vector(   0 downto 0);
        signal cVar1S25S3N043N067N034N051: std_logic_vector(   0 downto 0);
        signal cVar1S26S3N043N067N034N051: std_logic_vector(   0 downto 0);
        signal cVar1S27S3N043N067N034N051: std_logic_vector(   0 downto 0);
        signal cVar1S0S4P044P023P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S4P044P023N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S4P044P023N006N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S4P044N023P025P018: std_logic_vector(   0 downto 0);
        signal cVar1S4S4P044N023P025P018: std_logic_vector(   0 downto 0);
        signal cVar1S5S4P044N023P025P018psss: std_logic_vector(   0 downto 0);
        signal cVar1S6S4P044N023N025P022: std_logic_vector(   0 downto 0);
        signal cVar1S7S4P044N023N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S8S4P044N023N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S9S4N044P037P008P067: std_logic_vector(   0 downto 0);
        signal cVar1S10S4N044P037P008P067: std_logic_vector(   0 downto 0);
        signal cVar1S11S4N044P037P008P067: std_logic_vector(   0 downto 0);
        signal cVar1S12S4N044P037P008P067: std_logic_vector(   0 downto 0);
        signal cVar1S13S4N044P037P008P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S4N044P037P008P050: std_logic_vector(   0 downto 0);
        signal cVar1S15S4N044P037P008N050: std_logic_vector(   0 downto 0);
        signal cVar1S16S4N044P037P008N050: std_logic_vector(   0 downto 0);
        signal cVar1S17S4N044N037P031P066: std_logic_vector(   0 downto 0);
        signal cVar1S18S4N044N037P031P066: std_logic_vector(   0 downto 0);
        signal cVar1S19S4N044N037P031P066: std_logic_vector(   0 downto 0);
        signal cVar1S20S4N044N037P031P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S4N044N037P031P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S4N044N037N031P036: std_logic_vector(   0 downto 0);
        signal cVar1S23S4N044N037N031P036: std_logic_vector(   0 downto 0);
        signal cVar1S24S4N044N037N031P036: std_logic_vector(   0 downto 0);
        signal cVar1S25S4N044N037N031P036: std_logic_vector(   0 downto 0);
        signal cVar1S26S4N044N037N031N036: std_logic_vector(   0 downto 0);
        signal cVar1S27S4N044N037N031N036: std_logic_vector(   0 downto 0);
        signal cVar1S28S4N044N037N031N036: std_logic_vector(   0 downto 0);
        signal cVar1S0S5P027P048P052P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S5P027P048P052N050: std_logic_vector(   0 downto 0);
        signal cVar1S2S5P027P048P052N050: std_logic_vector(   0 downto 0);
        signal cVar1S3S5P027P048P052N050: std_logic_vector(   0 downto 0);
        signal cVar1S4S5P027P048P052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S5P027N048P050P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S5P027N048P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S7S5P027N048P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S8S5P027N048P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S9S5P027N048N050P049: std_logic_vector(   0 downto 0);
        signal cVar1S10S5P027N048N050N049: std_logic_vector(   0 downto 0);
        signal cVar1S11S5P027N048N050N049: std_logic_vector(   0 downto 0);
        signal cVar1S12S5P027N048N050N049: std_logic_vector(   0 downto 0);
        signal cVar1S13S5N027P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S5N027P043N022P007: std_logic_vector(   0 downto 0);
        signal cVar1S15S5N027P043N022N007: std_logic_vector(   0 downto 0);
        signal cVar1S16S5N027P043N022N007: std_logic_vector(   0 downto 0);
        signal cVar1S17S5N027P043N022N007: std_logic_vector(   0 downto 0);
        signal cVar1S18S5N027P043N022N007: std_logic_vector(   0 downto 0);
        signal cVar1S19S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S22S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S23S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S24S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S25S5N027N043P036P015: std_logic_vector(   0 downto 0);
        signal cVar1S26S5N027N043N036P068: std_logic_vector(   0 downto 0);
        signal cVar1S27S5N027N043N036P068: std_logic_vector(   0 downto 0);
        signal cVar1S28S5N027N043N036P068: std_logic_vector(   0 downto 0);
        signal cVar1S29S5N027N043N036N068: std_logic_vector(   0 downto 0);
        signal cVar1S30S5N027N043N036N068: std_logic_vector(   0 downto 0);
        signal cVar1S31S5N027N043N036N068: std_logic_vector(   0 downto 0);
        signal cVar1S32S5N027N043N036N068: std_logic_vector(   0 downto 0);
        signal cVar1S0S6P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S6P040N021P023P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S6P040N021P023N018: std_logic_vector(   0 downto 0);
        signal cVar1S3S6P040N021N023P020: std_logic_vector(   0 downto 0);
        signal cVar1S4S6P040N021N023P020: std_logic_vector(   0 downto 0);
        signal cVar1S5S6P040N021N023N020: std_logic_vector(   0 downto 0);
        signal cVar1S6S6P040N021N023N020: std_logic_vector(   0 downto 0);
        signal cVar1S7S6N040P025P046P016: std_logic_vector(   0 downto 0);
        signal cVar1S8S6N040P025P046P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S6N040P025N046P044nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S6N040P025N046N044: std_logic_vector(   0 downto 0);
        signal cVar1S11S6N040P025N046N044: std_logic_vector(   0 downto 0);
        signal cVar1S12S6N040P025N046N044: std_logic_vector(   0 downto 0);
        signal cVar1S13S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S14S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S15S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S6N040N025P056P055: std_logic_vector(   0 downto 0);
        signal cVar1S20S6N040N025N056P060: std_logic_vector(   0 downto 0);
        signal cVar1S21S6N040N025N056P060: std_logic_vector(   0 downto 0);
        signal cVar1S22S6N040N025N056P060: std_logic_vector(   0 downto 0);
        signal cVar1S23S6N040N025N056N060: std_logic_vector(   0 downto 0);
        signal cVar1S24S6N040N025N056N060: std_logic_vector(   0 downto 0);
        signal cVar1S25S6N040N025N056N060: std_logic_vector(   0 downto 0);
        signal cVar1S26S6N040N025N056N060: std_logic_vector(   0 downto 0);
        signal cVar1S0S7P066P028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S7P066P028N055P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S7P066P028N055N053: std_logic_vector(   0 downto 0);
        signal cVar1S3S7P066P028N055N053: std_logic_vector(   0 downto 0);
        signal cVar1S4S7P066P028N055N053: std_logic_vector(   0 downto 0);
        signal cVar1S5S7P066P028N055N053: std_logic_vector(   0 downto 0);
        signal cVar1S6S7P066N028P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S7P066N028P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S8S7P066N028P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S9S7P066N028P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S10S7P066N028P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S11S7P066N028N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S12S7P066N028N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S13S7P066N028N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S14S7P066N028N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S15S7P066N028N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S16S7P066N028N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S17S7P066P065P003P067: std_logic_vector(   0 downto 0);
        signal cVar1S18S7P066P065P003P067: std_logic_vector(   0 downto 0);
        signal cVar1S19S7P066P065P003P067: std_logic_vector(   0 downto 0);
        signal cVar1S20S7P066P065P003P067: std_logic_vector(   0 downto 0);
        signal cVar1S21S7P066P065P003P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S7P066P065P003N041: std_logic_vector(   0 downto 0);
        signal cVar1S23S7P066P065P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S24S7P066P065P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S25S7P066P065P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S26S7P066P065P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S27S7P066P065P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S28S7P066P065P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S29S7P066P065P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S0S8P043P045P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S8P043P045N064P031: std_logic_vector(   0 downto 0);
        signal cVar1S2S8P043P045N064P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S8P043P045N064P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S8P043N045P005P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S8P043N045P005N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S8P043N045N005P022: std_logic_vector(   0 downto 0);
        signal cVar1S7S8P043N045N005N022: std_logic_vector(   0 downto 0);
        signal cVar1S8S8P043N045N005N022: std_logic_vector(   0 downto 0);
        signal cVar1S9S8N043P003P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S8N043P003P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S11S8N043P003P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S12S8N043P003P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S13S8N043P003N040P026: std_logic_vector(   0 downto 0);
        signal cVar1S14S8N043P003N040P026: std_logic_vector(   0 downto 0);
        signal cVar1S15S8N043P003N040P026: std_logic_vector(   0 downto 0);
        signal cVar1S16S8N043P003N040N026: std_logic_vector(   0 downto 0);
        signal cVar1S17S8N043P003N040N026: std_logic_vector(   0 downto 0);
        signal cVar1S18S8N043P003N040N026: std_logic_vector(   0 downto 0);
        signal cVar1S19S8N043P003P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S8N043P003P039N020: std_logic_vector(   0 downto 0);
        signal cVar1S21S8N043P003P039N020: std_logic_vector(   0 downto 0);
        signal cVar1S22S8N043P003N039P036: std_logic_vector(   0 downto 0);
        signal cVar1S23S8N043P003N039N036: std_logic_vector(   0 downto 0);
        signal cVar1S24S8N043P003N039N036: std_logic_vector(   0 downto 0);
        signal cVar1S0S9P032P015P062P059: std_logic_vector(   0 downto 0);
        signal cVar1S1S9P032P015P062P059: std_logic_vector(   0 downto 0);
        signal cVar1S2S9P032P015P062P059: std_logic_vector(   0 downto 0);
        signal cVar1S3S9P032P015P062P059: std_logic_vector(   0 downto 0);
        signal cVar1S4S9P032P015P062N059: std_logic_vector(   0 downto 0);
        signal cVar1S5S9P032P015P062N059: std_logic_vector(   0 downto 0);
        signal cVar1S6S9P032P015P062N059: std_logic_vector(   0 downto 0);
        signal cVar1S7S9P032P015P062N059: std_logic_vector(   0 downto 0);
        signal cVar1S8S9P032P015P062P055: std_logic_vector(   0 downto 0);
        signal cVar1S9S9P032P015P062P055: std_logic_vector(   0 downto 0);
        signal cVar1S10S9P032P015P063P059nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S9P032P015P063N059: std_logic_vector(   0 downto 0);
        signal cVar1S12S9P032P015N063P068: std_logic_vector(   0 downto 0);
        signal cVar1S13S9P032P015N063P068: std_logic_vector(   0 downto 0);
        signal cVar1S14S9P032P015N063N068: std_logic_vector(   0 downto 0);
        signal cVar1S15S9P032P015N063N068: std_logic_vector(   0 downto 0);
        signal cVar1S16S9P032P015N063N068: std_logic_vector(   0 downto 0);
        signal cVar1S17S9P032P015N063N068: std_logic_vector(   0 downto 0);
        signal cVar1S18S9N032P043P045P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S9N032P043P045N062: std_logic_vector(   0 downto 0);
        signal cVar1S20S9N032P043P045N062: std_logic_vector(   0 downto 0);
        signal cVar1S21S9N032P043N045P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S9N032P043N045N005: std_logic_vector(   0 downto 0);
        signal cVar1S23S9N032P043N045N005: std_logic_vector(   0 downto 0);
        signal cVar1S24S9N032P043N045N005: std_logic_vector(   0 downto 0);
        signal cVar1S25S9N032N043P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S9N032N043P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S27S9N032N043P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S28S9N032N043P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S29S9N032N043N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S30S9N032N043N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S31S9N032N043N044P040: std_logic_vector(   0 downto 0);
        signal cVar1S32S9N032N043N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S33S9N032N043N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S34S9N032N043N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S35S9N032N043N044N040: std_logic_vector(   0 downto 0);
        signal cVar1S0S10P032P015P062P061: std_logic_vector(   0 downto 0);
        signal cVar1S1S10P032P015P062P061: std_logic_vector(   0 downto 0);
        signal cVar1S2S10P032P015P062P061: std_logic_vector(   0 downto 0);
        signal cVar1S3S10P032P015P062P061: std_logic_vector(   0 downto 0);
        signal cVar1S4S10P032P015P062N061: std_logic_vector(   0 downto 0);
        signal cVar1S5S10P032P015P062N061: std_logic_vector(   0 downto 0);
        signal cVar1S6S10P032P015P062P055: std_logic_vector(   0 downto 0);
        signal cVar1S7S10P032P015P062P055: std_logic_vector(   0 downto 0);
        signal cVar1S8S10P032P015P063P057: std_logic_vector(   0 downto 0);
        signal cVar1S9S10P032P015P063P057: std_logic_vector(   0 downto 0);
        signal cVar1S10S10P032P015P063P057: std_logic_vector(   0 downto 0);
        signal cVar1S11S10P032P015N063P018: std_logic_vector(   0 downto 0);
        signal cVar1S12S10P032P015N063P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S10P032P015N063N018: std_logic_vector(   0 downto 0);
        signal cVar1S14S10P032P015N063N018: std_logic_vector(   0 downto 0);
        signal cVar1S15S10P032P015N063N018: std_logic_vector(   0 downto 0);
        signal cVar1S16S10N032P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S18S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S19S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S20S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S21S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S22S10N032P040N021P010: std_logic_vector(   0 downto 0);
        signal cVar1S23S10N032N040P043P062: std_logic_vector(   0 downto 0);
        signal cVar1S24S10N032N040P043P062: std_logic_vector(   0 downto 0);
        signal cVar1S25S10N032N040P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S26S10N032N040P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S27S10N032N040P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S28S10N032N040P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S29S10N032N040N043P033: std_logic_vector(   0 downto 0);
        signal cVar1S30S10N032N040N043P033: std_logic_vector(   0 downto 0);
        signal cVar1S31S10N032N040N043P033: std_logic_vector(   0 downto 0);
        signal cVar1S32S10N032N040N043N033: std_logic_vector(   0 downto 0);
        signal cVar1S33S10N032N040N043N033: std_logic_vector(   0 downto 0);
        signal cVar1S34S10N032N040N043N033: std_logic_vector(   0 downto 0);
        signal cVar1S35S10N032N040N043N033: std_logic_vector(   0 downto 0);
        signal cVar1S0S11P027P008P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S11P027P008N046P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S11P027P008N046N050: std_logic_vector(   0 downto 0);
        signal cVar1S3S11P027N008P050P052: std_logic_vector(   0 downto 0);
        signal cVar1S4S11P027N008P050P052: std_logic_vector(   0 downto 0);
        signal cVar1S5S11P027N008P050P052: std_logic_vector(   0 downto 0);
        signal cVar1S6S11P027N008N050P018: std_logic_vector(   0 downto 0);
        signal cVar1S7S11P027N008N050P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S11P027N008N050N018: std_logic_vector(   0 downto 0);
        signal cVar1S9S11N027P039P020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S11N027P039P020N005: std_logic_vector(   0 downto 0);
        signal cVar1S11S11N027P039N020P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S11N027P039N020P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S11N027P039N020P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S11N027P039N020P013: std_logic_vector(   0 downto 0);
        signal cVar1S15S11N027N039P020P034: std_logic_vector(   0 downto 0);
        signal cVar1S16S11N027N039P020P034: std_logic_vector(   0 downto 0);
        signal cVar1S17S11N027N039P020N034: std_logic_vector(   0 downto 0);
        signal cVar1S18S11N027N039P020N034: std_logic_vector(   0 downto 0);
        signal cVar1S19S11N027N039P020N034: std_logic_vector(   0 downto 0);
        signal cVar1S20S11N027N039P020P040: std_logic_vector(   0 downto 0);
        signal cVar1S21S11N027N039P020P040: std_logic_vector(   0 downto 0);
        signal cVar1S22S11N027N039P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S23S11N027N039P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S0S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S1S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S2S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S3S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S4S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S5S12P035P068P032P015: std_logic_vector(   0 downto 0);
        signal cVar1S6S12P035P068N032P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S12P035P068N032P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S12P035P068N032P036: std_logic_vector(   0 downto 0);
        signal cVar1S9S12P035P068N032P036: std_logic_vector(   0 downto 0);
        signal cVar1S10S12P035P068N032N036: std_logic_vector(   0 downto 0);
        signal cVar1S11S12P035P068N032N036: std_logic_vector(   0 downto 0);
        signal cVar1S12S12P035P068N032N036: std_logic_vector(   0 downto 0);
        signal cVar1S13S12P035P068N032N036: std_logic_vector(   0 downto 0);
        signal cVar1S14S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S18S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S19S12P035P068P028P067: std_logic_vector(   0 downto 0);
        signal cVar1S20S12P035P068P028P018: std_logic_vector(   0 downto 0);
        signal cVar1S21S12P035P068P028P018: std_logic_vector(   0 downto 0);
        signal cVar1S22S12P035P068P028P018: std_logic_vector(   0 downto 0);
        signal cVar1S23S12P035P068P028P018: std_logic_vector(   0 downto 0);
        signal cVar1S24S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S25S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S26S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S28S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S29S12P035P067P066P061: std_logic_vector(   0 downto 0);
        signal cVar1S30S12P035P067P066P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S12P035P067P066P037: std_logic_vector(   0 downto 0);
        signal cVar1S32S12P035P067P066N037: std_logic_vector(   0 downto 0);
        signal cVar1S33S12P035P067P068P014: std_logic_vector(   0 downto 0);
        signal cVar1S34S12P035P067P068P014: std_logic_vector(   0 downto 0);
        signal cVar1S35S12P035P067P068P014: std_logic_vector(   0 downto 0);
        signal cVar1S36S12P035P067N068P018: std_logic_vector(   0 downto 0);
        signal cVar1S37S12P035P067N068P018: std_logic_vector(   0 downto 0);
        signal cVar1S38S12P035P067N068P018: std_logic_vector(   0 downto 0);
        signal cVar1S0S13P064P037P029P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S13P064P037P029P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S13P064P037P029N010: std_logic_vector(   0 downto 0);
        signal cVar1S3S13P064P037P029N010: std_logic_vector(   0 downto 0);
        signal cVar1S4S13P064P037P029N010: std_logic_vector(   0 downto 0);
        signal cVar1S5S13P064P037N029P046: std_logic_vector(   0 downto 0);
        signal cVar1S6S13P064P037N029P046: std_logic_vector(   0 downto 0);
        signal cVar1S7S13P064P037N029P046: std_logic_vector(   0 downto 0);
        signal cVar1S8S13P064P037N029N046: std_logic_vector(   0 downto 0);
        signal cVar1S9S13P064P037N029N046: std_logic_vector(   0 downto 0);
        signal cVar1S10S13P064P037N029N046: std_logic_vector(   0 downto 0);
        signal cVar1S11S13P064P037P067P066: std_logic_vector(   0 downto 0);
        signal cVar1S12S13P064P037P067P066: std_logic_vector(   0 downto 0);
        signal cVar1S13S13P064P037P067N066: std_logic_vector(   0 downto 0);
        signal cVar1S14S13P064P037P067N066: std_logic_vector(   0 downto 0);
        signal cVar1S15S13P064P037P067N066: std_logic_vector(   0 downto 0);
        signal cVar1S16S13P064P037N067P060: std_logic_vector(   0 downto 0);
        signal cVar1S17S13P064P037N067P060: std_logic_vector(   0 downto 0);
        signal cVar1S18S13P064P037N067N060: std_logic_vector(   0 downto 0);
        signal cVar1S19S13P064P037N067N060: std_logic_vector(   0 downto 0);
        signal cVar1S20S13P064P037N067N060: std_logic_vector(   0 downto 0);
        signal cVar1S21S13P064P010P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S22S13P064P010P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S23S13P064P010P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S24S13P064P010P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S25S13P064P010P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S26S13P064P010P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S27S13P064P010P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S28S13P064P010P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S29S13P064P010P063N018: std_logic_vector(   0 downto 0);
        signal cVar1S30S13P064P010P063N018: std_logic_vector(   0 downto 0);
        signal cVar1S31S13P064P010P063N018: std_logic_vector(   0 downto 0);
        signal cVar1S32S13P064P010P063N018: std_logic_vector(   0 downto 0);
        signal cVar1S33S13P064P010P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar1S34S13P064P010N032P061: std_logic_vector(   0 downto 0);
        signal cVar1S35S13P064P010N032P061: std_logic_vector(   0 downto 0);
        signal cVar1S36S13P064P010N032P061: std_logic_vector(   0 downto 0);
        signal cVar1S0S14P030P057P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S6S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S7S14P030P057N063P013: std_logic_vector(   0 downto 0);
        signal cVar1S8S14P030N057P056P037: std_logic_vector(   0 downto 0);
        signal cVar1S9S14P030N057P056P037: std_logic_vector(   0 downto 0);
        signal cVar1S10S14P030N057P056P037: std_logic_vector(   0 downto 0);
        signal cVar1S11S14P030N057N056P061: std_logic_vector(   0 downto 0);
        signal cVar1S12S14P030N057N056P061: std_logic_vector(   0 downto 0);
        signal cVar1S13S14P030N057N056N061: std_logic_vector(   0 downto 0);
        signal cVar1S14S14N030P029P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S15S14N030P029P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S16S14N030P029P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S17S14N030P029P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S18S14N030P029N010P053: std_logic_vector(   0 downto 0);
        signal cVar1S19S14N030P029N010P053: std_logic_vector(   0 downto 0);
        signal cVar1S20S14N030P029N010P053: std_logic_vector(   0 downto 0);
        signal cVar1S21S14N030P029N010N053: std_logic_vector(   0 downto 0);
        signal cVar1S22S14N030P029N010N053: std_logic_vector(   0 downto 0);
        signal cVar1S23S14N030N029P046P068: std_logic_vector(   0 downto 0);
        signal cVar1S24S14N030N029P046P068: std_logic_vector(   0 downto 0);
        signal cVar1S25S14N030N029P046P068: std_logic_vector(   0 downto 0);
        signal cVar1S26S14N030N029P046P068: std_logic_vector(   0 downto 0);
        signal cVar1S27S14N030N029P046P068: std_logic_vector(   0 downto 0);
        signal cVar1S28S14N030N029N046P037: std_logic_vector(   0 downto 0);
        signal cVar1S29S14N030N029N046P037: std_logic_vector(   0 downto 0);
        signal cVar1S30S14N030N029N046P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S14N030N029N046N037: std_logic_vector(   0 downto 0);
        signal cVar1S32S14N030N029N046N037: std_logic_vector(   0 downto 0);
        signal cVar1S33S14N030N029N046N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S15P037P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S15P037P039N020P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S15P037P039N020N022: std_logic_vector(   0 downto 0);
        signal cVar1S3S15P037P039N020N022: std_logic_vector(   0 downto 0);
        signal cVar1S4S15P037P039N020N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S15P037N039P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S6S15P037N039P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S15P037N039P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S8S15P037N039P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S9S15P037N039N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S10S15P037N039N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S11S15P037N039N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S15P037N039N027N026: std_logic_vector(   0 downto 0);
        signal cVar1S13S15P037N039N027N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S15P037N039N027N026: std_logic_vector(   0 downto 0);
        signal cVar1S15S15P037P030P057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S15P037P030P057N016: std_logic_vector(   0 downto 0);
        signal cVar1S17S15P037P030P057N016: std_logic_vector(   0 downto 0);
        signal cVar1S18S15P037P030P057N016: std_logic_vector(   0 downto 0);
        signal cVar1S19S15P037P030N057P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S15P037P030N057P065: std_logic_vector(   0 downto 0);
        signal cVar1S21S15P037N030P055P009: std_logic_vector(   0 downto 0);
        signal cVar1S22S15P037N030P055P009: std_logic_vector(   0 downto 0);
        signal cVar1S23S15P037N030P055P009: std_logic_vector(   0 downto 0);
        signal cVar1S24S15P037N030P055N009: std_logic_vector(   0 downto 0);
        signal cVar1S25S15P037N030P055N009: std_logic_vector(   0 downto 0);
        signal cVar1S26S15P037N030P055N009: std_logic_vector(   0 downto 0);
        signal cVar1S27S15P037N030P055P031: std_logic_vector(   0 downto 0);
        signal cVar1S28S15P037N030P055P031: std_logic_vector(   0 downto 0);
        signal cVar1S29S15P037N030P055N031: std_logic_vector(   0 downto 0);
        signal cVar1S30S15P037N030P055N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S16P043P022P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S16P043P022N007P019: std_logic_vector(   0 downto 0);
        signal cVar1S2S16P043P022N007P019: std_logic_vector(   0 downto 0);
        signal cVar1S3S16P043P022N007N019: std_logic_vector(   0 downto 0);
        signal cVar1S4S16P043P022N007N019: std_logic_vector(   0 downto 0);
        signal cVar1S5S16P043N022P062P016nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S16P043N022P062N016: std_logic_vector(   0 downto 0);
        signal cVar1S7S16P043N022N062P006: std_logic_vector(   0 downto 0);
        signal cVar1S8S16P043N022N062P006: std_logic_vector(   0 downto 0);
        signal cVar1S9S16P043N022N062N006: std_logic_vector(   0 downto 0);
        signal cVar1S10S16N043P030P057P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S16N043P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S16N043P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S13S16N043P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S14S16N043P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S15S16N043P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S16S16N043P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S17S16N043P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S18S16N043P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S19S16N043P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S20S16N043N030P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S21S16N043N030P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S22S16N043N030P039N020: std_logic_vector(   0 downto 0);
        signal cVar1S23S16N043N030P039N020: std_logic_vector(   0 downto 0);
        signal cVar1S24S16N043N030N039P034: std_logic_vector(   0 downto 0);
        signal cVar1S25S16N043N030N039P034: std_logic_vector(   0 downto 0);
        signal cVar1S26S16N043N030N039P034: std_logic_vector(   0 downto 0);
        signal cVar1S27S16N043N030N039P034: std_logic_vector(   0 downto 0);
        signal cVar1S28S16N043N030N039N034: std_logic_vector(   0 downto 0);
        signal cVar1S29S16N043N030N039N034: std_logic_vector(   0 downto 0);
        signal cVar1S30S16N043N030N039N034: std_logic_vector(   0 downto 0);
        signal cVar1S31S16N043N030N039N034: std_logic_vector(   0 downto 0);
        signal cVar1S0S17P001P032P068P031: std_logic_vector(   0 downto 0);
        signal cVar1S1S17P001P032P068P031: std_logic_vector(   0 downto 0);
        signal cVar1S2S17P001P032P068P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S17P001P032P068P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S17P001P032P068P031: std_logic_vector(   0 downto 0);
        signal cVar1S5S17P001P032P068P066: std_logic_vector(   0 downto 0);
        signal cVar1S6S17P001P032P068P066: std_logic_vector(   0 downto 0);
        signal cVar1S7S17P001P032P068P066: std_logic_vector(   0 downto 0);
        signal cVar1S8S17P001P032P068N066: std_logic_vector(   0 downto 0);
        signal cVar1S9S17P001N032P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S10S17P001N032P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S11S17P001N032P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S17P001N032P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S13S17P001N032P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S14S17P001N032P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S15S17P001N032P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S16S17P001N032P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S17S17P001N032P000P069: std_logic_vector(   0 downto 0);
        signal cVar1S18S17P001N032P000P069: std_logic_vector(   0 downto 0);
        signal cVar1S19S17P001N032P000P069: std_logic_vector(   0 downto 0);
        signal cVar1S20S17P001N032P000N069: std_logic_vector(   0 downto 0);
        signal cVar1S21S17P001N032P000N069: std_logic_vector(   0 downto 0);
        signal cVar1S22S17P001N032P000N069: std_logic_vector(   0 downto 0);
        signal cVar1S23S17P001N032P000N069: std_logic_vector(   0 downto 0);
        signal cVar1S24S17P001P015P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S17P001P015N041P059: std_logic_vector(   0 downto 0);
        signal cVar1S26S17P001P015N041P059: std_logic_vector(   0 downto 0);
        signal cVar1S27S17P001P015N041P059: std_logic_vector(   0 downto 0);
        signal cVar1S28S17P001P015N041P059: std_logic_vector(   0 downto 0);
        signal cVar1S29S17P001P015P012P066: std_logic_vector(   0 downto 0);
        signal cVar1S30S17P001P015P012P066: std_logic_vector(   0 downto 0);
        signal cVar1S31S17P001P015P012P066: std_logic_vector(   0 downto 0);
        signal cVar1S32S17P001P015N012P063: std_logic_vector(   0 downto 0);
        signal cVar1S0S18P067P037P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S1S18P067P037P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S2S18P067P037P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S18P067P037P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S18P067P037P069N031: std_logic_vector(   0 downto 0);
        signal cVar1S5S18P067P037P069N031: std_logic_vector(   0 downto 0);
        signal cVar1S6S18P067P037P069N031: std_logic_vector(   0 downto 0);
        signal cVar1S7S18P067P037P069N031: std_logic_vector(   0 downto 0);
        signal cVar1S8S18P067P037P069P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S18P067P037P069P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S18P067P037P069N017: std_logic_vector(   0 downto 0);
        signal cVar1S11S18P067P037P069N017: std_logic_vector(   0 downto 0);
        signal cVar1S12S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S14S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S15S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S18P067P037P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S18S18P067P037N016P019: std_logic_vector(   0 downto 0);
        signal cVar1S19S18P067P037N016P019: std_logic_vector(   0 downto 0);
        signal cVar1S20S18P067P037N016N019: std_logic_vector(   0 downto 0);
        signal cVar1S21S18P067P037N016N019: std_logic_vector(   0 downto 0);
        signal cVar1S22S18P067P037N016N019: std_logic_vector(   0 downto 0);
        signal cVar1S23S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S24S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S25S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S26S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S27S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S28S18P067P007P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S29S18P067P007N069P018: std_logic_vector(   0 downto 0);
        signal cVar1S30S18P067P007N069P018: std_logic_vector(   0 downto 0);
        signal cVar1S31S18P067P007N069N018: std_logic_vector(   0 downto 0);
        signal cVar1S32S18P067P007N069N018: std_logic_vector(   0 downto 0);
        signal cVar1S33S18P067P007P049nsss: std_logic_vector(   0 downto 0);
        signal cVar1S34S18P067P007N049P044: std_logic_vector(   0 downto 0);
        signal cVar1S0S19P031P012P008P060: std_logic_vector(   0 downto 0);
        signal cVar1S1S19P031P012P008P060: std_logic_vector(   0 downto 0);
        signal cVar1S2S19P031P012P008N060: std_logic_vector(   0 downto 0);
        signal cVar1S3S19P031P012P008N060: std_logic_vector(   0 downto 0);
        signal cVar1S4S19P031P012P008N060: std_logic_vector(   0 downto 0);
        signal cVar1S5S19P031P012P008P033: std_logic_vector(   0 downto 0);
        signal cVar1S6S19P031P012P008P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S19P031N012P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S8S19P031N012P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S19P031N012P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S19P031N012P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S11S19P031N012P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S12S19P031N012N013P054: std_logic_vector(   0 downto 0);
        signal cVar1S13S19P031N012N013P054: std_logic_vector(   0 downto 0);
        signal cVar1S14S19P031N012N013N054: std_logic_vector(   0 downto 0);
        signal cVar1S15S19P031N012N013N054: std_logic_vector(   0 downto 0);
        signal cVar1S16S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S17S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S18S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S19S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S20S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S19N031P036P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S19N031P036P007P008: std_logic_vector(   0 downto 0);
        signal cVar1S23S19N031P036P007P008: std_logic_vector(   0 downto 0);
        signal cVar1S24S19N031P036P007P008: std_logic_vector(   0 downto 0);
        signal cVar1S25S19N031N036P045P007: std_logic_vector(   0 downto 0);
        signal cVar1S26S19N031N036P045P007: std_logic_vector(   0 downto 0);
        signal cVar1S27S19N031N036P045P007: std_logic_vector(   0 downto 0);
        signal cVar1S28S19N031N036P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S29S19N031N036P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S30S19N031N036P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S31S19N031N036N045P053: std_logic_vector(   0 downto 0);
        signal cVar1S32S19N031N036N045P053: std_logic_vector(   0 downto 0);
        signal cVar1S33S19N031N036N045P053: std_logic_vector(   0 downto 0);
        signal cVar1S34S19N031N036N045N053: std_logic_vector(   0 downto 0);
        signal cVar1S35S19N031N036N045N053: std_logic_vector(   0 downto 0);
        signal cVar1S36S19N031N036N045N053: std_logic_vector(   0 downto 0);
        signal cVar1S0S20P032P031P016P013: std_logic_vector(   0 downto 0);
        signal cVar1S1S20P032P031P016P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S20P032P031P016P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S20P032P031P016P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S20P032P031P016P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S20P032P031N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S6S20P032P031N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S7S20P032P031N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S20P032P031N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S9S20P032P031N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S10S20P032P031N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S11S20P032P031P003P018: std_logic_vector(   0 downto 0);
        signal cVar1S12S20P032P031P003N018: std_logic_vector(   0 downto 0);
        signal cVar1S13S20N032P036P024P047: std_logic_vector(   0 downto 0);
        signal cVar1S14S20N032P036P024P047: std_logic_vector(   0 downto 0);
        signal cVar1S15S20N032P036P024P047: std_logic_vector(   0 downto 0);
        signal cVar1S16S20N032P036P024N047: std_logic_vector(   0 downto 0);
        signal cVar1S17S20N032P036P024N047: std_logic_vector(   0 downto 0);
        signal cVar1S18S20N032P036P024N047: std_logic_vector(   0 downto 0);
        signal cVar1S19S20N032P036N024P019: std_logic_vector(   0 downto 0);
        signal cVar1S20S20N032P036N024P019: std_logic_vector(   0 downto 0);
        signal cVar1S21S20N032P036N024P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S20N032P036N024P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S20N032P036N024N019: std_logic_vector(   0 downto 0);
        signal cVar1S24S20N032P036N024N019: std_logic_vector(   0 downto 0);
        signal cVar1S25S20N032P036N024N019: std_logic_vector(   0 downto 0);
        signal cVar1S26S20N032P036N024N019: std_logic_vector(   0 downto 0);
        signal cVar1S27S20N032P036P010P029: std_logic_vector(   0 downto 0);
        signal cVar1S28S20N032P036P010P029: std_logic_vector(   0 downto 0);
        signal cVar1S29S20N032P036P010P029: std_logic_vector(   0 downto 0);
        signal cVar1S30S20N032P036P010P029: std_logic_vector(   0 downto 0);
        signal cVar1S31S20N032P036P010P029: std_logic_vector(   0 downto 0);
        signal cVar1S32S20N032P036P010P055: std_logic_vector(   0 downto 0);
        signal cVar1S33S20N032P036P010P055: std_logic_vector(   0 downto 0);
        signal cVar1S34S20N032P036P010N055: std_logic_vector(   0 downto 0);
        signal cVar1S0S21P024P047P066P063: std_logic_vector(   0 downto 0);
        signal cVar1S1S21P024P047P066P063: std_logic_vector(   0 downto 0);
        signal cVar1S2S21P024P047P066P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S21P024P047P066P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S21P024P047P066N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S21P024N047P010P043: std_logic_vector(   0 downto 0);
        signal cVar1S6S21P024N047P010P043: std_logic_vector(   0 downto 0);
        signal cVar1S7S21P024N047P010N043: std_logic_vector(   0 downto 0);
        signal cVar1S8S21P024N047P010N043: std_logic_vector(   0 downto 0);
        signal cVar1S9S21P024N047P010N043: std_logic_vector(   0 downto 0);
        signal cVar1S10S21P024N047P010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S21P024N047P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S12S21N024P030P057P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S21N024P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S14S21N024P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S15S21N024P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S16S21N024P030P057N063: std_logic_vector(   0 downto 0);
        signal cVar1S17S21N024P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S18S21N024P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S19S21N024P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S20S21N024P030N057P029: std_logic_vector(   0 downto 0);
        signal cVar1S21S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S24S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S25S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S21N024N030P031P019: std_logic_vector(   0 downto 0);
        signal cVar1S27S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S28S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S29S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S30S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S31S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S32S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S33S21N024N030N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S0S22P024P047P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S22P024P047P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S22P024P047P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S22P024N047P010P001: std_logic_vector(   0 downto 0);
        signal cVar1S4S22P024N047P010P001: std_logic_vector(   0 downto 0);
        signal cVar1S5S22P024N047P010P001: std_logic_vector(   0 downto 0);
        signal cVar1S6S22P024N047P010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S22P024N047P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S8S22N024P067P017P022: std_logic_vector(   0 downto 0);
        signal cVar1S9S22N024P067P017P022: std_logic_vector(   0 downto 0);
        signal cVar1S10S22N024P067P017P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S22N024P067P017N022: std_logic_vector(   0 downto 0);
        signal cVar1S12S22N024P067P017N022: std_logic_vector(   0 downto 0);
        signal cVar1S13S22N024P067P017P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S22N024P067P017P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S22N024P067P017N014: std_logic_vector(   0 downto 0);
        signal cVar1S16S22N024P067P017N014: std_logic_vector(   0 downto 0);
        signal cVar1S17S22N024P067P017N014: std_logic_vector(   0 downto 0);
        signal cVar1S18S22N024P067P017N014: std_logic_vector(   0 downto 0);
        signal cVar1S19S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S20S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S21S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S22S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S23S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S24S22N024P067P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S25S22N024P067N060P064: std_logic_vector(   0 downto 0);
        signal cVar1S26S22N024P067N060P064: std_logic_vector(   0 downto 0);
        signal cVar1S27S22N024P067N060P064: std_logic_vector(   0 downto 0);
        signal cVar1S28S22N024P067N060N064: std_logic_vector(   0 downto 0);
        signal cVar1S29S22N024P067N060N064: std_logic_vector(   0 downto 0);
        signal cVar1S30S22N024P067N060N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S23P024P047P066P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S23P024P047P066P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S23P024P047P066N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S23P024P047P066N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S23P024N047P010P049: std_logic_vector(   0 downto 0);
        signal cVar1S5S23P024N047P010P049: std_logic_vector(   0 downto 0);
        signal cVar1S6S23P024N047P010P049: std_logic_vector(   0 downto 0);
        signal cVar1S7S23P024N047P010P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S23N024P069P047P007: std_logic_vector(   0 downto 0);
        signal cVar1S9S23N024P069P047P007: std_logic_vector(   0 downto 0);
        signal cVar1S10S23N024P069P047P007: std_logic_vector(   0 downto 0);
        signal cVar1S11S23N024P069P047P007: std_logic_vector(   0 downto 0);
        signal cVar1S12S23N024P069P047P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S23N024P069P047P063: std_logic_vector(   0 downto 0);
        signal cVar1S14S23N024P069P047P063: std_logic_vector(   0 downto 0);
        signal cVar1S15S23N024N069P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S23N024N069P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S17S23N024N069P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S18S23N024N069N022P036: std_logic_vector(   0 downto 0);
        signal cVar1S19S23N024N069N022P036: std_logic_vector(   0 downto 0);
        signal cVar1S20S23N024N069N022N036: std_logic_vector(   0 downto 0);
        signal cVar1S21S23N024N069N022N036: std_logic_vector(   0 downto 0);
        signal cVar1S22S23N024N069N022N036: std_logic_vector(   0 downto 0);
        signal cVar1S0S24P024P047P066P060: std_logic_vector(   0 downto 0);
        signal cVar1S1S24P024P047P066P060: std_logic_vector(   0 downto 0);
        signal cVar1S2S24P024P047P066P060psss: std_logic_vector(   0 downto 0);
        signal cVar1S3S24P024P047P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S24P024P047P066N069: std_logic_vector(   0 downto 0);
        signal cVar1S5S24P024P047P066N069: std_logic_vector(   0 downto 0);
        signal cVar1S6S24P024N047P010P064: std_logic_vector(   0 downto 0);
        signal cVar1S7S24P024N047P010P064: std_logic_vector(   0 downto 0);
        signal cVar1S8S24P024N047P010P064: std_logic_vector(   0 downto 0);
        signal cVar1S9S24P024N047P010N064: std_logic_vector(   0 downto 0);
        signal cVar1S10S24P024N047P010N064: std_logic_vector(   0 downto 0);
        signal cVar1S11S24P024N047P010N064: std_logic_vector(   0 downto 0);
        signal cVar1S12S24P024N047P010P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S24P024N047P010N025: std_logic_vector(   0 downto 0);
        signal cVar1S14S24N024P040P021P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S24N024P040N021P037: std_logic_vector(   0 downto 0);
        signal cVar1S16S24N024P040N021P037: std_logic_vector(   0 downto 0);
        signal cVar1S17S24N024P040N021P037: std_logic_vector(   0 downto 0);
        signal cVar1S18S24N024P040N021N037: std_logic_vector(   0 downto 0);
        signal cVar1S19S24N024P040N021N037: std_logic_vector(   0 downto 0);
        signal cVar1S20S24N024P040N021N037: std_logic_vector(   0 downto 0);
        signal cVar1S21S24N024N040P002P039: std_logic_vector(   0 downto 0);
        signal cVar1S22S24N024N040P002P039: std_logic_vector(   0 downto 0);
        signal cVar1S23S24N024N040P002P039: std_logic_vector(   0 downto 0);
        signal cVar1S24S24N024N040P002N039: std_logic_vector(   0 downto 0);
        signal cVar1S25S24N024N040P002N039: std_logic_vector(   0 downto 0);
        signal cVar1S26S24N024N040P002P053: std_logic_vector(   0 downto 0);
        signal cVar1S27S24N024N040P002N053: std_logic_vector(   0 downto 0);
        signal cVar1S28S24N024N040P002N053: std_logic_vector(   0 downto 0);
        signal cVar1S0S25P001P031P012P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S25P001P031P012P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S25P001P031P012P062: std_logic_vector(   0 downto 0);
        signal cVar1S3S25P001P031P012P062: std_logic_vector(   0 downto 0);
        signal cVar1S4S25P001P031P012P062: std_logic_vector(   0 downto 0);
        signal cVar1S5S25P001P031N012P013: std_logic_vector(   0 downto 0);
        signal cVar1S6S25P001P031N012P013: std_logic_vector(   0 downto 0);
        signal cVar1S7S25P001P031N012N013: std_logic_vector(   0 downto 0);
        signal cVar1S8S25P001P031N012N013: std_logic_vector(   0 downto 0);
        signal cVar1S9S25P001N031P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S25P001N031P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S25P001N031P030N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S25P001N031P030N063: std_logic_vector(   0 downto 0);
        signal cVar1S13S25P001N031P030N063: std_logic_vector(   0 downto 0);
        signal cVar1S14S25P001N031P030N063: std_logic_vector(   0 downto 0);
        signal cVar1S15S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S20S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S21S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S22S25P001N031N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S23S25P001P023P067P012: std_logic_vector(   0 downto 0);
        signal cVar1S24S25P001P023P067N012: std_logic_vector(   0 downto 0);
        signal cVar1S25S25P001P023P067N012: std_logic_vector(   0 downto 0);
        signal cVar1S26S25P001P023N067P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S27S25P001P023N067N041: std_logic_vector(   0 downto 0);
        signal cVar1S28S25P001P023N067N041: std_logic_vector(   0 downto 0);
        signal cVar1S29S25P001P023N067N041: std_logic_vector(   0 downto 0);
        signal cVar1S0S26P015P017P034P058: std_logic_vector(   0 downto 0);
        signal cVar1S1S26P015P017P034P058: std_logic_vector(   0 downto 0);
        signal cVar1S2S26P015P017P034P058: std_logic_vector(   0 downto 0);
        signal cVar1S3S26P015P017N034P033: std_logic_vector(   0 downto 0);
        signal cVar1S4S26P015P017N034N033: std_logic_vector(   0 downto 0);
        signal cVar1S5S26P015P017N034N033: std_logic_vector(   0 downto 0);
        signal cVar1S6S26P015P017N034N033: std_logic_vector(   0 downto 0);
        signal cVar1S7S26P015P017N034N033: std_logic_vector(   0 downto 0);
        signal cVar1S8S26P015P017P006P001: std_logic_vector(   0 downto 0);
        signal cVar1S9S26P015P017P006P001: std_logic_vector(   0 downto 0);
        signal cVar1S10S26P015P017P006P001: std_logic_vector(   0 downto 0);
        signal cVar1S11S26P015P017P006P001: std_logic_vector(   0 downto 0);
        signal cVar1S12S26P015P017P006P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S26P015P017P006P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S26P015P017P006N062: std_logic_vector(   0 downto 0);
        signal cVar1S15S26P015P017P006N062: std_logic_vector(   0 downto 0);
        signal cVar1S16S26P015P017P006N062: std_logic_vector(   0 downto 0);
        signal cVar1S17S26N015P031P012P017: std_logic_vector(   0 downto 0);
        signal cVar1S18S26N015P031P012P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S26N015P031P012N017: std_logic_vector(   0 downto 0);
        signal cVar1S20S26N015P031P012N017: std_logic_vector(   0 downto 0);
        signal cVar1S21S26N015P031P012N017: std_logic_vector(   0 downto 0);
        signal cVar1S22S26N015P031N012P014: std_logic_vector(   0 downto 0);
        signal cVar1S23S26N015P031N012P014: std_logic_vector(   0 downto 0);
        signal cVar1S24S26N015P031N012P014: std_logic_vector(   0 downto 0);
        signal cVar1S25S26N015P031N012N014: std_logic_vector(   0 downto 0);
        signal cVar1S26S26N015P031N012N014: std_logic_vector(   0 downto 0);
        signal cVar1S27S26N015P031N012N014: std_logic_vector(   0 downto 0);
        signal cVar1S28S26N015P031N012N014: std_logic_vector(   0 downto 0);
        signal cVar1S29S26N015N031P030P059: std_logic_vector(   0 downto 0);
        signal cVar1S30S26N015N031P030P059: std_logic_vector(   0 downto 0);
        signal cVar1S31S26N015N031P030P059: std_logic_vector(   0 downto 0);
        signal cVar1S32S26N015N031P030N059: std_logic_vector(   0 downto 0);
        signal cVar1S33S26N015N031P030N059: std_logic_vector(   0 downto 0);
        signal cVar1S34S26N015N031P030N059: std_logic_vector(   0 downto 0);
        signal cVar1S35S26N015N031N030P007: std_logic_vector(   0 downto 0);
        signal cVar1S36S26N015N031N030P007: std_logic_vector(   0 downto 0);
        signal cVar1S37S26N015N031N030P007: std_logic_vector(   0 downto 0);
        signal cVar1S38S26N015N031N030N007: std_logic_vector(   0 downto 0);
        signal cVar1S39S26N015N031N030N007: std_logic_vector(   0 downto 0);
        signal cVar1S40S26N015N031N030N007: std_logic_vector(   0 downto 0);
        signal cVar1S0S27P002P022P043P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S27P002P022P043N007: std_logic_vector(   0 downto 0);
        signal cVar1S2S27P002P022P043N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S27P002P022P043N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S27P002P022N043P042: std_logic_vector(   0 downto 0);
        signal cVar1S5S27P002P022N043P042: std_logic_vector(   0 downto 0);
        signal cVar1S6S27P002P022N043N042: std_logic_vector(   0 downto 0);
        signal cVar1S7S27P002P022N043N042: std_logic_vector(   0 downto 0);
        signal cVar1S8S27P002N022P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S9S27P002N022P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S10S27P002N022P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S11S27P002N022P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S27P002N022N027P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S27P002N022N027P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S27P002N022N027P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S27P002N022N027N032: std_logic_vector(   0 downto 0);
        signal cVar1S16S27P002N022N027N032: std_logic_vector(   0 downto 0);
        signal cVar1S17S27P002N022N027N032: std_logic_vector(   0 downto 0);
        signal cVar1S18S27P002N022N027N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S27P002P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S27P002P040N021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S27P002N040P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S22S27P002N040P050N048: std_logic_vector(   0 downto 0);
        signal cVar1S23S27P002N040P050N048: std_logic_vector(   0 downto 0);
        signal cVar1S0S28P032P002P016P049: std_logic_vector(   0 downto 0);
        signal cVar1S1S28P032P002P016P049: std_logic_vector(   0 downto 0);
        signal cVar1S2S28P032P002N016P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S28P032P002N016P063: std_logic_vector(   0 downto 0);
        signal cVar1S4S28P032P002N016P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S28P032P002N016N063: std_logic_vector(   0 downto 0);
        signal cVar1S6S28P032P002N016N063: std_logic_vector(   0 downto 0);
        signal cVar1S7S28P032P002N016N063: std_logic_vector(   0 downto 0);
        signal cVar1S8S28P032P002N016N063: std_logic_vector(   0 downto 0);
        signal cVar1S9S28P032P002P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S28N032P027P026P000: std_logic_vector(   0 downto 0);
        signal cVar1S11S28N032P027P026P000: std_logic_vector(   0 downto 0);
        signal cVar1S12S28N032P027P026P000: std_logic_vector(   0 downto 0);
        signal cVar1S13S28N032P027P026P036: std_logic_vector(   0 downto 0);
        signal cVar1S14S28N032P027P026P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S28N032N027P022P069: std_logic_vector(   0 downto 0);
        signal cVar1S16S28N032N027P022P069: std_logic_vector(   0 downto 0);
        signal cVar1S17S28N032N027P022P069: std_logic_vector(   0 downto 0);
        signal cVar1S18S28N032N027P022P069: std_logic_vector(   0 downto 0);
        signal cVar1S19S28N032N027N022P030: std_logic_vector(   0 downto 0);
        signal cVar1S20S28N032N027N022P030: std_logic_vector(   0 downto 0);
        signal cVar1S21S28N032N027N022P030: std_logic_vector(   0 downto 0);
        signal cVar1S22S28N032N027N022N030: std_logic_vector(   0 downto 0);
        signal cVar1S23S28N032N027N022N030: std_logic_vector(   0 downto 0);
        signal cVar1S24S28N032N027N022N030: std_logic_vector(   0 downto 0);
        signal cVar1S0S29P040P021P035P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S29P040P021P035N002: std_logic_vector(   0 downto 0);
        signal cVar1S2S29P040P021P035N002: std_logic_vector(   0 downto 0);
        signal cVar1S3S29P040P021P035N002: std_logic_vector(   0 downto 0);
        signal cVar1S4S29P040N021P037P005: std_logic_vector(   0 downto 0);
        signal cVar1S5S29P040N021P037P005: std_logic_vector(   0 downto 0);
        signal cVar1S6S29P040N021P037P005: std_logic_vector(   0 downto 0);
        signal cVar1S7S29P040N021N037P017: std_logic_vector(   0 downto 0);
        signal cVar1S8S29P040N021N037P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S29P040N021N037N017: std_logic_vector(   0 downto 0);
        signal cVar1S10S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S11S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S12S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S13S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S14S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S15S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S16S29N040P038P021P002: std_logic_vector(   0 downto 0);
        signal cVar1S17S29N040P038P021P010: std_logic_vector(   0 downto 0);
        signal cVar1S18S29N040P038P021P010: std_logic_vector(   0 downto 0);
        signal cVar1S19S29N040P038P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S29N040P038N026N059: std_logic_vector(   0 downto 0);
        signal cVar1S0S30P068P047P049P065: std_logic_vector(   0 downto 0);
        signal cVar1S1S30P068P047P049P065: std_logic_vector(   0 downto 0);
        signal cVar1S2S30P068P047P049P065: std_logic_vector(   0 downto 0);
        signal cVar1S3S30P068P047P049P065: std_logic_vector(   0 downto 0);
        signal cVar1S4S30P068P047P049P065: std_logic_vector(   0 downto 0);
        signal cVar1S5S30P068P047N049P024: std_logic_vector(   0 downto 0);
        signal cVar1S6S30P068P047N049N024: std_logic_vector(   0 downto 0);
        signal cVar1S7S30P068P047N049N024: std_logic_vector(   0 downto 0);
        signal cVar1S8S30P068N047P052P066: std_logic_vector(   0 downto 0);
        signal cVar1S9S30P068N047P052P066: std_logic_vector(   0 downto 0);
        signal cVar1S10S30P068N047P052P066: std_logic_vector(   0 downto 0);
        signal cVar1S11S30P068N047P052P066: std_logic_vector(   0 downto 0);
        signal cVar1S12S30P068N047P052P066: std_logic_vector(   0 downto 0);
        signal cVar1S13S30P068N047N052P036: std_logic_vector(   0 downto 0);
        signal cVar1S14S30P068N047N052P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S30P068N047N052P036: std_logic_vector(   0 downto 0);
        signal cVar1S16S30P068N047N052N036: std_logic_vector(   0 downto 0);
        signal cVar1S17S30P068N047N052N036: std_logic_vector(   0 downto 0);
        signal cVar1S18S30P068N047N052N036: std_logic_vector(   0 downto 0);
        signal cVar1S19S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S23S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S24S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S25S30P068P055P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S26S30P068P055N019P051: std_logic_vector(   0 downto 0);
        signal cVar1S27S30P068P055N019P051: std_logic_vector(   0 downto 0);
        signal cVar1S28S30P068P055N019N051: std_logic_vector(   0 downto 0);
        signal cVar1S29S30P068P055N019N051: std_logic_vector(   0 downto 0);
        signal cVar1S30S30P068P055N019N051: std_logic_vector(   0 downto 0);
        signal cVar1S31S30P068P055P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S32S30P068P055P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S33S30P068P055P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S34S30P068P055N016P049: std_logic_vector(   0 downto 0);
        signal cVar1S35S30P068P055N016P049: std_logic_vector(   0 downto 0);
        signal cVar1S36S30P068P055N016P049: std_logic_vector(   0 downto 0);
        signal cVar1S37S30P068P055N016P049: std_logic_vector(   0 downto 0);
        signal cVar1S0S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S1S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S2S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S3S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S4S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S5S31P036P063P005P048: std_logic_vector(   0 downto 0);
        signal cVar1S6S31P036P063P005P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S31P036P063P005N035: std_logic_vector(   0 downto 0);
        signal cVar1S8S31P036N063P016P064: std_logic_vector(   0 downto 0);
        signal cVar1S9S31P036N063P016P064: std_logic_vector(   0 downto 0);
        signal cVar1S10S31P036N063P016P064: std_logic_vector(   0 downto 0);
        signal cVar1S11S31P036N063P016P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S31P036N063P016N064: std_logic_vector(   0 downto 0);
        signal cVar1S13S31P036N063P016N064: std_logic_vector(   0 downto 0);
        signal cVar1S14S31P036N063P016N064: std_logic_vector(   0 downto 0);
        signal cVar1S15S31P036N063P016N064: std_logic_vector(   0 downto 0);
        signal cVar1S16S31P036N063N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S31P036N063N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S18S31P036N063N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S19S31P036N063N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S20S31P036N063N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S31P036N063N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S22S31N036P052P068P048: std_logic_vector(   0 downto 0);
        signal cVar1S23S31N036P052P068P048: std_logic_vector(   0 downto 0);
        signal cVar1S24S31N036P052P068P048: std_logic_vector(   0 downto 0);
        signal cVar1S25S31N036P052P068P048: std_logic_vector(   0 downto 0);
        signal cVar1S26S31N036P052P068P048: std_logic_vector(   0 downto 0);
        signal cVar1S27S31N036P052P068P055: std_logic_vector(   0 downto 0);
        signal cVar1S28S31N036P052P068P055: std_logic_vector(   0 downto 0);
        signal cVar1S29S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S30S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S31S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S32S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S33S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S34S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S35S31N036N052P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S36S31N036N052N018P014: std_logic_vector(   0 downto 0);
        signal cVar1S37S31N036N052N018P014: std_logic_vector(   0 downto 0);
        signal cVar1S38S31N036N052N018P014: std_logic_vector(   0 downto 0);
        signal cVar1S39S31N036N052N018P014: std_logic_vector(   0 downto 0);
        signal cVar1S40S31N036N052N018N014: std_logic_vector(   0 downto 0);
        signal cVar1S41S31N036N052N018N014: std_logic_vector(   0 downto 0);
        signal cVar1S42S31N036N052N018N014: std_logic_vector(   0 downto 0);
        signal cVar1S43S31N036N052N018N014: std_logic_vector(   0 downto 0);
        signal cVar1S0S32P036P066P006P027: std_logic_vector(   0 downto 0);
        signal cVar1S1S32P036P066P006P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S32P036P066P006P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S32P036P066P006P059: std_logic_vector(   0 downto 0);
        signal cVar1S4S32P036N066P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S5S32P036N066P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S6S32P036N066P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S7S32P036N066P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S32P036N066P016P018: std_logic_vector(   0 downto 0);
        signal cVar1S9S32P036N066N016P068: std_logic_vector(   0 downto 0);
        signal cVar1S10S32P036N066N016P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S32P036N066N016P068: std_logic_vector(   0 downto 0);
        signal cVar1S12S32P036N066N016P068: std_logic_vector(   0 downto 0);
        signal cVar1S13S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S14S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S15S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S18S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S19S32N036P060P048P063: std_logic_vector(   0 downto 0);
        signal cVar1S20S32N036P060P048P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S32N036P060P048N006: std_logic_vector(   0 downto 0);
        signal cVar1S22S32N036N060P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S23S32N036N060P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S24S32N036N060P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S25S32N036N060P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S26S32N036N060P058N054: std_logic_vector(   0 downto 0);
        signal cVar1S27S32N036N060P058N054: std_logic_vector(   0 downto 0);
        signal cVar1S28S32N036N060P058N054: std_logic_vector(   0 downto 0);
        signal cVar1S29S32N036N060P058P056: std_logic_vector(   0 downto 0);
        signal cVar1S30S32N036N060P058P056: std_logic_vector(   0 downto 0);
        signal cVar1S31S32N036N060P058P056: std_logic_vector(   0 downto 0);
        signal cVar1S32S32N036N060P058N056: std_logic_vector(   0 downto 0);
        signal cVar1S0S33P034P049P026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S33P034P049P026N018: std_logic_vector(   0 downto 0);
        signal cVar1S2S33P034P049P026N018: std_logic_vector(   0 downto 0);
        signal cVar1S3S33P034P049N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S33P034P049N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S5S33P034P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S33P034P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S7S33P034P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S8S33P034N049P028P011: std_logic_vector(   0 downto 0);
        signal cVar1S9S33P034N049P028P011: std_logic_vector(   0 downto 0);
        signal cVar1S10S33P034N049P028N011: std_logic_vector(   0 downto 0);
        signal cVar1S11S33P034N049P028N011: std_logic_vector(   0 downto 0);
        signal cVar1S12S33P034N049P028N011: std_logic_vector(   0 downto 0);
        signal cVar1S13S33P034N049P028N011: std_logic_vector(   0 downto 0);
        signal cVar1S14S33P034N049N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S33P034N049N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S33P034N049N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S17S33P034N049N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S18S33P034N049N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S19S33P034N049N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S20S33P034N049N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S21S33P034P014P044P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S33P034P014P044P069: std_logic_vector(   0 downto 0);
        signal cVar1S23S33P034P014P044P069: std_logic_vector(   0 downto 0);
        signal cVar1S24S33P034P014P044N069: std_logic_vector(   0 downto 0);
        signal cVar1S25S33P034P014P044N069: std_logic_vector(   0 downto 0);
        signal cVar1S26S33P034P014P044N069: std_logic_vector(   0 downto 0);
        signal cVar1S27S33P034N014P045P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S33P034N014P045N062: std_logic_vector(   0 downto 0);
        signal cVar1S29S33P034N014N045P046: std_logic_vector(   0 downto 0);
        signal cVar1S30S33P034N014N045P046: std_logic_vector(   0 downto 0);
        signal cVar1S31S33P034N014N045P046: std_logic_vector(   0 downto 0);
        signal cVar1S0S34P034P068P032P054: std_logic_vector(   0 downto 0);
        signal cVar1S1S34P034P068P032P054: std_logic_vector(   0 downto 0);
        signal cVar1S2S34P034P068P032P054: std_logic_vector(   0 downto 0);
        signal cVar1S3S34P034P068P032P054: std_logic_vector(   0 downto 0);
        signal cVar1S4S34P034P068P032P054: std_logic_vector(   0 downto 0);
        signal cVar1S5S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S6S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S7S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S8S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S34P034P068N032P059: std_logic_vector(   0 downto 0);
        signal cVar1S11S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S16S34P034P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S17S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S18S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S19S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S20S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S21S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S22S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S23S34P034P068P019P036: std_logic_vector(   0 downto 0);
        signal cVar1S24S34P034P062P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S25S34P034P062P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S26S34P034P062P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S27S34P034P062P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S28S34P034P062P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S29S34P034P062P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S30S34P034P062P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S31S34P034P062P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S32S34P034P062P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S33S34P034P062P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S34S34P034P062P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S35S34P034P062P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S36S34P034N062P008P063: std_logic_vector(   0 downto 0);
        signal cVar1S37S34P034N062P008P063: std_logic_vector(   0 downto 0);
        signal cVar1S38S34P034N062P008P063: std_logic_vector(   0 downto 0);
        signal cVar1S39S34P034N062P008N063: std_logic_vector(   0 downto 0);
        signal cVar1S40S34P034N062P008N063: std_logic_vector(   0 downto 0);
        signal cVar1S41S34P034N062P008N063: std_logic_vector(   0 downto 0);
        signal cVar1S42S34P034N062P008P026: std_logic_vector(   0 downto 0);
        signal cVar1S43S34P034N062P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S44S34P034N062P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S0S35P061P064P030P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S35P061P064P030N013: std_logic_vector(   0 downto 0);
        signal cVar1S2S35P061P064P030N013: std_logic_vector(   0 downto 0);
        signal cVar1S3S35P061P064N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S4S35P061P064N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S5S35P061P064N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S6S35P061P064N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S7S35P061P064N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S8S35P061P064P058P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S35P061P064P058N008: std_logic_vector(   0 downto 0);
        signal cVar1S10S35P061P064P058N008: std_logic_vector(   0 downto 0);
        signal cVar1S11S35P061P064P058N008: std_logic_vector(   0 downto 0);
        signal cVar1S12S35P061P064P058P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S35N061P057P026P007: std_logic_vector(   0 downto 0);
        signal cVar1S14S35N061P057P026P007: std_logic_vector(   0 downto 0);
        signal cVar1S15S35N061P057P026P007: std_logic_vector(   0 downto 0);
        signal cVar1S16S35N061P057P026P007: std_logic_vector(   0 downto 0);
        signal cVar1S17S35N061P057P026N030: std_logic_vector(   0 downto 0);
        signal cVar1S18S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S19S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S21S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S22S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S23S35N061N057P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S35N061N057N064P063: std_logic_vector(   0 downto 0);
        signal cVar1S25S35N061N057N064P063: std_logic_vector(   0 downto 0);
        signal cVar1S26S35N061N057N064N063: std_logic_vector(   0 downto 0);
        signal cVar1S27S35N061N057N064N063: std_logic_vector(   0 downto 0);
        signal cVar1S0S36P063P062P065P066: std_logic_vector(   0 downto 0);
        signal cVar1S1S36P063P062P065P066: std_logic_vector(   0 downto 0);
        signal cVar1S2S36P063P062P065P066: std_logic_vector(   0 downto 0);
        signal cVar1S3S36P063P062P065P066: std_logic_vector(   0 downto 0);
        signal cVar1S4S36P063P062P065P066: std_logic_vector(   0 downto 0);
        signal cVar1S5S36P063P062N065P007: std_logic_vector(   0 downto 0);
        signal cVar1S6S36P063P062N065P007: std_logic_vector(   0 downto 0);
        signal cVar1S7S36P063P062N065P007: std_logic_vector(   0 downto 0);
        signal cVar1S8S36P063P062N065P007: std_logic_vector(   0 downto 0);
        signal cVar1S9S36P063P062P048P054: std_logic_vector(   0 downto 0);
        signal cVar1S10S36P063P062P048P054: std_logic_vector(   0 downto 0);
        signal cVar1S11S36P063P062P048P054: std_logic_vector(   0 downto 0);
        signal cVar1S12S36P063P062P048P054: std_logic_vector(   0 downto 0);
        signal cVar1S13S36P063P062P048P054: std_logic_vector(   0 downto 0);
        signal cVar1S14S36P063P062P048P046: std_logic_vector(   0 downto 0);
        signal cVar1S15S36N063P067P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S16S36N063P067P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S17S36N063P067P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S18S36N063P067P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S19S36N063P067P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S20S36N063P067P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S21S36N063P067P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S22S36N063P067P064P037: std_logic_vector(   0 downto 0);
        signal cVar1S23S36N063P067P064P037: std_logic_vector(   0 downto 0);
        signal cVar1S24S36N063P067P064N037: std_logic_vector(   0 downto 0);
        signal cVar1S25S36N063P067P064N037: std_logic_vector(   0 downto 0);
        signal cVar1S26S36N063N067P053P051: std_logic_vector(   0 downto 0);
        signal cVar1S27S36N063N067P053P051: std_logic_vector(   0 downto 0);
        signal cVar1S28S36N063N067P053P051: std_logic_vector(   0 downto 0);
        signal cVar1S29S36N063N067P053N051: std_logic_vector(   0 downto 0);
        signal cVar1S30S36N063N067N053P022: std_logic_vector(   0 downto 0);
        signal cVar1S31S36N063N067N053P022: std_logic_vector(   0 downto 0);
        signal cVar1S32S36N063N067N053N022: std_logic_vector(   0 downto 0);
        signal cVar1S33S36N063N067N053N022: std_logic_vector(   0 downto 0);
        signal cVar1S0S37P065P067P000P068: std_logic_vector(   0 downto 0);
        signal cVar1S1S37P065P067P000P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S37P065P067P000P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S37P065P067P000N068: std_logic_vector(   0 downto 0);
        signal cVar1S4S37P065P067P000N068: std_logic_vector(   0 downto 0);
        signal cVar1S5S37P065P067P000N068: std_logic_vector(   0 downto 0);
        signal cVar1S6S37P065P067P000P053: std_logic_vector(   0 downto 0);
        signal cVar1S7S37P065P067P062P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S37P065P067P062N056: std_logic_vector(   0 downto 0);
        signal cVar1S9S37P065P067P062N056: std_logic_vector(   0 downto 0);
        signal cVar1S10S37P065P067P062N056: std_logic_vector(   0 downto 0);
        signal cVar1S11S37P065P067P062N056: std_logic_vector(   0 downto 0);
        signal cVar1S12S37P065P067P062P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S37P065P067P062P018: std_logic_vector(   0 downto 0);
        signal cVar1S14S37P065P067P062P018: std_logic_vector(   0 downto 0);
        signal cVar1S15S37P065P067P062P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S37P065P067P062P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S37P065P060P058P069: std_logic_vector(   0 downto 0);
        signal cVar1S18S37P065P060P058N069: std_logic_vector(   0 downto 0);
        signal cVar1S19S37P065P060P058N069: std_logic_vector(   0 downto 0);
        signal cVar1S20S37P065P060P058N069: std_logic_vector(   0 downto 0);
        signal cVar1S21S37P065P060P058N069: std_logic_vector(   0 downto 0);
        signal cVar1S22S37P065P060N058P018: std_logic_vector(   0 downto 0);
        signal cVar1S23S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S24S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S25S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S26S37P065N060P062N063: std_logic_vector(   0 downto 0);
        signal cVar1S27S37P065N060P062N063: std_logic_vector(   0 downto 0);
        signal cVar1S28S37P065N060P062N063: std_logic_vector(   0 downto 0);
        signal cVar1S29S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S30S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S31S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S32S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S33S37P065N060P062P063: std_logic_vector(   0 downto 0);
        signal cVar1S0S38P019P069P015P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S38P019P069P015P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S38P019P069P015P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S38P019P069P015P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S38P019P069N015P009: std_logic_vector(   0 downto 0);
        signal cVar1S5S38P019P069N015P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S38P019P069N015N009: std_logic_vector(   0 downto 0);
        signal cVar1S7S38P019P069N015N009: std_logic_vector(   0 downto 0);
        signal cVar1S8S38P019P069N015N009: std_logic_vector(   0 downto 0);
        signal cVar1S9S38P019P069N015N009: std_logic_vector(   0 downto 0);
        signal cVar1S10S38P019N069P008P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S38P019N069P008P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S38P019N069P008P034: std_logic_vector(   0 downto 0);
        signal cVar1S13S38P019N069P008P034: std_logic_vector(   0 downto 0);
        signal cVar1S14S38P019N069P008P034: std_logic_vector(   0 downto 0);
        signal cVar1S15S38P019N069N008P016: std_logic_vector(   0 downto 0);
        signal cVar1S16S38P019N069N008P016: std_logic_vector(   0 downto 0);
        signal cVar1S17S38P019N069N008P016: std_logic_vector(   0 downto 0);
        signal cVar1S18S38P019N069N008N016: std_logic_vector(   0 downto 0);
        signal cVar1S19S38P019N069N008N016: std_logic_vector(   0 downto 0);
        signal cVar1S20S38P019N069N008N016: std_logic_vector(   0 downto 0);
        signal cVar1S21S38N019P069P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S22S38N019P069P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S23S38N019P069P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S38N019P069P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S38N019P069P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S26S38N019P069N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S27S38N019P069N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S28S38N019P069N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S29S38N019P069N033N041: std_logic_vector(   0 downto 0);
        signal cVar1S30S38N019P069N033N041: std_logic_vector(   0 downto 0);
        signal cVar1S31S38N019P069N033N041: std_logic_vector(   0 downto 0);
        signal cVar1S32S38N019P069P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S33S38N019P069P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S34S38N019P069P058P054: std_logic_vector(   0 downto 0);
        signal cVar1S35S38N019P069N058P011: std_logic_vector(   0 downto 0);
        signal cVar1S36S38N019P069N058P011: std_logic_vector(   0 downto 0);
        signal cVar1S37S38N019P069N058P011: std_logic_vector(   0 downto 0);
        signal cVar1S38S38N019P069N058P011: std_logic_vector(   0 downto 0);
        signal cVar1S0S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S5S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S6S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S7S39P011P069P058P067: std_logic_vector(   0 downto 0);
        signal cVar1S8S39P011P069P058P062: std_logic_vector(   0 downto 0);
        signal cVar1S9S39P011P069P058P062: std_logic_vector(   0 downto 0);
        signal cVar1S10S39P011P069P058P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S39P011P069P058P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S39P011P069P058P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S39P011P069P017P068: std_logic_vector(   0 downto 0);
        signal cVar1S14S39P011P069P017P068: std_logic_vector(   0 downto 0);
        signal cVar1S15S39P011P069P017P068: std_logic_vector(   0 downto 0);
        signal cVar1S16S39P011P069P017P068: std_logic_vector(   0 downto 0);
        signal cVar1S17S39P011P069P017N068: std_logic_vector(   0 downto 0);
        signal cVar1S18S39P011P069P017N068: std_logic_vector(   0 downto 0);
        signal cVar1S19S39P011P069N017P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S39P011P069N017N047: std_logic_vector(   0 downto 0);
        signal cVar1S21S39P011P069N017N047: std_logic_vector(   0 downto 0);
        signal cVar1S22S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S23S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S24S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S25S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S26S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S27S39P011P019P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S28S39P011P019N062P064: std_logic_vector(   0 downto 0);
        signal cVar1S29S39P011P019N062P064: std_logic_vector(   0 downto 0);
        signal cVar1S30S39P011P019N062P064: std_logic_vector(   0 downto 0);
        signal cVar1S31S39P011P019N062P064: std_logic_vector(   0 downto 0);
        signal cVar1S32S39P011N019P060P061: std_logic_vector(   0 downto 0);
        signal cVar1S33S39P011N019P060P061: std_logic_vector(   0 downto 0);
        signal cVar1S34S39P011N019P060P061: std_logic_vector(   0 downto 0);
        signal cVar1S35S39P011N019P060N061: std_logic_vector(   0 downto 0);
        signal cVar1S36S39P011N019P060N061: std_logic_vector(   0 downto 0);
        signal cVar1S37S39P011N019N060P049: std_logic_vector(   0 downto 0);
        signal cVar1S38S39P011N019N060P049: std_logic_vector(   0 downto 0);
        signal cVar1S39S39P011N019N060N049: std_logic_vector(   0 downto 0);
        signal cVar1S40S39P011N019N060N049: std_logic_vector(   0 downto 0);
        signal cVar1S0S40P069P053P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S1S40P069P053P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S2S40P069P053P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S40P069P053P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S40P069P053P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S5S40P069P053N067P064: std_logic_vector(   0 downto 0);
        signal cVar1S6S40P069P053N067P064: std_logic_vector(   0 downto 0);
        signal cVar1S7S40P069P053N067P064: std_logic_vector(   0 downto 0);
        signal cVar1S8S40P069P053N067N064: std_logic_vector(   0 downto 0);
        signal cVar1S9S40P069P053N067N064: std_logic_vector(   0 downto 0);
        signal cVar1S10S40P069P053N067N064: std_logic_vector(   0 downto 0);
        signal cVar1S11S40P069P053N067N064: std_logic_vector(   0 downto 0);
        signal cVar1S12S40P069P053P059P060nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S40P069P053P059N060: std_logic_vector(   0 downto 0);
        signal cVar1S14S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S15S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S19S40N069P031P013P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S40N069P031N013P058: std_logic_vector(   0 downto 0);
        signal cVar1S21S40N069P031N013P058: std_logic_vector(   0 downto 0);
        signal cVar1S22S40N069P031N013N058: std_logic_vector(   0 downto 0);
        signal cVar1S23S40N069P031N013N058: std_logic_vector(   0 downto 0);
        signal cVar1S24S40N069P031N013N058: std_logic_vector(   0 downto 0);
        signal cVar1S25S40N069N031P030P061: std_logic_vector(   0 downto 0);
        signal cVar1S26S40N069N031P030P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S40N069N031P030N061: std_logic_vector(   0 downto 0);
        signal cVar1S28S40N069N031P030N061: std_logic_vector(   0 downto 0);
        signal cVar1S29S40N069N031P030N061: std_logic_vector(   0 downto 0);
        signal cVar1S30S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S31S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S32S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S33S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S34S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S35S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S36S40N069N031N030P000: std_logic_vector(   0 downto 0);
        signal cVar1S0S41P025P004P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S41P025P004N048P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S41P025N004P007P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S41P025N004P007P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S41P025N004P007P067: std_logic_vector(   0 downto 0);
        signal cVar1S5S41P025N004N007P037: std_logic_vector(   0 downto 0);
        signal cVar1S6S41P025N004N007P037: std_logic_vector(   0 downto 0);
        signal cVar1S7S41P025N004N007N037: std_logic_vector(   0 downto 0);
        signal cVar1S8S41P025N004N007N037: std_logic_vector(   0 downto 0);
        signal cVar1S9S41P025N004N007N037: std_logic_vector(   0 downto 0);
        signal cVar1S10S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S11S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S12S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S13S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S14S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S15S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S41N025P062P058P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S41N025P062P058P049: std_logic_vector(   0 downto 0);
        signal cVar1S18S41N025P062P058P049: std_logic_vector(   0 downto 0);
        signal cVar1S19S41N025N062P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S20S41N025N062P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S41N025N062P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S41N025N062P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S23S41N025N062P027P026: std_logic_vector(   0 downto 0);
        signal cVar1S24S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S25S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S26S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S27S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S28S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S29S41N025N062N027P048: std_logic_vector(   0 downto 0);
        signal cVar1S0S42P068P004P025P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S42P068P004P025N048: std_logic_vector(   0 downto 0);
        signal cVar1S2S42P068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S3S42P068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S4S42P068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S5S42P068P004N025N040: std_logic_vector(   0 downto 0);
        signal cVar1S6S42P068P004N025N040: std_logic_vector(   0 downto 0);
        signal cVar1S7S42P068N004P055P013: std_logic_vector(   0 downto 0);
        signal cVar1S8S42P068N004P055P013: std_logic_vector(   0 downto 0);
        signal cVar1S9S42P068N004P055P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S42P068N004P055P013: std_logic_vector(   0 downto 0);
        signal cVar1S11S42P068N004P055P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S42P068N004P055P066: std_logic_vector(   0 downto 0);
        signal cVar1S13S42P068N004P055P066: std_logic_vector(   0 downto 0);
        signal cVar1S14S42P068N004P055P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S42P068N004P055P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S42P068N004P055P066: std_logic_vector(   0 downto 0);
        signal cVar1S17S42P068P015P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S18S42P068P015P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S19S42P068P015P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S20S42P068P015P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S21S42P068P015P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S42P068P015N061P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S42P068P015N061N025: std_logic_vector(   0 downto 0);
        signal cVar1S24S42P068P015N061N025: std_logic_vector(   0 downto 0);
        signal cVar1S25S42P068P015N061N025: std_logic_vector(   0 downto 0);
        signal cVar1S26S42P068N015P059P069: std_logic_vector(   0 downto 0);
        signal cVar1S27S42P068N015P059P069: std_logic_vector(   0 downto 0);
        signal cVar1S28S42P068N015P059P069: std_logic_vector(   0 downto 0);
        signal cVar1S29S42P068N015P059P069: std_logic_vector(   0 downto 0);
        signal cVar1S30S42P068N015P059P069: std_logic_vector(   0 downto 0);
        signal cVar1S31S42P068N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S32S42P068N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S33S42P068N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S34S42P068N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S35S42P068N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S36S42P068N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S1S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S2S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S3S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S4S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S5S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S43P068P069P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S7S43P068P069P000P064: std_logic_vector(   0 downto 0);
        signal cVar1S8S43P068P069P000N064: std_logic_vector(   0 downto 0);
        signal cVar1S9S43P068P069P000N064: std_logic_vector(   0 downto 0);
        signal cVar1S10S43P068P069P023P019: std_logic_vector(   0 downto 0);
        signal cVar1S11S43P068P069P023P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S43P068P069P023P019: std_logic_vector(   0 downto 0);
        signal cVar1S13S43P068P069P023P019: std_logic_vector(   0 downto 0);
        signal cVar1S14S43P068P069P023P019: std_logic_vector(   0 downto 0);
        signal cVar1S15S43N068P004P025P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S43N068P004P025N048: std_logic_vector(   0 downto 0);
        signal cVar1S17S43N068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S18S43N068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S19S43N068P004N025P040: std_logic_vector(   0 downto 0);
        signal cVar1S20S43N068P004N025N040: std_logic_vector(   0 downto 0);
        signal cVar1S21S43N068P004N025N040: std_logic_vector(   0 downto 0);
        signal cVar1S22S43N068P004N025N040: std_logic_vector(   0 downto 0);
        signal cVar1S23S43N068N004P013P064: std_logic_vector(   0 downto 0);
        signal cVar1S24S43N068N004P013P064: std_logic_vector(   0 downto 0);
        signal cVar1S25S43N068N004P013N064: std_logic_vector(   0 downto 0);
        signal cVar1S26S43N068N004P013N064: std_logic_vector(   0 downto 0);
        signal cVar1S27S43N068N004P013N064: std_logic_vector(   0 downto 0);
        signal cVar1S28S43N068N004N013P032: std_logic_vector(   0 downto 0);
        signal cVar1S29S43N068N004N013P032: std_logic_vector(   0 downto 0);
        signal cVar1S30S43N068N004N013P032: std_logic_vector(   0 downto 0);
        signal cVar1S31S43N068N004N013P032: std_logic_vector(   0 downto 0);
        signal cVar1S32S43N068N004N013N032: std_logic_vector(   0 downto 0);
        signal cVar1S33S43N068N004N013N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S44P068P001P018P065: std_logic_vector(   0 downto 0);
        signal cVar1S1S44P068P001P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S2S44P068P001P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S3S44P068P001P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S4S44P068P001P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S5S44P068P001N018P046: std_logic_vector(   0 downto 0);
        signal cVar1S6S44P068P001N018P046: std_logic_vector(   0 downto 0);
        signal cVar1S7S44P068P001N018N046: std_logic_vector(   0 downto 0);
        signal cVar1S8S44P068P001N018N046: std_logic_vector(   0 downto 0);
        signal cVar1S9S44P068P001N018N046: std_logic_vector(   0 downto 0);
        signal cVar1S10S44P068P001N018N046: std_logic_vector(   0 downto 0);
        signal cVar1S11S44P068P001P054P036: std_logic_vector(   0 downto 0);
        signal cVar1S12S44P068P001P054P036: std_logic_vector(   0 downto 0);
        signal cVar1S13S44P068P001P054P036: std_logic_vector(   0 downto 0);
        signal cVar1S14S44P068P001P054P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S44P068P067P057P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S44P068P067P057P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S44P068P067P057N032: std_logic_vector(   0 downto 0);
        signal cVar1S18S44P068P067P057N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S44P068N067P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S20S44P068N067P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S21S44P068N067P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S22S44P068N067P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S44P068N067N025P066: std_logic_vector(   0 downto 0);
        signal cVar1S24S44P068N067N025N066: std_logic_vector(   0 downto 0);
        signal cVar1S25S44P068N067N025N066: std_logic_vector(   0 downto 0);
        signal cVar1S0S45P014P068P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S45P014P068P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S45P014P068P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S45P014P068P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S45P014P068P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S5S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S6S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S9S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S10S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S11S45P014P068N016P036: std_logic_vector(   0 downto 0);
        signal cVar1S12S45P014P068P067P045: std_logic_vector(   0 downto 0);
        signal cVar1S13S45P014P068P067P045: std_logic_vector(   0 downto 0);
        signal cVar1S14S45P014P068P067N045: std_logic_vector(   0 downto 0);
        signal cVar1S15S45P014P068P067N045: std_logic_vector(   0 downto 0);
        signal cVar1S16S45P014P068P067N045: std_logic_vector(   0 downto 0);
        signal cVar1S17S45P014P068P067P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S45P014P068P067P035: std_logic_vector(   0 downto 0);
        signal cVar1S19S45P014P015P021P034: std_logic_vector(   0 downto 0);
        signal cVar1S20S45P014P015P021P034: std_logic_vector(   0 downto 0);
        signal cVar1S21S45P014P015P021N034: std_logic_vector(   0 downto 0);
        signal cVar1S22S45P014P015P021N034: std_logic_vector(   0 downto 0);
        signal cVar1S23S45P014P015P021N034: std_logic_vector(   0 downto 0);
        signal cVar1S24S45P014P015P021P037: std_logic_vector(   0 downto 0);
        signal cVar1S25S45P014P015P021N037: std_logic_vector(   0 downto 0);
        signal cVar1S26S45P014P015P018P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S45P014P015P018P061: std_logic_vector(   0 downto 0);
        signal cVar1S28S45P014P015P018N061: std_logic_vector(   0 downto 0);
        signal cVar1S29S45P014P015P018N061: std_logic_vector(   0 downto 0);
        signal cVar1S30S45P014P015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S0S46P016P038P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S46P016P038N021P019: std_logic_vector(   0 downto 0);
        signal cVar1S2S46P016P038N021P019: std_logic_vector(   0 downto 0);
        signal cVar1S3S46P016P038N021P019: std_logic_vector(   0 downto 0);
        signal cVar1S4S46P016P038N021P019: std_logic_vector(   0 downto 0);
        signal cVar1S5S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S6S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S9S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S10S46P016N038P010P036: std_logic_vector(   0 downto 0);
        signal cVar1S11S46P016N038N010P008: std_logic_vector(   0 downto 0);
        signal cVar1S12S46P016N038N010P008: std_logic_vector(   0 downto 0);
        signal cVar1S13S46P016N038N010P008: std_logic_vector(   0 downto 0);
        signal cVar1S14S46P016N038N010N008: std_logic_vector(   0 downto 0);
        signal cVar1S15S46P016N038N010N008: std_logic_vector(   0 downto 0);
        signal cVar1S16S46P016N038N010N008: std_logic_vector(   0 downto 0);
        signal cVar1S17S46P016P032P049P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S46P016P032P049P056: std_logic_vector(   0 downto 0);
        signal cVar1S19S46P016P032P049P056: std_logic_vector(   0 downto 0);
        signal cVar1S20S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S21S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S22S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S23S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S24S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S25S46P016N032P018P035: std_logic_vector(   0 downto 0);
        signal cVar1S26S46P016N032P018P058: std_logic_vector(   0 downto 0);
        signal cVar1S27S46P016N032P018P058: std_logic_vector(   0 downto 0);
        signal cVar1S28S46P016N032P018P058: std_logic_vector(   0 downto 0);
        signal cVar1S29S46P016N032P018N058: std_logic_vector(   0 downto 0);
        signal cVar1S30S46P016N032P018N058: std_logic_vector(   0 downto 0);
        signal cVar1S31S46P016N032P018N058: std_logic_vector(   0 downto 0);
        signal cVar1S32S46P016N032P018N058: std_logic_vector(   0 downto 0);
        signal cVar1S0S47P067P016P064P047: std_logic_vector(   0 downto 0);
        signal cVar1S1S47P067P016P064P047: std_logic_vector(   0 downto 0);
        signal cVar1S2S47P067P016P064P047: std_logic_vector(   0 downto 0);
        signal cVar1S3S47P067P016P064N047: std_logic_vector(   0 downto 0);
        signal cVar1S4S47P067P016P064N047: std_logic_vector(   0 downto 0);
        signal cVar1S5S47P067P016P064N047: std_logic_vector(   0 downto 0);
        signal cVar1S6S47P067P016P064N047: std_logic_vector(   0 downto 0);
        signal cVar1S7S47P067P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S8S47P067P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S47P067P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S47P067P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S11S47P067P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S12S47P067P016P002P006: std_logic_vector(   0 downto 0);
        signal cVar1S13S47P067P016P002P006: std_logic_vector(   0 downto 0);
        signal cVar1S14S47P067P016P002P006: std_logic_vector(   0 downto 0);
        signal cVar1S15S47P067P016P002P006: std_logic_vector(   0 downto 0);
        signal cVar1S16S47P067P016P002P006: std_logic_vector(   0 downto 0);
        signal cVar1S17S47P067P016P002P050: std_logic_vector(   0 downto 0);
        signal cVar1S18S47P067P016P002P050: std_logic_vector(   0 downto 0);
        signal cVar1S19S47P067P062P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S20S47P067P062P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S21S47P067P062P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S22S47P067P062P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S23S47P067P062P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S24S47P067P062P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S25S47P067P062N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S26S47P067P062N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S27S47P067P062N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S28S47P067P062N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S29S47P067P062N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S30S47P067P062P044P035: std_logic_vector(   0 downto 0);
        signal cVar1S31S47P067P062P044P035: std_logic_vector(   0 downto 0);
        signal cVar1S32S47P067P062P044N035: std_logic_vector(   0 downto 0);
        signal cVar1S33S47P067P062P044N035: std_logic_vector(   0 downto 0);
        signal cVar1S0S48P067P062P057P049: std_logic_vector(   0 downto 0);
        signal cVar1S1S48P067P062P057P049: std_logic_vector(   0 downto 0);
        signal cVar1S2S48P067P062P057N049: std_logic_vector(   0 downto 0);
        signal cVar1S3S48P067P062P057N049: std_logic_vector(   0 downto 0);
        signal cVar1S4S48P067P062P057N049: std_logic_vector(   0 downto 0);
        signal cVar1S5S48P067P062P057P051: std_logic_vector(   0 downto 0);
        signal cVar1S6S48P067P062P057P051: std_logic_vector(   0 downto 0);
        signal cVar1S7S48P067P062P057P051: std_logic_vector(   0 downto 0);
        signal cVar1S8S48P067P062P057P051: std_logic_vector(   0 downto 0);
        signal cVar1S9S48P067P062P044P042: std_logic_vector(   0 downto 0);
        signal cVar1S10S48N067P036P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S48N067P036P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S12S48N067P036P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S13S48N067P036P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S14S48N067P036P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S15S48N067P036N027P016: std_logic_vector(   0 downto 0);
        signal cVar1S16S48N067P036N027P016: std_logic_vector(   0 downto 0);
        signal cVar1S17S48N067P036N027P016: std_logic_vector(   0 downto 0);
        signal cVar1S18S48N067P036N027N016: std_logic_vector(   0 downto 0);
        signal cVar1S19S48N067P036N027N016: std_logic_vector(   0 downto 0);
        signal cVar1S20S48N067P036N027N016: std_logic_vector(   0 downto 0);
        signal cVar1S21S48N067P036N027N016: std_logic_vector(   0 downto 0);
        signal cVar1S22S48N067P036P005P043: std_logic_vector(   0 downto 0);
        signal cVar1S23S48N067P036P005P043: std_logic_vector(   0 downto 0);
        signal cVar1S24S48N067P036P005N043: std_logic_vector(   0 downto 0);
        signal cVar1S25S48N067P036P005P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S48N067P036P005N032: std_logic_vector(   0 downto 0);
        signal cVar1S27S48N067P036P005N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S1S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S49P036P011P010P013: std_logic_vector(   0 downto 0);
        signal cVar1S6S49P036P011P010P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S49P036P011P010N042: std_logic_vector(   0 downto 0);
        signal cVar1S8S49P036P011P010N042: std_logic_vector(   0 downto 0);
        signal cVar1S9S49P036N011P005P039: std_logic_vector(   0 downto 0);
        signal cVar1S10S49P036N011P005P039: std_logic_vector(   0 downto 0);
        signal cVar1S11S49P036N011P005P039: std_logic_vector(   0 downto 0);
        signal cVar1S12S49P036N011P005N039: std_logic_vector(   0 downto 0);
        signal cVar1S13S49P036N011P005N039: std_logic_vector(   0 downto 0);
        signal cVar1S14S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S15S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S16S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S17S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S18S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S19S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S20S49P036N011N005P016: std_logic_vector(   0 downto 0);
        signal cVar1S21S49P036P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S49P036P043N022P015: std_logic_vector(   0 downto 0);
        signal cVar1S23S49P036P043N022P015: std_logic_vector(   0 downto 0);
        signal cVar1S24S49P036P043N022P015: std_logic_vector(   0 downto 0);
        signal cVar1S25S49P036N043P045P016: std_logic_vector(   0 downto 0);
        signal cVar1S26S49P036N043P045P016: std_logic_vector(   0 downto 0);
        signal cVar1S27S49P036N043P045N016: std_logic_vector(   0 downto 0);
        signal cVar1S28S49P036N043P045N016: std_logic_vector(   0 downto 0);
        signal cVar1S29S49P036N043P045N016: std_logic_vector(   0 downto 0);
        signal cVar1S30S49P036N043P045P016: std_logic_vector(   0 downto 0);
        signal cVar1S0S50P036P033P015P038: std_logic_vector(   0 downto 0);
        signal cVar1S1S50P036P033P015P038: std_logic_vector(   0 downto 0);
        signal cVar1S2S50P036P033P015P038: std_logic_vector(   0 downto 0);
        signal cVar1S3S50P036P033P015N038: std_logic_vector(   0 downto 0);
        signal cVar1S4S50P036P033P015N038: std_logic_vector(   0 downto 0);
        signal cVar1S5S50P036P033P015N038: std_logic_vector(   0 downto 0);
        signal cVar1S6S50P036P033P015N038: std_logic_vector(   0 downto 0);
        signal cVar1S7S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S8S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S9S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S10S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S11S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S12S50P036P033P015P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S50P036P033P026P001: std_logic_vector(   0 downto 0);
        signal cVar1S14S50P036P033P026P001: std_logic_vector(   0 downto 0);
        signal cVar1S15S50P036P033P026P001: std_logic_vector(   0 downto 0);
        signal cVar1S16S50P036P033P026P001: std_logic_vector(   0 downto 0);
        signal cVar1S17S50P036P033P026P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S50P036P033P026N047: std_logic_vector(   0 downto 0);
        signal cVar1S19S50P036P068P065P018: std_logic_vector(   0 downto 0);
        signal cVar1S20S50P036P068P065N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S50P036P068P065N018: std_logic_vector(   0 downto 0);
        signal cVar1S22S50P036P068P065N018: std_logic_vector(   0 downto 0);
        signal cVar1S23S50P036P068N065P018: std_logic_vector(   0 downto 0);
        signal cVar1S24S50P036P068N065P018: std_logic_vector(   0 downto 0);
        signal cVar1S25S50P036P068N065P018: std_logic_vector(   0 downto 0);
        signal cVar1S26S50P036P068N065P018: std_logic_vector(   0 downto 0);
        signal cVar1S27S50P036P068P019P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S50P036P068P019N025: std_logic_vector(   0 downto 0);
        signal cVar1S29S50P036P068P019N025: std_logic_vector(   0 downto 0);
        signal cVar1S30S50P036P068N019P066: std_logic_vector(   0 downto 0);
        signal cVar1S31S50P036P068N019P066: std_logic_vector(   0 downto 0);
        signal cVar1S32S50P036P068N019P066: std_logic_vector(   0 downto 0);
        signal cVar1S33S50P036P068N019P066: std_logic_vector(   0 downto 0);
        signal cVar1S34S50P036P068N019N066: std_logic_vector(   0 downto 0);
        signal cVar1S0S51P033P015P032P035: std_logic_vector(   0 downto 0);
        signal cVar1S1S51P033P015P032P035: std_logic_vector(   0 downto 0);
        signal cVar1S2S51P033P015P032P035: std_logic_vector(   0 downto 0);
        signal cVar1S3S51P033P015P032P035: std_logic_vector(   0 downto 0);
        signal cVar1S4S51P033P015P032P035: std_logic_vector(   0 downto 0);
        signal cVar1S5S51P033P015N032P017: std_logic_vector(   0 downto 0);
        signal cVar1S6S51P033P015N032P017: std_logic_vector(   0 downto 0);
        signal cVar1S7S51P033P015N032P017: std_logic_vector(   0 downto 0);
        signal cVar1S8S51P033P015N032P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S51P033P015N032P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S51P033N015P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S11S51P033N015P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S12S51P033N015P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S51P033N015P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S14S51P033N015P059N049: std_logic_vector(   0 downto 0);
        signal cVar1S15S51P033N015P059N049: std_logic_vector(   0 downto 0);
        signal cVar1S16S51P033N015P059N049: std_logic_vector(   0 downto 0);
        signal cVar1S17S51P033N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S51P033N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S19S51P033N015P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S20S51P033N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S21S51P033N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S22S51P033N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S23S51P033N015P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S24S51P033P056P016P060: std_logic_vector(   0 downto 0);
        signal cVar1S25S51P033P056P016P060: std_logic_vector(   0 downto 0);
        signal cVar1S26S51P033P056P016P060: std_logic_vector(   0 downto 0);
        signal cVar1S27S51P033P056P016P060: std_logic_vector(   0 downto 0);
        signal cVar1S28S51P033P056P016P058: std_logic_vector(   0 downto 0);
        signal cVar1S29S51P033N056P006P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S51P033N056P006N042: std_logic_vector(   0 downto 0);
        signal cVar1S31S51P033N056P006N042: std_logic_vector(   0 downto 0);
        signal cVar1S0S52P006P017P064P037: std_logic_vector(   0 downto 0);
        signal cVar1S1S52P006P017P064P037: std_logic_vector(   0 downto 0);
        signal cVar1S2S52P006P017P064N037: std_logic_vector(   0 downto 0);
        signal cVar1S3S52P006P017P064N037: std_logic_vector(   0 downto 0);
        signal cVar1S4S52P006P017P064N037: std_logic_vector(   0 downto 0);
        signal cVar1S5S52P006P017N064P005: std_logic_vector(   0 downto 0);
        signal cVar1S6S52P006P017N064P005: std_logic_vector(   0 downto 0);
        signal cVar1S7S52P006P017N064P005: std_logic_vector(   0 downto 0);
        signal cVar1S8S52P006P017N064P005: std_logic_vector(   0 downto 0);
        signal cVar1S9S52P006P017N064P005: std_logic_vector(   0 downto 0);
        signal cVar1S10S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S11S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S12S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S13S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S14S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S15S52P006N017P059P044: std_logic_vector(   0 downto 0);
        signal cVar1S16S52P006N017P059P060: std_logic_vector(   0 downto 0);
        signal cVar1S17S52P006N017P059P060: std_logic_vector(   0 downto 0);
        signal cVar1S18S52P006N017P059P060: std_logic_vector(   0 downto 0);
        signal cVar1S19S52P006N017P059P060: std_logic_vector(   0 downto 0);
        signal cVar1S20S52P006P042P044nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S52P006P042N044P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S52P006N042P047P064: std_logic_vector(   0 downto 0);
        signal cVar1S23S52P006N042P047P064: std_logic_vector(   0 downto 0);
        signal cVar1S24S52P006N042P047P064: std_logic_vector(   0 downto 0);
        signal cVar1S25S52P006N042N047P043: std_logic_vector(   0 downto 0);
        signal cVar1S26S52P006N042N047N043: std_logic_vector(   0 downto 0);
        signal cVar1S27S52P006N042N047N043: std_logic_vector(   0 downto 0);
        signal cVar1S0S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S1S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S2S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S3S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S4S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S5S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S6S53P016P059P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S8S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S9S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S10S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S12S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S13S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S14S53P016P059P017P015: std_logic_vector(   0 downto 0);
        signal cVar1S15S53P016P059P015P019: std_logic_vector(   0 downto 0);
        signal cVar1S16S53P016P059P015P019: std_logic_vector(   0 downto 0);
        signal cVar1S17S53P016P059P015P019: std_logic_vector(   0 downto 0);
        signal cVar1S18S53P016P059P015N019: std_logic_vector(   0 downto 0);
        signal cVar1S19S53P016P059P015N019: std_logic_vector(   0 downto 0);
        signal cVar1S20S53P016P059P015N019: std_logic_vector(   0 downto 0);
        signal cVar1S21S53P016P059N015P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S53P016P059N015P066: std_logic_vector(   0 downto 0);
        signal cVar1S23S53P016P059N015P066: std_logic_vector(   0 downto 0);
        signal cVar1S24S53P016P059N015P066: std_logic_vector(   0 downto 0);
        signal cVar1S25S53P016P059N015P066: std_logic_vector(   0 downto 0);
        signal cVar1S26S53P016P038P002P021: std_logic_vector(   0 downto 0);
        signal cVar1S27S53P016P038P002P021: std_logic_vector(   0 downto 0);
        signal cVar1S28S53P016P038P002P021: std_logic_vector(   0 downto 0);
        signal cVar1S29S53P016P038P002P021: std_logic_vector(   0 downto 0);
        signal cVar1S30S53P016P038P002P021: std_logic_vector(   0 downto 0);
        signal cVar1S31S53P016P038P002P019: std_logic_vector(   0 downto 0);
        signal cVar1S32S53P016P038P002P019: std_logic_vector(   0 downto 0);
        signal cVar1S33S53P016P038P002N019: std_logic_vector(   0 downto 0);
        signal cVar1S34S53P016P038P002N019: std_logic_vector(   0 downto 0);
        signal cVar1S35S53P016P038P033P064: std_logic_vector(   0 downto 0);
        signal cVar1S36S53P016P038P033P064: std_logic_vector(   0 downto 0);
        signal cVar1S37S53P016P038P033P064: std_logic_vector(   0 downto 0);
        signal cVar1S0S54P037P016P038P002: std_logic_vector(   0 downto 0);
        signal cVar1S1S54P037P016P038P002: std_logic_vector(   0 downto 0);
        signal cVar1S2S54P037P016P038P002: std_logic_vector(   0 downto 0);
        signal cVar1S3S54P037P016P038P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S54P037P016P038P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S54P037P016P038P033: std_logic_vector(   0 downto 0);
        signal cVar1S6S54P037P016P038P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S54P037N016P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S8S54P037N016P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S9S54P037N016P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S10S54P037N016N050P039: std_logic_vector(   0 downto 0);
        signal cVar1S11S54P037N016N050P039: std_logic_vector(   0 downto 0);
        signal cVar1S12S54P037N016N050P039: std_logic_vector(   0 downto 0);
        signal cVar1S13S54P037N016N050N039: std_logic_vector(   0 downto 0);
        signal cVar1S14S54P037N016N050N039: std_logic_vector(   0 downto 0);
        signal cVar1S15S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S16S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S17S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S18S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S19S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S20S54P037P018P060P031: std_logic_vector(   0 downto 0);
        signal cVar1S21S54P037P018P060P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S54P037P018P060P066: std_logic_vector(   0 downto 0);
        signal cVar1S23S54P037P018P060P066: std_logic_vector(   0 downto 0);
        signal cVar1S24S54P037P018P060N066: std_logic_vector(   0 downto 0);
        signal cVar1S25S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S26S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S27S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S28S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S29S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S30S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S31S54P037N018P017P065: std_logic_vector(   0 downto 0);
        signal cVar1S32S54P037N018N017P064: std_logic_vector(   0 downto 0);
        signal cVar1S33S54P037N018N017P064: std_logic_vector(   0 downto 0);
        signal cVar1S34S54P037N018N017P064: std_logic_vector(   0 downto 0);
        signal cVar1S35S54P037N018N017P064: std_logic_vector(   0 downto 0);
        signal cVar1S0S55P016P037P062P001: std_logic_vector(   0 downto 0);
        signal cVar1S1S55P016P037P062P001: std_logic_vector(   0 downto 0);
        signal cVar1S2S55P016P037P062P001: std_logic_vector(   0 downto 0);
        signal cVar1S3S55P016P037P062P001: std_logic_vector(   0 downto 0);
        signal cVar1S4S55P016P037P062P001: std_logic_vector(   0 downto 0);
        signal cVar1S5S55P016P037P062P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S55P016P037P062P047: std_logic_vector(   0 downto 0);
        signal cVar1S7S55P016P037P062P047: std_logic_vector(   0 downto 0);
        signal cVar1S8S55P016P037P017P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S55P016P037P017N008: std_logic_vector(   0 downto 0);
        signal cVar1S10S55P016P037P017N008: std_logic_vector(   0 downto 0);
        signal cVar1S11S55P016P037P017N008: std_logic_vector(   0 downto 0);
        signal cVar1S12S55P016P037P017N008: std_logic_vector(   0 downto 0);
        signal cVar1S13S55P016P037N017P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S55P016P037N017P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S55P016P037N017N067: std_logic_vector(   0 downto 0);
        signal cVar1S16S55P016P037N017N067: std_logic_vector(   0 downto 0);
        signal cVar1S17S55P016P037N017N067: std_logic_vector(   0 downto 0);
        signal cVar1S18S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S19S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S20S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S23S55P016P036P038P037: std_logic_vector(   0 downto 0);
        signal cVar1S24S55P016N036P046P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S55P016N036P046N024: std_logic_vector(   0 downto 0);
        signal cVar1S26S55P016N036P046N024: std_logic_vector(   0 downto 0);
        signal cVar1S27S55P016N036N046P025: std_logic_vector(   0 downto 0);
        signal cVar1S28S55P016N036N046P025: std_logic_vector(   0 downto 0);
        signal cVar1S29S55P016N036N046P025: std_logic_vector(   0 downto 0);
        signal cVar1S30S55P016N036N046P025: std_logic_vector(   0 downto 0);
        signal cVar1S31S55P016N036N046P025: std_logic_vector(   0 downto 0);
        signal cVar1S0S56P016P036P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S1S56P016P036P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S2S56P016P036P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S56P016P036P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S4S56P016P036P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S5S56P016P036P054P052: std_logic_vector(   0 downto 0);
        signal cVar1S6S56P016P036P054P052: std_logic_vector(   0 downto 0);
        signal cVar1S7S56P016P036P054P052: std_logic_vector(   0 downto 0);
        signal cVar1S8S56P016P036P054P052: std_logic_vector(   0 downto 0);
        signal cVar1S9S56P016P036P054P052: std_logic_vector(   0 downto 0);
        signal cVar1S10S56P016P036P043P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S56P016P036N043P005: std_logic_vector(   0 downto 0);
        signal cVar1S12S56P016P036N043P005: std_logic_vector(   0 downto 0);
        signal cVar1S13S56P016P036N043P005: std_logic_vector(   0 downto 0);
        signal cVar1S14S56N016P053P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S15S56N016P053P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S16S56N016P053P051N057: std_logic_vector(   0 downto 0);
        signal cVar1S17S56N016P053P051N057: std_logic_vector(   0 downto 0);
        signal cVar1S18S56N016P053P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S19S56N016P053P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S20S56N016P053P028P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S56N016P053P028P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S56N016P053P028P066: std_logic_vector(   0 downto 0);
        signal cVar1S23S56N016P053P028P066: std_logic_vector(   0 downto 0);
        signal cVar1S24S56N016P053P028P066: std_logic_vector(   0 downto 0);
        signal cVar1S25S56N016P053N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S26S56N016P053N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S27S56N016P053N028P066: std_logic_vector(   0 downto 0);
        signal cVar1S28S56N016P053N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S29S56N016P053N028N066: std_logic_vector(   0 downto 0);
        signal cVar1S0S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S1S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S2S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S3S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S4S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S5S57P056P051P016P053: std_logic_vector(   0 downto 0);
        signal cVar1S6S57P056P051P016P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S57P056P051P016P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S57P056P051P016P036: std_logic_vector(   0 downto 0);
        signal cVar1S9S57P056P051P016N036: std_logic_vector(   0 downto 0);
        signal cVar1S10S57P056P051P016N036: std_logic_vector(   0 downto 0);
        signal cVar1S11S57P056P051P016N036: std_logic_vector(   0 downto 0);
        signal cVar1S12S57P056P051P016N036: std_logic_vector(   0 downto 0);
        signal cVar1S13S57P056P051P008P036: std_logic_vector(   0 downto 0);
        signal cVar1S14S57P056P051P008P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S57P056P051P008N036: std_logic_vector(   0 downto 0);
        signal cVar1S16S57P056P051P008N036: std_logic_vector(   0 downto 0);
        signal cVar1S17S57P056P051P008N036: std_logic_vector(   0 downto 0);
        signal cVar1S18S57P056P051N008P064: std_logic_vector(   0 downto 0);
        signal cVar1S19S57P056P051N008P064: std_logic_vector(   0 downto 0);
        signal cVar1S20S57P056P051N008P064: std_logic_vector(   0 downto 0);
        signal cVar1S21S57P056P051N008P064: std_logic_vector(   0 downto 0);
        signal cVar1S22S57P056P052P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S23S57P056P052P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S24S57P056P052P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S25S57P056P052P027P050: std_logic_vector(   0 downto 0);
        signal cVar1S26S57P056P052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S27S57P056P052N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S57P056P052N009N008: std_logic_vector(   0 downto 0);
        signal cVar1S0S58P017P065P041P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S58P017P065P041P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S58P017P065P041P062: std_logic_vector(   0 downto 0);
        signal cVar1S3S58P017P065P041P062: std_logic_vector(   0 downto 0);
        signal cVar1S4S58P017P065N041P038: std_logic_vector(   0 downto 0);
        signal cVar1S5S58P017P065N041P038: std_logic_vector(   0 downto 0);
        signal cVar1S6S58P017P065N041N038: std_logic_vector(   0 downto 0);
        signal cVar1S7S58P017P065N041N038: std_logic_vector(   0 downto 0);
        signal cVar1S8S58P017P065N041N038: std_logic_vector(   0 downto 0);
        signal cVar1S9S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S11S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S12S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S13S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S14S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S15S58P017P065P063P056: std_logic_vector(   0 downto 0);
        signal cVar1S16S58P017P065N063P000: std_logic_vector(   0 downto 0);
        signal cVar1S17S58P017P065N063N000: std_logic_vector(   0 downto 0);
        signal cVar1S18S58P017P065N063N000: std_logic_vector(   0 downto 0);
        signal cVar1S19S58P017P065N063N000: std_logic_vector(   0 downto 0);
        signal cVar1S20S58P017P064P037P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S58P017P064P037P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S58P017P064P037P026: std_logic_vector(   0 downto 0);
        signal cVar1S23S58P017P064P037P026: std_logic_vector(   0 downto 0);
        signal cVar1S24S58P017P064N037P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S58P017P064N037P003: std_logic_vector(   0 downto 0);
        signal cVar1S26S58P017P064N037P003: std_logic_vector(   0 downto 0);
        signal cVar1S27S58P017P064N037N003: std_logic_vector(   0 downto 0);
        signal cVar1S28S58P017N064P063P068: std_logic_vector(   0 downto 0);
        signal cVar1S29S58P017N064P063P068: std_logic_vector(   0 downto 0);
        signal cVar1S30S58P017N064P063P068: std_logic_vector(   0 downto 0);
        signal cVar1S31S58P017N064P063P068: std_logic_vector(   0 downto 0);
        signal cVar1S32S58P017N064P063P068: std_logic_vector(   0 downto 0);
        signal cVar1S33S58P017N064N063P036: std_logic_vector(   0 downto 0);
        signal cVar1S34S58P017N064N063P036: std_logic_vector(   0 downto 0);
        signal cVar1S35S58P017N064N063N036: std_logic_vector(   0 downto 0);
        signal cVar1S36S58P017N064N063N036: std_logic_vector(   0 downto 0);
        signal cVar1S37S58P017N064N063N036: std_logic_vector(   0 downto 0);
        signal cVar1S0S59P063P001P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S1S59P063P001P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S2S59P063P001P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S3S59P063P001P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S4S59P063P001P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S5S59P063P001N035P057: std_logic_vector(   0 downto 0);
        signal cVar1S6S59P063P001N035P057: std_logic_vector(   0 downto 0);
        signal cVar1S7S59P063P001N035P057: std_logic_vector(   0 downto 0);
        signal cVar1S8S59P063P001N035P057: std_logic_vector(   0 downto 0);
        signal cVar1S9S59P063P001N035P057: std_logic_vector(   0 downto 0);
        signal cVar1S10S59P063P001P034P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S59N063P060P054P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S59N063P060P054P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S59N063P060P054P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S59N063P060P054P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S59N063P060P054P064: std_logic_vector(   0 downto 0);
        signal cVar1S16S59N063P060P054P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S59N063N060P064P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S59N063N060P064N065: std_logic_vector(   0 downto 0);
        signal cVar1S19S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S20S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S21S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S22S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S23S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S24S59N063N060N064P062: std_logic_vector(   0 downto 0);
        signal cVar1S0S60P037P063P033P017: std_logic_vector(   0 downto 0);
        signal cVar1S1S60P037P063P033P017: std_logic_vector(   0 downto 0);
        signal cVar1S2S60P037P063P033P017: std_logic_vector(   0 downto 0);
        signal cVar1S3S60P037P063P033N017: std_logic_vector(   0 downto 0);
        signal cVar1S4S60P037P063P033N017: std_logic_vector(   0 downto 0);
        signal cVar1S5S60P037P063P033N017: std_logic_vector(   0 downto 0);
        signal cVar1S6S60P037P063P033P059: std_logic_vector(   0 downto 0);
        signal cVar1S7S60P037P063P033P059: std_logic_vector(   0 downto 0);
        signal cVar1S8S60P037P063P033N059: std_logic_vector(   0 downto 0);
        signal cVar1S9S60P037P063P033N059: std_logic_vector(   0 downto 0);
        signal cVar1S10S60P037P063P033N059: std_logic_vector(   0 downto 0);
        signal cVar1S11S60P037P063P068P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S60P037P063P068P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S60P037P063P068P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S60P037P063P068N013: std_logic_vector(   0 downto 0);
        signal cVar1S15S60P037P063P068N013: std_logic_vector(   0 downto 0);
        signal cVar1S16S60P037P063P068N013: std_logic_vector(   0 downto 0);
        signal cVar1S17S60P037P063P068P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S60P037P063P068N052: std_logic_vector(   0 downto 0);
        signal cVar1S19S60P037P063P068N052: std_logic_vector(   0 downto 0);
        signal cVar1S20S60N037P035P065P022: std_logic_vector(   0 downto 0);
        signal cVar1S21S60N037P035P065P022: std_logic_vector(   0 downto 0);
        signal cVar1S22S60N037P035P065N022: std_logic_vector(   0 downto 0);
        signal cVar1S23S60N037P035P065N022: std_logic_vector(   0 downto 0);
        signal cVar1S24S60N037P035P065N022: std_logic_vector(   0 downto 0);
        signal cVar1S25S60N037P035P065P002: std_logic_vector(   0 downto 0);
        signal cVar1S26S60N037P035P065P002: std_logic_vector(   0 downto 0);
        signal cVar1S27S60N037P035P065P002: std_logic_vector(   0 downto 0);
        signal cVar1S28S60N037P035P065P041: std_logic_vector(   0 downto 0);
        signal cVar1S29S60N037P035P065P041: std_logic_vector(   0 downto 0);
        signal cVar1S30S60N037P035P065P041: std_logic_vector(   0 downto 0);
        signal cVar1S31S60N037P035N065P054: std_logic_vector(   0 downto 0);
        signal cVar1S32S60N037P035N065P054: std_logic_vector(   0 downto 0);
        signal cVar1S33S60N037P035N065P054: std_logic_vector(   0 downto 0);
        signal cVar1S34S60N037P035N065N054: std_logic_vector(   0 downto 0);
        signal cVar1S35S60N037P035N065N054: std_logic_vector(   0 downto 0);
        signal cVar1S36S60N037P035N065N054: std_logic_vector(   0 downto 0);
        signal cVar1S0S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S1S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S2S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S3S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S4S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S5S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S6S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S7S61P063P035P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S8S61P063P035P015P025: std_logic_vector(   0 downto 0);
        signal cVar1S9S61P063P035P015P025: std_logic_vector(   0 downto 0);
        signal cVar1S10S61P063P035P015N025: std_logic_vector(   0 downto 0);
        signal cVar1S11S61P063P035P015N025: std_logic_vector(   0 downto 0);
        signal cVar1S12S61P063P035P015N025: std_logic_vector(   0 downto 0);
        signal cVar1S13S61P063P035P014P047: std_logic_vector(   0 downto 0);
        signal cVar1S14S61P063P035P014P047: std_logic_vector(   0 downto 0);
        signal cVar1S15S61P063P035P014P047: std_logic_vector(   0 downto 0);
        signal cVar1S16S61P063P035N014P061: std_logic_vector(   0 downto 0);
        signal cVar1S17S61P063P035N014P061: std_logic_vector(   0 downto 0);
        signal cVar1S18S61P063P035N014P061: std_logic_vector(   0 downto 0);
        signal cVar1S19S61P063P035N014N061: std_logic_vector(   0 downto 0);
        signal cVar1S20S61P063P035N014N061: std_logic_vector(   0 downto 0);
        signal cVar1S21S61P063P035N014N061: std_logic_vector(   0 downto 0);
        signal cVar1S22S61P063P062P068P060nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S61P063P062P068N060: std_logic_vector(   0 downto 0);
        signal cVar1S24S61P063P062P068N060: std_logic_vector(   0 downto 0);
        signal cVar1S25S61P063P062P068N060: std_logic_vector(   0 downto 0);
        signal cVar1S26S61P063P062N068P022: std_logic_vector(   0 downto 0);
        signal cVar1S27S61P063P062N068P022: std_logic_vector(   0 downto 0);
        signal cVar1S28S61P063P062N068P022: std_logic_vector(   0 downto 0);
        signal cVar1S29S61P063P062N068P022: std_logic_vector(   0 downto 0);
        signal cVar1S30S61P063N062P002P035: std_logic_vector(   0 downto 0);
        signal cVar1S31S61P063N062P002N035: std_logic_vector(   0 downto 0);
        signal cVar1S32S61P063N062P002N035: std_logic_vector(   0 downto 0);
        signal cVar1S33S61P063N062P002P037: std_logic_vector(   0 downto 0);
        signal cVar1S34S61P063N062P002N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S62P062P017P048P022: std_logic_vector(   0 downto 0);
        signal cVar1S1S62P062P017P048P022: std_logic_vector(   0 downto 0);
        signal cVar1S2S62P062P017P048P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S62P062P017P048P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S62P062P017P048P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S62P062P017P048N046: std_logic_vector(   0 downto 0);
        signal cVar1S6S62P062N017P047P005: std_logic_vector(   0 downto 0);
        signal cVar1S7S62P062N017P047P005: std_logic_vector(   0 downto 0);
        signal cVar1S8S62P062N017P047P005: std_logic_vector(   0 downto 0);
        signal cVar1S9S62P062N017P047P005: std_logic_vector(   0 downto 0);
        signal cVar1S10S62P062N017P047P005: std_logic_vector(   0 downto 0);
        signal cVar1S11S62P062N017P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S62P062N017P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S13S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S14S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S15S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S17S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S18S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S19S62N062P066P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S20S62N062P066P067P016: std_logic_vector(   0 downto 0);
        signal cVar1S21S62N062P066P067P016: std_logic_vector(   0 downto 0);
        signal cVar1S22S62N062P066P067P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S62N062P066P067N016: std_logic_vector(   0 downto 0);
        signal cVar1S24S62N062P066P067N016: std_logic_vector(   0 downto 0);
        signal cVar1S25S62N062P066P067N016: std_logic_vector(   0 downto 0);
        signal cVar1S26S62N062N066P034P010: std_logic_vector(   0 downto 0);
        signal cVar1S27S62N062N066P034P010: std_logic_vector(   0 downto 0);
        signal cVar1S28S62N062N066P034P010: std_logic_vector(   0 downto 0);
        signal cVar1S29S62N062N066P034N010: std_logic_vector(   0 downto 0);
        signal cVar1S30S62N062N066P034N010: std_logic_vector(   0 downto 0);
        signal cVar1S31S62N062N066P034N010: std_logic_vector(   0 downto 0);
        signal cVar1S32S62N062N066P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S33S62N062N066P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S34S62N062N066P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S35S62N062N066P034N016: std_logic_vector(   0 downto 0);
        signal cVar1S36S62N062N066P034N016: std_logic_vector(   0 downto 0);
        signal cVar1S37S62N062N066P034N016: std_logic_vector(   0 downto 0);
        signal cVar1S0S63P067P018P050P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S63P067P018P050P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S63P067P018P050P062: std_logic_vector(   0 downto 0);
        signal cVar1S3S63P067P018P050P062: std_logic_vector(   0 downto 0);
        signal cVar1S4S63P067P018P050P062: std_logic_vector(   0 downto 0);
        signal cVar1S5S63P067P018P050P010: std_logic_vector(   0 downto 0);
        signal cVar1S6S63P067P018P050N010: std_logic_vector(   0 downto 0);
        signal cVar1S7S63P067P018P050N010: std_logic_vector(   0 downto 0);
        signal cVar1S8S63P067N018P068P049: std_logic_vector(   0 downto 0);
        signal cVar1S9S63P067N018P068P049: std_logic_vector(   0 downto 0);
        signal cVar1S10S63P067N018N068P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S63P067N018N068P015: std_logic_vector(   0 downto 0);
        signal cVar1S12S63P067N018N068P015: std_logic_vector(   0 downto 0);
        signal cVar1S13S63P067N018N068N015: std_logic_vector(   0 downto 0);
        signal cVar1S14S63P067N018N068N015: std_logic_vector(   0 downto 0);
        signal cVar1S15S63P067N018N068N015: std_logic_vector(   0 downto 0);
        signal cVar1S16S63N067P044P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S63N067P044N028P023: std_logic_vector(   0 downto 0);
        signal cVar1S18S63N067P044N028N023: std_logic_vector(   0 downto 0);
        signal cVar1S19S63N067P044N028N023: std_logic_vector(   0 downto 0);
        signal cVar1S20S63N067P044N028N023: std_logic_vector(   0 downto 0);
        signal cVar1S21S63N067P044N028N023: std_logic_vector(   0 downto 0);
        signal cVar1S22S63N067N044P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S23S63N067N044P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S24S63N067N044P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S25S63N067N044P059P049: std_logic_vector(   0 downto 0);
        signal cVar1S26S63N067N044N059P031: std_logic_vector(   0 downto 0);
        signal cVar1S27S63N067N044N059P031: std_logic_vector(   0 downto 0);
        signal cVar1S28S63N067N044N059P031: std_logic_vector(   0 downto 0);
        signal cVar1S29S63N067N044N059N031: std_logic_vector(   0 downto 0);
        signal cVar1S30S63N067N044N059N031: std_logic_vector(   0 downto 0);
        signal cVar1S31S63N067N044N059N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S64P059P061P058P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S64P059P061P058P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S64P059P061P058N032: std_logic_vector(   0 downto 0);
        signal cVar1S3S64P059P061P058N032: std_logic_vector(   0 downto 0);
        signal cVar1S4S64P059P061P058N032: std_logic_vector(   0 downto 0);
        signal cVar1S5S64P059P061N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S6S64P059P061N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S64P059P061N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S8S64P059P061N058P033: std_logic_vector(   0 downto 0);
        signal cVar1S9S64P059P061P067P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S64P059P061P067N069: std_logic_vector(   0 downto 0);
        signal cVar1S11S64P059P061P067P037: std_logic_vector(   0 downto 0);
        signal cVar1S12S64P059P049P030P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S64P059P049P030P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S64P059P049P030P004: std_logic_vector(   0 downto 0);
        signal cVar1S15S64P059P049N030P005: std_logic_vector(   0 downto 0);
        signal cVar1S16S64P059P049N030P005: std_logic_vector(   0 downto 0);
        signal cVar1S17S64P059P049N030P005: std_logic_vector(   0 downto 0);
        signal cVar1S18S64P059P049N030P005: std_logic_vector(   0 downto 0);
        signal cVar1S19S64P059P049N030P005: std_logic_vector(   0 downto 0);
        signal cVar1S20S64P059P049P055P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S64P059P049P055N051: std_logic_vector(   0 downto 0);
        signal cVar1S0S65P058P054P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S65P058P054P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S2S65P058P054N047P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S65P058P054N047P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S65P058P054N047P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S65P058P054N047N013: std_logic_vector(   0 downto 0);
        signal cVar1S6S65P058P054N047N013: std_logic_vector(   0 downto 0);
        signal cVar1S7S65P058P054N047N013: std_logic_vector(   0 downto 0);
        signal cVar1S8S65P058P054P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S65P058P054P015N013: std_logic_vector(   0 downto 0);
        signal cVar1S10S65P058P054N015P033: std_logic_vector(   0 downto 0);
        signal cVar1S11S65P058P054N015P033: std_logic_vector(   0 downto 0);
        signal cVar1S12S65P058P054N015N033: std_logic_vector(   0 downto 0);
        signal cVar1S13S65N058P043P022P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S65N058P043P022N003: std_logic_vector(   0 downto 0);
        signal cVar1S15S65N058P043P022N003: std_logic_vector(   0 downto 0);
        signal cVar1S16S65N058P043N022P047: std_logic_vector(   0 downto 0);
        signal cVar1S17S65N058P043N022P047: std_logic_vector(   0 downto 0);
        signal cVar1S18S65N058P043N022P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S65N058N043P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S20S65N058N043P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S21S65N058N043P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S22S65N058N043P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S23S65N058N043P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S24S65N058N043N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S25S65N058N043N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S26S65N058N043N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S27S65N058N043N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S0S66P015P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S66P015P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S66P015P044N025N023: std_logic_vector(   0 downto 0);
        signal cVar1S3S66P015P044N025N023: std_logic_vector(   0 downto 0);
        signal cVar1S4S66P015N044P003P055: std_logic_vector(   0 downto 0);
        signal cVar1S5S66P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S6S66P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S7S66P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S8S66P015N044N003P027: std_logic_vector(   0 downto 0);
        signal cVar1S9S66P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S10S66P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S66P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S12S66N015P063P037P067: std_logic_vector(   0 downto 0);
        signal cVar1S13S66N015P063P037P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S66N015P063P037P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S66N015P063P037P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S66N015P063P037P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S66N015P063N037P017: std_logic_vector(   0 downto 0);
        signal cVar1S18S66N015P063N037P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S66N015P063N037P017: std_logic_vector(   0 downto 0);
        signal cVar1S20S66N015P063N037N017: std_logic_vector(   0 downto 0);
        signal cVar1S21S66N015P063N037N017: std_logic_vector(   0 downto 0);
        signal cVar1S22S66N015P063N037N017: std_logic_vector(   0 downto 0);
        signal cVar1S23S66N015N063P029P058: std_logic_vector(   0 downto 0);
        signal cVar1S24S66N015N063P029P058: std_logic_vector(   0 downto 0);
        signal cVar1S25S66N015N063P029P058: std_logic_vector(   0 downto 0);
        signal cVar1S26S66N015N063P029P058: std_logic_vector(   0 downto 0);
        signal cVar1S27S66N015N063P029P058: std_logic_vector(   0 downto 0);
        signal cVar1S28S66N015N063N029P028: std_logic_vector(   0 downto 0);
        signal cVar1S29S66N015N063N029P028: std_logic_vector(   0 downto 0);
        signal cVar1S30S66N015N063N029N028: std_logic_vector(   0 downto 0);
        signal cVar1S31S66N015N063N029N028: std_logic_vector(   0 downto 0);
        signal cVar1S32S66N015N063N029N028: std_logic_vector(   0 downto 0);
        signal cVar1S33S66N015N063N029N028: std_logic_vector(   0 downto 0);
        signal cVar1S0S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S1S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S2S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S3S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S4S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S5S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S6S67P015P014P050P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S67P015P014P050P011: std_logic_vector(   0 downto 0);
        signal cVar1S8S67P015P014P050P011: std_logic_vector(   0 downto 0);
        signal cVar1S9S67P015P014P050N011: std_logic_vector(   0 downto 0);
        signal cVar1S10S67P015P014P050N011: std_logic_vector(   0 downto 0);
        signal cVar1S11S67P015P014P050N011: std_logic_vector(   0 downto 0);
        signal cVar1S12S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S14S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S15S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S16S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S17S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S18S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S19S67P015P014P021P012: std_logic_vector(   0 downto 0);
        signal cVar1S20S67P015P044P031P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S67P015P044P031N006: std_logic_vector(   0 downto 0);
        signal cVar1S22S67P015P044P031N006: std_logic_vector(   0 downto 0);
        signal cVar1S23S67P015N044P003P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S24S67P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S25S67P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S26S67P015N044P003N055: std_logic_vector(   0 downto 0);
        signal cVar1S27S67P015N044N003P027: std_logic_vector(   0 downto 0);
        signal cVar1S28S67P015N044N003P027: std_logic_vector(   0 downto 0);
        signal cVar1S29S67P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S30S67P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S31S67P015N044N003N027: std_logic_vector(   0 downto 0);
        signal cVar1S0S68P014P012P021P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S68P014P012P021P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S68P014P012P021P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S68P014P012P021N032: std_logic_vector(   0 downto 0);
        signal cVar1S4S68P014P012P021N032: std_logic_vector(   0 downto 0);
        signal cVar1S5S68P014P012P021N032: std_logic_vector(   0 downto 0);
        signal cVar1S6S68P014P012P021N032: std_logic_vector(   0 downto 0);
        signal cVar1S7S68P014P012P021P026: std_logic_vector(   0 downto 0);
        signal cVar1S8S68P014P012P001P010nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S68P014P012P001N010: std_logic_vector(   0 downto 0);
        signal cVar1S10S68P014P012P001N010: std_logic_vector(   0 downto 0);
        signal cVar1S11S68P014P012N001P009: std_logic_vector(   0 downto 0);
        signal cVar1S12S68P014P012N001P009: std_logic_vector(   0 downto 0);
        signal cVar1S13S68P014P012N001P009: std_logic_vector(   0 downto 0);
        signal cVar1S14S68P014P012N001P009: std_logic_vector(   0 downto 0);
        signal cVar1S15S68N014P027P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S68N014P027P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S68N014P027P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S18S68N014P027P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S19S68N014P027N009P026: std_logic_vector(   0 downto 0);
        signal cVar1S20S68N014P027N009P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S68N014P027N009P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S68N014N027P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S23S68N014N027P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S24S68N014N027P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S25S68N014N027P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S26S68N014N027P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S27S68N014N027P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S28S68N014N027P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S29S68N014N027P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S30S68N014N027P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S31S68N014N027P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S32S68N014N027P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S33S68N014N027P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S0S69P017P062P034P064: std_logic_vector(   0 downto 0);
        signal cVar1S1S69P017P062P034P064: std_logic_vector(   0 downto 0);
        signal cVar1S2S69P017P062P034P064: std_logic_vector(   0 downto 0);
        signal cVar1S3S69P017P062P034P064: std_logic_vector(   0 downto 0);
        signal cVar1S4S69P017P062P034N064: std_logic_vector(   0 downto 0);
        signal cVar1S5S69P017P062P034N064: std_logic_vector(   0 downto 0);
        signal cVar1S6S69P017P062P034N064: std_logic_vector(   0 downto 0);
        signal cVar1S7S69P017P062P034P060: std_logic_vector(   0 downto 0);
        signal cVar1S8S69P017P062P034P060: std_logic_vector(   0 downto 0);
        signal cVar1S9S69P017P062P034N060: std_logic_vector(   0 downto 0);
        signal cVar1S10S69P017P062P034N060: std_logic_vector(   0 downto 0);
        signal cVar1S11S69P017P062P034N060: std_logic_vector(   0 downto 0);
        signal cVar1S12S69P017P062P034N060: std_logic_vector(   0 downto 0);
        signal cVar1S13S69P017N062P014P054: std_logic_vector(   0 downto 0);
        signal cVar1S14S69P017N062P014P054: std_logic_vector(   0 downto 0);
        signal cVar1S15S69P017N062P014P054: std_logic_vector(   0 downto 0);
        signal cVar1S16S69P017N062P014N054: std_logic_vector(   0 downto 0);
        signal cVar1S17S69P017N062P014N054: std_logic_vector(   0 downto 0);
        signal cVar1S18S69P017N062P014N054: std_logic_vector(   0 downto 0);
        signal cVar1S19S69P017N062P014P035: std_logic_vector(   0 downto 0);
        signal cVar1S20S69P017N062P014P035: std_logic_vector(   0 downto 0);
        signal cVar1S21S69P017N062P014P035: std_logic_vector(   0 downto 0);
        signal cVar1S22S69P017N062P014P035: std_logic_vector(   0 downto 0);
        signal cVar1S23S69P017N062P014P035: std_logic_vector(   0 downto 0);
        signal cVar1S24S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S25S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S26S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S27S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S28S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S29S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S30S69N017P066P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S31S69N017P066P028P030: std_logic_vector(   0 downto 0);
        signal cVar1S32S69N017N066P047P049: std_logic_vector(   0 downto 0);
        signal cVar1S33S69N017N066P047P049: std_logic_vector(   0 downto 0);
        signal cVar1S34S69N017N066P047P049: std_logic_vector(   0 downto 0);
        signal cVar1S35S69N017N066P047N049: std_logic_vector(   0 downto 0);
        signal cVar1S36S69N017N066P047N049: std_logic_vector(   0 downto 0);
        signal cVar1S37S69N017N066P047N049: std_logic_vector(   0 downto 0);
        signal cVar1S38S69N017N066N047P023: std_logic_vector(   0 downto 0);
        signal cVar1S39S69N017N066N047P023: std_logic_vector(   0 downto 0);
        signal cVar1S40S69N017N066N047N023: std_logic_vector(   0 downto 0);
        signal cVar1S41S69N017N066N047N023: std_logic_vector(   0 downto 0);
        signal cVar1S42S69N017N066N047N023: std_logic_vector(   0 downto 0);
        signal cVar1S43S69N017N066N047N023: std_logic_vector(   0 downto 0);
        signal cVar1S0S70P017P014P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S70P017P014P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S70P017P014P062N010: std_logic_vector(   0 downto 0);
        signal cVar1S3S70P017P014P062N010: std_logic_vector(   0 downto 0);
        signal cVar1S4S70P017P014P062N010: std_logic_vector(   0 downto 0);
        signal cVar1S5S70P017P014P062P033: std_logic_vector(   0 downto 0);
        signal cVar1S6S70P017P014P062N033: std_logic_vector(   0 downto 0);
        signal cVar1S7S70P017P014P062N033: std_logic_vector(   0 downto 0);
        signal cVar1S8S70P017P014P012P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S70P017P014P012N041: std_logic_vector(   0 downto 0);
        signal cVar1S10S70P017P014P012P049: std_logic_vector(   0 downto 0);
        signal cVar1S11S70P017P014P012P049: std_logic_vector(   0 downto 0);
        signal cVar1S12S70P017P014P012P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S70N017P066P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S70N017P066P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S70N017P066P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S16S70N017P066P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S17S70N017P066P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S18S70N017P066P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S70N017P066P044P045: std_logic_vector(   0 downto 0);
        signal cVar1S20S70N017P066P044P045: std_logic_vector(   0 downto 0);
        signal cVar1S21S70N017P066P044P045: std_logic_vector(   0 downto 0);
        signal cVar1S22S70N017P066P004P034: std_logic_vector(   0 downto 0);
        signal cVar1S23S70N017P066P004N034: std_logic_vector(   0 downto 0);
        signal cVar1S24S70N017P066P004N034: std_logic_vector(   0 downto 0);
        signal cVar1S25S70N017P066P004P061nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S70N017P066P004N061: std_logic_vector(   0 downto 0);
        signal cVar1S27S70N017P066P004N061: std_logic_vector(   0 downto 0);
        signal cVar1S0S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S1S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S2S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S3S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S4S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S5S71P067P015P018P069: std_logic_vector(   0 downto 0);
        signal cVar1S6S71P067P015N018P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S71P067P015N018P002: std_logic_vector(   0 downto 0);
        signal cVar1S8S71P067P015N018N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S71P067P015N018N002: std_logic_vector(   0 downto 0);
        signal cVar1S10S71P067P015N018N002: std_logic_vector(   0 downto 0);
        signal cVar1S11S71P067P015N018N002: std_logic_vector(   0 downto 0);
        signal cVar1S12S71P067P015P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S13S71P067P015P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S14S71P067P015P017P069: std_logic_vector(   0 downto 0);
        signal cVar1S15S71P067P015P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S16S71P067P015P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S17S71P067P015P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S18S71P067P015P017N069: std_logic_vector(   0 downto 0);
        signal cVar1S19S71P067P015N017P026: std_logic_vector(   0 downto 0);
        signal cVar1S20S71P067P015N017P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S71P067P015N017P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S71P067P015N017P026: std_logic_vector(   0 downto 0);
        signal cVar1S23S71P067P001P057P037: std_logic_vector(   0 downto 0);
        signal cVar1S24S71P067P001P057P037: std_logic_vector(   0 downto 0);
        signal cVar1S25S71P067P001P057P037: std_logic_vector(   0 downto 0);
        signal cVar1S26S71P067P001P057P037: std_logic_vector(   0 downto 0);
        signal cVar1S27S71P067N001P003P054: std_logic_vector(   0 downto 0);
        signal cVar1S28S71P067N001P003P054: std_logic_vector(   0 downto 0);
        signal cVar1S29S71P067N001N003P045: std_logic_vector(   0 downto 0);
        signal cVar1S30S71P067N001N003P045: std_logic_vector(   0 downto 0);
        signal cVar1S31S71P067N001N003P045: std_logic_vector(   0 downto 0);
        signal cVar1S32S71P067N001N003P045: std_logic_vector(   0 downto 0);
        signal cVar1S0S72P069P045P052P056: std_logic_vector(   0 downto 0);
        signal cVar1S1S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S2S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S3S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S4S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S5S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S6S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S7S72P069P045N052P029: std_logic_vector(   0 downto 0);
        signal cVar1S8S72P069P045P018P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S72P069P045P018N006: std_logic_vector(   0 downto 0);
        signal cVar1S10S72P069P045P018P047: std_logic_vector(   0 downto 0);
        signal cVar1S11S72N069P015P027P008: std_logic_vector(   0 downto 0);
        signal cVar1S12S72N069P015P027P008: std_logic_vector(   0 downto 0);
        signal cVar1S13S72N069P015P027N008: std_logic_vector(   0 downto 0);
        signal cVar1S14S72N069P015P027N008: std_logic_vector(   0 downto 0);
        signal cVar1S15S72N069P015N027P000: std_logic_vector(   0 downto 0);
        signal cVar1S16S72N069P015N027P000: std_logic_vector(   0 downto 0);
        signal cVar1S17S72N069P015N027P000: std_logic_vector(   0 downto 0);
        signal cVar1S18S72N069P015N027P000: std_logic_vector(   0 downto 0);
        signal cVar1S19S72N069P015N027P000: std_logic_vector(   0 downto 0);
        signal cVar1S20S72N069P015P028P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S72N069P015P028P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S72N069P015P028P026: std_logic_vector(   0 downto 0);
        signal cVar1S23S72N069P015N028P020: std_logic_vector(   0 downto 0);
        signal cVar1S24S72N069P015N028P020: std_logic_vector(   0 downto 0);
        signal cVar1S25S72N069P015N028P020: std_logic_vector(   0 downto 0);
        signal cVar1S26S72N069P015N028P020: std_logic_vector(   0 downto 0);
        signal cVar1S27S72N069P015N028P020: std_logic_vector(   0 downto 0);
        signal cVar1S0S73P016P038P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S1S73P016P038P043N045: std_logic_vector(   0 downto 0);
        signal cVar1S2S73P016P038P043N045: std_logic_vector(   0 downto 0);
        signal cVar1S3S73P016P038P043N045: std_logic_vector(   0 downto 0);
        signal cVar1S4S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S5S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S6S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S7S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S8S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S73P016P038N043P045: std_logic_vector(   0 downto 0);
        signal cVar1S11S73P016P038P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S12S73P016P038P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S16S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S18S73N016P036P027P014: std_logic_vector(   0 downto 0);
        signal cVar1S19S73N016P036N027P038: std_logic_vector(   0 downto 0);
        signal cVar1S20S73N016P036N027P038: std_logic_vector(   0 downto 0);
        signal cVar1S21S73N016P036N027P038: std_logic_vector(   0 downto 0);
        signal cVar1S22S73N016P036N027N038: std_logic_vector(   0 downto 0);
        signal cVar1S23S73N016P036N027N038: std_logic_vector(   0 downto 0);
        signal cVar1S24S73N016P036N027N038: std_logic_vector(   0 downto 0);
        signal cVar1S25S73N016P036N027N038: std_logic_vector(   0 downto 0);
        signal cVar1S26S73N016P036P045P068: std_logic_vector(   0 downto 0);
        signal cVar1S27S73N016P036P045P068: std_logic_vector(   0 downto 0);
        signal cVar1S28S73N016P036P045P068: std_logic_vector(   0 downto 0);
        signal cVar1S29S73N016P036P045P068: std_logic_vector(   0 downto 0);
        signal cVar1S30S73N016P036P045P043: std_logic_vector(   0 downto 0);
        signal cVar1S0S74P016P053P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S1S74P016P053P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S2S74P016P053P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S3S74P016P053P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S4S74P016P053P035N026: std_logic_vector(   0 downto 0);
        signal cVar1S5S74P016P053P035N026: std_logic_vector(   0 downto 0);
        signal cVar1S6S74P016P053P035N026: std_logic_vector(   0 downto 0);
        signal cVar1S7S74P016P053P035P052: std_logic_vector(   0 downto 0);
        signal cVar1S8S74P016P053P035P052: std_logic_vector(   0 downto 0);
        signal cVar1S9S74P016P053P035P052: std_logic_vector(   0 downto 0);
        signal cVar1S10S74P016P053P035N052: std_logic_vector(   0 downto 0);
        signal cVar1S11S74P016P053P030P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S74P016P053P030P019: std_logic_vector(   0 downto 0);
        signal cVar1S13S74P016P053P030P019: std_logic_vector(   0 downto 0);
        signal cVar1S14S74P016P053N030P059: std_logic_vector(   0 downto 0);
        signal cVar1S15S74P016P053N030P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S74P016P053N030P059: std_logic_vector(   0 downto 0);
        signal cVar1S17S74P016P043P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S74P016P043N062P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S74P016P043N062N022: std_logic_vector(   0 downto 0);
        signal cVar1S20S74P016P043N062N022: std_logic_vector(   0 downto 0);
        signal cVar1S21S74P016N043P038P056: std_logic_vector(   0 downto 0);
        signal cVar1S22S74P016N043P038P056: std_logic_vector(   0 downto 0);
        signal cVar1S23S74P016N043P038P056: std_logic_vector(   0 downto 0);
        signal cVar1S24S74P016N043P038P056: std_logic_vector(   0 downto 0);
        signal cVar1S25S74P016N043P038P056: std_logic_vector(   0 downto 0);
        signal cVar1S26S74P016N043P038P033: std_logic_vector(   0 downto 0);
        signal cVar1S27S74P016N043P038P033: std_logic_vector(   0 downto 0);
        signal cVar1S0S75P064P027P026P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S75P064P027P026P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S75P064P027P026N006: std_logic_vector(   0 downto 0);
        signal cVar1S3S75P064P027P026N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S75P064P027P026P010: std_logic_vector(   0 downto 0);
        signal cVar1S5S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S6S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S7S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S8S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S9S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S10S75P064N027P060P054: std_logic_vector(   0 downto 0);
        signal cVar1S11S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S15S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S16S75P064N027N060P062: std_logic_vector(   0 downto 0);
        signal cVar1S17S75P064P003P046P058: std_logic_vector(   0 downto 0);
        signal cVar1S18S75P064P003P046N058: std_logic_vector(   0 downto 0);
        signal cVar1S19S75P064P003P046N058: std_logic_vector(   0 downto 0);
        signal cVar1S20S75P064P003P046N058: std_logic_vector(   0 downto 0);
        signal cVar1S21S75P064N003P018P065: std_logic_vector(   0 downto 0);
        signal cVar1S22S75P064N003P018P065: std_logic_vector(   0 downto 0);
        signal cVar1S23S75P064N003P018P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S75P064N003P018P065: std_logic_vector(   0 downto 0);
        signal cVar1S25S75P064N003P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S26S75P064N003P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S27S75P064N003P018N065: std_logic_vector(   0 downto 0);
        signal cVar1S28S75P064N003N018P013: std_logic_vector(   0 downto 0);
        signal cVar1S29S75P064N003N018P013: std_logic_vector(   0 downto 0);
        signal cVar1S30S75P064N003N018P013: std_logic_vector(   0 downto 0);
        signal cVar1S31S75P064N003N018N013: std_logic_vector(   0 downto 0);
        signal cVar1S32S75P064N003N018N013: std_logic_vector(   0 downto 0);
        signal cVar1S33S75P064N003N018N013: std_logic_vector(   0 downto 0);
        signal cVar1S0S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S5S76P016P060P056P067: std_logic_vector(   0 downto 0);
        signal cVar1S6S76P016P060P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S76P016P060P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S8S76P016P060P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S9S76P016P060P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S10S76P016P060P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S11S76P016P060P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S76P016P060P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S76P016P060P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S76P016P060P015P020: std_logic_vector(   0 downto 0);
        signal cVar1S15S76P016P060P015P020: std_logic_vector(   0 downto 0);
        signal cVar1S16S76N016P064P048P062: std_logic_vector(   0 downto 0);
        signal cVar1S17S76N016P064P048P062: std_logic_vector(   0 downto 0);
        signal cVar1S18S76N016P064P048P062: std_logic_vector(   0 downto 0);
        signal cVar1S19S76N016P064P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S20S76N016P064P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S21S76N016P064P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S22S76N016P064P048P058: std_logic_vector(   0 downto 0);
        signal cVar1S23S76N016P064P048P058: std_logic_vector(   0 downto 0);
        signal cVar1S24S76N016N064P027P006: std_logic_vector(   0 downto 0);
        signal cVar1S25S76N016N064P027N006: std_logic_vector(   0 downto 0);
        signal cVar1S26S76N016N064P027N006: std_logic_vector(   0 downto 0);
        signal cVar1S27S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S28S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S29S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S30S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S31S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S32S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S33S76N016N064N027P057: std_logic_vector(   0 downto 0);
        signal cVar1S0S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S1S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S2S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S3S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S4S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S5S77P035P053P016P057: std_logic_vector(   0 downto 0);
        signal cVar1S6S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S7S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S8S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S9S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S10S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S11S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S12S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S13S77P035P053P016P028: std_logic_vector(   0 downto 0);
        signal cVar1S14S77P035P053P016N028: std_logic_vector(   0 downto 0);
        signal cVar1S15S77P035P053N016P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S77P035P053N016P059: std_logic_vector(   0 downto 0);
        signal cVar1S17S77P035P053N016P059: std_logic_vector(   0 downto 0);
        signal cVar1S18S77P035P053N016P059: std_logic_vector(   0 downto 0);
        signal cVar1S19S77P035P053N016P059: std_logic_vector(   0 downto 0);
        signal cVar1S20S77P035P052P012P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S77P035P052P012N029: std_logic_vector(   0 downto 0);
        signal cVar1S22S77P035P052P012N029: std_logic_vector(   0 downto 0);
        signal cVar1S23S77P035P052P012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S24S77P035N052P046P033: std_logic_vector(   0 downto 0);
        signal cVar1S25S77P035N052P046P033: std_logic_vector(   0 downto 0);
        signal cVar1S26S77P035N052N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S27S77P035N052N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S28S77P035N052N046N051: std_logic_vector(   0 downto 0);
        signal cVar1S29S77P035N052N046N051: std_logic_vector(   0 downto 0);
        signal cVar1S30S77P035N052N046N051: std_logic_vector(   0 downto 0);
        signal cVar1S0S78P035P064P052P036nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S78P035P064P052N036: std_logic_vector(   0 downto 0);
        signal cVar1S2S78P035P064P052N036: std_logic_vector(   0 downto 0);
        signal cVar1S3S78P035P064P052N036: std_logic_vector(   0 downto 0);
        signal cVar1S4S78P035P064N052P037: std_logic_vector(   0 downto 0);
        signal cVar1S5S78P035P064N052P037: std_logic_vector(   0 downto 0);
        signal cVar1S6S78P035P064N052P037: std_logic_vector(   0 downto 0);
        signal cVar1S7S78P035P064N052P037: std_logic_vector(   0 downto 0);
        signal cVar1S8S78P035P064N052N037: std_logic_vector(   0 downto 0);
        signal cVar1S9S78P035P064N052N037: std_logic_vector(   0 downto 0);
        signal cVar1S10S78P035P064N052N037: std_logic_vector(   0 downto 0);
        signal cVar1S11S78P035N064P012P001: std_logic_vector(   0 downto 0);
        signal cVar1S12S78P035N064P012P001: std_logic_vector(   0 downto 0);
        signal cVar1S13S78P035N064P012P001: std_logic_vector(   0 downto 0);
        signal cVar1S14S78P035N064P012P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S78P035N064P012P036: std_logic_vector(   0 downto 0);
        signal cVar1S16S78P035N064P012N036: std_logic_vector(   0 downto 0);
        signal cVar1S17S78N035P016P064P015: std_logic_vector(   0 downto 0);
        signal cVar1S18S78N035P016P064P015: std_logic_vector(   0 downto 0);
        signal cVar1S19S78N035P016P064N015: std_logic_vector(   0 downto 0);
        signal cVar1S20S78N035P016P064N015: std_logic_vector(   0 downto 0);
        signal cVar1S21S78N035P016P064N015: std_logic_vector(   0 downto 0);
        signal cVar1S22S78N035P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S23S78N035P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S24S78N035P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S25S78N035P016P064P048: std_logic_vector(   0 downto 0);
        signal cVar1S26S78N035P016P053P004: std_logic_vector(   0 downto 0);
        signal cVar1S27S78N035P016P053P004: std_logic_vector(   0 downto 0);
        signal cVar1S28S78N035P016P053P004: std_logic_vector(   0 downto 0);
        signal cVar1S29S78N035P016N053P028: std_logic_vector(   0 downto 0);
        signal cVar1S30S78N035P016N053P028: std_logic_vector(   0 downto 0);
        signal cVar1S31S78N035P016N053P028: std_logic_vector(   0 downto 0);
        signal cVar1S32S78N035P016N053P028: std_logic_vector(   0 downto 0);
        signal cVar1S33S78N035P016N053P028: std_logic_vector(   0 downto 0);
        signal cVar1S0S79P064P035P052P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S79P064P035N052P055: std_logic_vector(   0 downto 0);
        signal cVar1S2S79P064P035N052P055: std_logic_vector(   0 downto 0);
        signal cVar1S3S79P064P035N052P055: std_logic_vector(   0 downto 0);
        signal cVar1S4S79P064P035N052P055: std_logic_vector(   0 downto 0);
        signal cVar1S5S79P064P035N052P055: std_logic_vector(   0 downto 0);
        signal cVar1S6S79P064N035P051P048: std_logic_vector(   0 downto 0);
        signal cVar1S7S79P064N035P051P048: std_logic_vector(   0 downto 0);
        signal cVar1S8S79P064N035P051P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S79P064N035P051P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S79P064N035P051P069: std_logic_vector(   0 downto 0);
        signal cVar1S11S79N064P035P016P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S79N064P035P016P026: std_logic_vector(   0 downto 0);
        signal cVar1S13S79N064P035P016N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S79N064P035P016N026: std_logic_vector(   0 downto 0);
        signal cVar1S15S79N064P035P016N026: std_logic_vector(   0 downto 0);
        signal cVar1S16S79N064P035P016N026: std_logic_vector(   0 downto 0);
        signal cVar1S17S79N064P035P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S18S79N064P035P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S19S79N064P035P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S20S79N064P035P016N052: std_logic_vector(   0 downto 0);
        signal cVar1S21S79N064P035P016N052: std_logic_vector(   0 downto 0);
        signal cVar1S22S79N064P035P013P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S79N064P035P013N016: std_logic_vector(   0 downto 0);
        signal cVar1S24S79N064P035P013N016: std_logic_vector(   0 downto 0);
        signal cVar1S25S79N064P035P013N016: std_logic_vector(   0 downto 0);
        signal cVar1S26S79N064P035P013P030: std_logic_vector(   0 downto 0);
        signal cVar1S27S79N064P035P013P030: std_logic_vector(   0 downto 0);
        signal cVar1S28S79N064P035P013N030: std_logic_vector(   0 downto 0);
        signal cVar1S29S79N064P035P013N030: std_logic_vector(   0 downto 0);
        signal cVar1S0S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S1S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S2S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S3S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S4S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S5S80P037P034P057P058: std_logic_vector(   0 downto 0);
        signal cVar1S6S80P037P034P057P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S80P037P034P057P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S80P037P034P057N014: std_logic_vector(   0 downto 0);
        signal cVar1S9S80P037N034P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S10S80P037N034P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S11S80P037N034P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S12S80P037N034P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S80P037N034P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S14S80P037N034N017P012: std_logic_vector(   0 downto 0);
        signal cVar1S15S80P037N034N017P012: std_logic_vector(   0 downto 0);
        signal cVar1S16S80P037N034N017P012: std_logic_vector(   0 downto 0);
        signal cVar1S17S80P037N034N017N012: std_logic_vector(   0 downto 0);
        signal cVar1S18S80P037N034N017N012: std_logic_vector(   0 downto 0);
        signal cVar1S19S80P037N034N017N012: std_logic_vector(   0 downto 0);
        signal cVar1S20S80P037P015P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S80P037P015P052N029: std_logic_vector(   0 downto 0);
        signal cVar1S22S80P037P015N052P025: std_logic_vector(   0 downto 0);
        signal cVar1S23S80P037P015N052P025: std_logic_vector(   0 downto 0);
        signal cVar1S24S80P037P015N052N025: std_logic_vector(   0 downto 0);
        signal cVar1S25S80P037P015N052N025: std_logic_vector(   0 downto 0);
        signal cVar1S26S80P037N015P018P055: std_logic_vector(   0 downto 0);
        signal cVar1S27S80P037N015P018P055: std_logic_vector(   0 downto 0);
        signal cVar1S28S80P037N015P018P055: std_logic_vector(   0 downto 0);
        signal cVar1S29S80P037N015P018P055: std_logic_vector(   0 downto 0);
        signal cVar1S30S80P037N015P018P055: std_logic_vector(   0 downto 0);
        signal cVar1S31S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S32S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S33S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S34S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S35S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S36S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S37S80P037N015N018P034: std_logic_vector(   0 downto 0);
        signal cVar1S0S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S1S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S2S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S3S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S5S81P037P032P017P056: std_logic_vector(   0 downto 0);
        signal cVar1S6S81P037P032P017P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S81P037P032P017P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S81P037P032P017N036: std_logic_vector(   0 downto 0);
        signal cVar1S9S81P037P032P017N036: std_logic_vector(   0 downto 0);
        signal cVar1S10S81P037P032P013P031: std_logic_vector(   0 downto 0);
        signal cVar1S11S81P037P032P013P031: std_logic_vector(   0 downto 0);
        signal cVar1S12S81P037P032P013P031: std_logic_vector(   0 downto 0);
        signal cVar1S13S81P037P032P013P031: std_logic_vector(   0 downto 0);
        signal cVar1S14S81P037P032P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S15S81P037P032P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S81P037P032P013P059: std_logic_vector(   0 downto 0);
        signal cVar1S17S81P037P032P013N059: std_logic_vector(   0 downto 0);
        signal cVar1S18S81P037P032P013N059: std_logic_vector(   0 downto 0);
        signal cVar1S19S81P037P052P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S81P037P052P008N013: std_logic_vector(   0 downto 0);
        signal cVar1S21S81P037P052P008N013: std_logic_vector(   0 downto 0);
        signal cVar1S22S81P037P052P008N013: std_logic_vector(   0 downto 0);
        signal cVar1S23S81P037P052N008P068: std_logic_vector(   0 downto 0);
        signal cVar1S24S81P037P052N008P068: std_logic_vector(   0 downto 0);
        signal cVar1S25S81P037P052N008P068: std_logic_vector(   0 downto 0);
        signal cVar1S26S81P037P052N008N068: std_logic_vector(   0 downto 0);
        signal cVar1S27S81P037P052N008N068: std_logic_vector(   0 downto 0);
        signal cVar1S28S81P037P052N008N068: std_logic_vector(   0 downto 0);
        signal cVar1S29S81P037N052P025P044nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S81P037N052P025N044: std_logic_vector(   0 downto 0);
        signal cVar1S31S81P037N052P025N044: std_logic_vector(   0 downto 0);
        signal cVar1S32S81P037N052N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S33S81P037N052N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S34S81P037N052N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S35S81P037N052N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S36S81P037N052N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S37S81P037N052N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S38S81P037N052N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S0S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S1S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S2S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S3S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S4S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S5S82P037P031P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S6S82P037P031P054P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S82P037P031P054N065: std_logic_vector(   0 downto 0);
        signal cVar1S8S82P037P031P054N065: std_logic_vector(   0 downto 0);
        signal cVar1S9S82P037P031P054N065: std_logic_vector(   0 downto 0);
        signal cVar1S10S82P037P031P058P007: std_logic_vector(   0 downto 0);
        signal cVar1S11S82P037P031N058P054: std_logic_vector(   0 downto 0);
        signal cVar1S12S82P037P031N058P054: std_logic_vector(   0 downto 0);
        signal cVar1S13S82P037P031N058N054: std_logic_vector(   0 downto 0);
        signal cVar1S14S82N037P017P044P060: std_logic_vector(   0 downto 0);
        signal cVar1S15S82N037P017N044P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S82N037P017N044P023: std_logic_vector(   0 downto 0);
        signal cVar1S17S82N037P017N044P023: std_logic_vector(   0 downto 0);
        signal cVar1S18S82N037P017N044P023: std_logic_vector(   0 downto 0);
        signal cVar1S19S82N037P017N044P023: std_logic_vector(   0 downto 0);
        signal cVar1S20S82N037N017P029P009: std_logic_vector(   0 downto 0);
        signal cVar1S21S82N037N017P029P009: std_logic_vector(   0 downto 0);
        signal cVar1S22S82N037N017P029N009: std_logic_vector(   0 downto 0);
        signal cVar1S23S82N037N017P029N009: std_logic_vector(   0 downto 0);
        signal cVar1S24S82N037N017N029P067: std_logic_vector(   0 downto 0);
        signal cVar1S25S82N037N017N029N067: std_logic_vector(   0 downto 0);
        signal cVar1S0S83P017P037P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S1S83P017P037P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S2S83P017P037P000P047: std_logic_vector(   0 downto 0);
        signal cVar1S3S83P017P037P000N047: std_logic_vector(   0 downto 0);
        signal cVar1S4S83P017P037P000N047: std_logic_vector(   0 downto 0);
        signal cVar1S5S83P017P037P000N047: std_logic_vector(   0 downto 0);
        signal cVar1S6S83P017P037P000P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S83P017P037P000N021: std_logic_vector(   0 downto 0);
        signal cVar1S8S83P017P037P019P003: std_logic_vector(   0 downto 0);
        signal cVar1S9S83P017P037P019N003: std_logic_vector(   0 downto 0);
        signal cVar1S10S83P017P037P019N003: std_logic_vector(   0 downto 0);
        signal cVar1S11S83P017P037P019N003: std_logic_vector(   0 downto 0);
        signal cVar1S12S83P017P037N019P001: std_logic_vector(   0 downto 0);
        signal cVar1S13S83P017P037N019P001: std_logic_vector(   0 downto 0);
        signal cVar1S14S83P017P037N019P001: std_logic_vector(   0 downto 0);
        signal cVar1S15S83P017P044P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S16S83P017P044P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S17S83P017N044P023P052: std_logic_vector(   0 downto 0);
        signal cVar1S18S83P017N044P023P052: std_logic_vector(   0 downto 0);
        signal cVar1S19S83P017N044P023N052: std_logic_vector(   0 downto 0);
        signal cVar1S20S83P017N044P023N052: std_logic_vector(   0 downto 0);
        signal cVar1S21S83P017N044P023N052: std_logic_vector(   0 downto 0);
        signal cVar1S22S83P017N044P023P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S83P017N044P023N065: std_logic_vector(   0 downto 0);
        signal cVar1S0S84P019P018P057P064: std_logic_vector(   0 downto 0);
        signal cVar1S1S84P019P018P057P064: std_logic_vector(   0 downto 0);
        signal cVar1S2S84P019P018P057P064: std_logic_vector(   0 downto 0);
        signal cVar1S3S84P019P018P057P064: std_logic_vector(   0 downto 0);
        signal cVar1S4S84P019P018P057P064: std_logic_vector(   0 downto 0);
        signal cVar1S5S84P019P018P057P003: std_logic_vector(   0 downto 0);
        signal cVar1S6S84P019P018P057N003: std_logic_vector(   0 downto 0);
        signal cVar1S7S84P019P018P057N003: std_logic_vector(   0 downto 0);
        signal cVar1S8S84P019P018P057N003: std_logic_vector(   0 downto 0);
        signal cVar1S9S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S10S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S11S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S12S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S84P019P018P033P014: std_logic_vector(   0 downto 0);
        signal cVar1S16S84P019P018P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S17S84P019P018P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S18S84P019P018P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S19S84P019P018P033N013: std_logic_vector(   0 downto 0);
        signal cVar1S20S84P019P018P033N013: std_logic_vector(   0 downto 0);
        signal cVar1S21S84N019P047P006P064: std_logic_vector(   0 downto 0);
        signal cVar1S22S84N019P047P006P064: std_logic_vector(   0 downto 0);
        signal cVar1S23S84N019P047N006P066: std_logic_vector(   0 downto 0);
        signal cVar1S24S84N019P047N006P066: std_logic_vector(   0 downto 0);
        signal cVar1S25S84N019P047N006P066: std_logic_vector(   0 downto 0);
        signal cVar1S26S84N019P047N006P066: std_logic_vector(   0 downto 0);
        signal cVar1S27S84N019P047N006P066: std_logic_vector(   0 downto 0);
        signal cVar1S28S84N019N047P043P044: std_logic_vector(   0 downto 0);
        signal cVar1S29S84N019N047P043P044: std_logic_vector(   0 downto 0);
        signal cVar1S30S84N019N047P043P044: std_logic_vector(   0 downto 0);
        signal cVar1S31S84N019N047P043P044: std_logic_vector(   0 downto 0);
        signal cVar1S32S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S33S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S34S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S35S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S36S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S37S84N019N047N043P024: std_logic_vector(   0 downto 0);
        signal cVar1S0S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S1S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S3S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S4S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S5S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S6S85P019P051P067P007: std_logic_vector(   0 downto 0);
        signal cVar1S7S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S8S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S9S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S10S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S11S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S12S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S13S85P019P051N067P001: std_logic_vector(   0 downto 0);
        signal cVar1S14S85P019P051P008P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S85P019P051P008N027: std_logic_vector(   0 downto 0);
        signal cVar1S16S85P019P051P008N027: std_logic_vector(   0 downto 0);
        signal cVar1S17S85P019P051N008P057: std_logic_vector(   0 downto 0);
        signal cVar1S18S85P019P051N008P057: std_logic_vector(   0 downto 0);
        signal cVar1S19S85P019P051N008P057: std_logic_vector(   0 downto 0);
        signal cVar1S20S85P019P051N008P057: std_logic_vector(   0 downto 0);
        signal cVar1S21S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S22S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S23S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S24S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S25S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S26S85P019P018P014P033: std_logic_vector(   0 downto 0);
        signal cVar1S27S85P019P018P014P023: std_logic_vector(   0 downto 0);
        signal cVar1S28S85P019P018P014N023: std_logic_vector(   0 downto 0);
        signal cVar1S29S85P019P018P014N023: std_logic_vector(   0 downto 0);
        signal cVar1S30S85P019P018P014N023: std_logic_vector(   0 downto 0);
        signal cVar1S31S85P019P018P014N023: std_logic_vector(   0 downto 0);
        signal cVar1S32S85P019N018P033P012: std_logic_vector(   0 downto 0);
        signal cVar1S33S85P019N018P033P012: std_logic_vector(   0 downto 0);
        signal cVar1S34S85P019N018P033N012: std_logic_vector(   0 downto 0);
        signal cVar1S35S85P019N018P033N012: std_logic_vector(   0 downto 0);
        signal cVar1S36S85P019N018N033P010: std_logic_vector(   0 downto 0);
        signal cVar1S37S85P019N018N033P010: std_logic_vector(   0 downto 0);
        signal cVar1S38S85P019N018N033P010: std_logic_vector(   0 downto 0);
        signal cVar1S39S85P019N018N033N010: std_logic_vector(   0 downto 0);
        signal cVar1S40S85P019N018N033N010: std_logic_vector(   0 downto 0);
        signal cVar1S41S85P019N018N033N010: std_logic_vector(   0 downto 0);
        signal cVar1S0S86P019P018P036P014: std_logic_vector(   0 downto 0);
        signal cVar1S1S86P019P018P036P014: std_logic_vector(   0 downto 0);
        signal cVar1S2S86P019P018P036P014: std_logic_vector(   0 downto 0);
        signal cVar1S3S86P019P018P036N014: std_logic_vector(   0 downto 0);
        signal cVar1S4S86P019P018P036N014: std_logic_vector(   0 downto 0);
        signal cVar1S5S86P019P018P036N014: std_logic_vector(   0 downto 0);
        signal cVar1S6S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S7S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S8S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S9S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S10S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S11S86P019P018N036P069: std_logic_vector(   0 downto 0);
        signal cVar1S12S86P019P018P055P030: std_logic_vector(   0 downto 0);
        signal cVar1S13S86P019P018P055P030: std_logic_vector(   0 downto 0);
        signal cVar1S14S86P019P018P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S15S86P019P018P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S16S86P019P018P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S17S86P019P018N055P046: std_logic_vector(   0 downto 0);
        signal cVar1S18S86P019P018N055P046: std_logic_vector(   0 downto 0);
        signal cVar1S19S86P019P018N055P046: std_logic_vector(   0 downto 0);
        signal cVar1S20S86P019P018N055P046: std_logic_vector(   0 downto 0);
        signal cVar1S21S86N019P067P002P031: std_logic_vector(   0 downto 0);
        signal cVar1S22S86N019P067P002P031: std_logic_vector(   0 downto 0);
        signal cVar1S23S86N019P067P002P031: std_logic_vector(   0 downto 0);
        signal cVar1S24S86N019P067P002P031: std_logic_vector(   0 downto 0);
        signal cVar1S25S86N019P067P002P031: std_logic_vector(   0 downto 0);
        signal cVar1S26S86N019P067P002P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S27S86N019P067P002N064: std_logic_vector(   0 downto 0);
        signal cVar1S28S86N019N067P017P011: std_logic_vector(   0 downto 0);
        signal cVar1S29S86N019N067P017P011: std_logic_vector(   0 downto 0);
        signal cVar1S30S86N019N067P017N011: std_logic_vector(   0 downto 0);
        signal cVar1S31S86N019N067P017N011: std_logic_vector(   0 downto 0);
        signal cVar1S32S86N019N067P017N011: std_logic_vector(   0 downto 0);
        signal cVar1S33S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S34S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S35S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S36S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S37S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S38S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S39S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S40S86N019N067N017P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S87P017P002P038P066: std_logic_vector(   0 downto 0);
        signal cVar1S1S87P017P002P038P066: std_logic_vector(   0 downto 0);
        signal cVar1S2S87P017P002P038P066: std_logic_vector(   0 downto 0);
        signal cVar1S3S87P017P002P038P066: std_logic_vector(   0 downto 0);
        signal cVar1S4S87P017P002P038N066: std_logic_vector(   0 downto 0);
        signal cVar1S5S87P017P002P038N066: std_logic_vector(   0 downto 0);
        signal cVar1S6S87P017P002P038N066: std_logic_vector(   0 downto 0);
        signal cVar1S7S87P017P002P038P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S87P017P002P038N004: std_logic_vector(   0 downto 0);
        signal cVar1S9S87P017P002P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S87P017P002N040P013: std_logic_vector(   0 downto 0);
        signal cVar1S11S87P017P002N040P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S87P017P002N040N013: std_logic_vector(   0 downto 0);
        signal cVar1S13S87P017P002N040N013: std_logic_vector(   0 downto 0);
        signal cVar1S14S87P017P002N040N013: std_logic_vector(   0 downto 0);
        signal cVar1S15S87N017P019P052P003: std_logic_vector(   0 downto 0);
        signal cVar1S16S87N017P019P052P003: std_logic_vector(   0 downto 0);
        signal cVar1S17S87N017P019P052P003: std_logic_vector(   0 downto 0);
        signal cVar1S18S87N017P019P052N003: std_logic_vector(   0 downto 0);
        signal cVar1S19S87N017P019P052N003: std_logic_vector(   0 downto 0);
        signal cVar1S20S87N017P019P052N003: std_logic_vector(   0 downto 0);
        signal cVar1S21S87N017P019P052P009: std_logic_vector(   0 downto 0);
        signal cVar1S22S87N017P019P052P009: std_logic_vector(   0 downto 0);
        signal cVar1S23S87N017P019P052N009: std_logic_vector(   0 downto 0);
        signal cVar1S24S87N017P019P052N009: std_logic_vector(   0 downto 0);
        signal cVar1S25S87N017P019P052N009: std_logic_vector(   0 downto 0);
        signal cVar1S26S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S27S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S28S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S29S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S30S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S31S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S32S87N017N019P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S33S87N017N019P069P064: std_logic_vector(   0 downto 0);
        signal cVar1S34S87N017N019P069P064: std_logic_vector(   0 downto 0);
        signal cVar1S35S87N017N019P069P064: std_logic_vector(   0 downto 0);
        signal cVar1S36S87N017N019P069P064: std_logic_vector(   0 downto 0);
        signal cVar1S37S87N017N019P069N064: std_logic_vector(   0 downto 0);
        signal cVar1S38S87N017N019P069N064: std_logic_vector(   0 downto 0);
        signal cVar1S39S87N017N019P069N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S1S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S3S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S4S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S5S88P014P016P018P012: std_logic_vector(   0 downto 0);
        signal cVar1S6S88P014P016P018P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S88P014P016P018P033: std_logic_vector(   0 downto 0);
        signal cVar1S8S88P014P016P018P033: std_logic_vector(   0 downto 0);
        signal cVar1S9S88P014P016P018N033: std_logic_vector(   0 downto 0);
        signal cVar1S10S88P014P016P018N033: std_logic_vector(   0 downto 0);
        signal cVar1S11S88P014P016P018N033: std_logic_vector(   0 downto 0);
        signal cVar1S12S88P014P016P018N033: std_logic_vector(   0 downto 0);
        signal cVar1S13S88P014N016P021P040: std_logic_vector(   0 downto 0);
        signal cVar1S14S88P014N016P021P040: std_logic_vector(   0 downto 0);
        signal cVar1S15S88P014N016P021P040: std_logic_vector(   0 downto 0);
        signal cVar1S16S88P014N016P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S17S88P014N016P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S18S88P014N016N021P054: std_logic_vector(   0 downto 0);
        signal cVar1S19S88P014N016N021P054: std_logic_vector(   0 downto 0);
        signal cVar1S20S88P014N016N021P054: std_logic_vector(   0 downto 0);
        signal cVar1S21S88P014N016N021N054: std_logic_vector(   0 downto 0);
        signal cVar1S22S88P014P021P003P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S88P014P021P003N019: std_logic_vector(   0 downto 0);
        signal cVar1S24S88P014P021N003P023: std_logic_vector(   0 downto 0);
        signal cVar1S25S88P014P021N003P023: std_logic_vector(   0 downto 0);
        signal cVar1S26S88P014P021N003P023: std_logic_vector(   0 downto 0);
        signal cVar1S27S88P014P021N003N023: std_logic_vector(   0 downto 0);
        signal cVar1S28S88P014P021N003N023: std_logic_vector(   0 downto 0);
        signal cVar1S29S88P014P021N003N023: std_logic_vector(   0 downto 0);
        signal cVar1S30S88P014P021P026P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S88P014P021P026P037: std_logic_vector(   0 downto 0);
        signal cVar1S32S88P014P021P026N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S89P014P017P015P037: std_logic_vector(   0 downto 0);
        signal cVar1S1S89P014P017P015P037: std_logic_vector(   0 downto 0);
        signal cVar1S2S89P014P017P015P037: std_logic_vector(   0 downto 0);
        signal cVar1S3S89P014P017P015N037: std_logic_vector(   0 downto 0);
        signal cVar1S4S89P014P017P015N037: std_logic_vector(   0 downto 0);
        signal cVar1S5S89P014P017P015N037: std_logic_vector(   0 downto 0);
        signal cVar1S6S89P014P017P015P030: std_logic_vector(   0 downto 0);
        signal cVar1S7S89P014P017P015P030: std_logic_vector(   0 downto 0);
        signal cVar1S8S89P014P017P015P030: std_logic_vector(   0 downto 0);
        signal cVar1S9S89P014P017P015N030: std_logic_vector(   0 downto 0);
        signal cVar1S10S89P014P017P015N030: std_logic_vector(   0 downto 0);
        signal cVar1S11S89P014N017P044P015: std_logic_vector(   0 downto 0);
        signal cVar1S12S89P014N017P044P015: std_logic_vector(   0 downto 0);
        signal cVar1S13S89P014N017P044P015: std_logic_vector(   0 downto 0);
        signal cVar1S14S89P014N017P044N015: std_logic_vector(   0 downto 0);
        signal cVar1S15S89P014N017P044N015: std_logic_vector(   0 downto 0);
        signal cVar1S16S89P014N017P044N015: std_logic_vector(   0 downto 0);
        signal cVar1S17S89P014N017N044P027: std_logic_vector(   0 downto 0);
        signal cVar1S18S89P014N017N044P027: std_logic_vector(   0 downto 0);
        signal cVar1S19S89P014N017N044N027: std_logic_vector(   0 downto 0);
        signal cVar1S20S89P014N017N044N027: std_logic_vector(   0 downto 0);
        signal cVar1S21S89P014P021P012P040: std_logic_vector(   0 downto 0);
        signal cVar1S22S89P014P021P012P040: std_logic_vector(   0 downto 0);
        signal cVar1S23S89P014P021P012P040: std_logic_vector(   0 downto 0);
        signal cVar1S24S89P014P021P012P040: std_logic_vector(   0 downto 0);
        signal cVar1S25S89P014P021P012P040: std_logic_vector(   0 downto 0);
        signal cVar1S26S89P014P021P012P039: std_logic_vector(   0 downto 0);
        signal cVar1S27S89P014P021P012P039: std_logic_vector(   0 downto 0);
        signal cVar1S28S89P014P021P012P039: std_logic_vector(   0 downto 0);
        signal cVar1S29S89P014P021P012P039: std_logic_vector(   0 downto 0);
        signal cVar1S30S89P014P021P026P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S89P014P021P026P037: std_logic_vector(   0 downto 0);
        signal cVar1S32S89P014P021P026N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S1S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S2S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S3S90P017P014P019N042: std_logic_vector(   0 downto 0);
        signal cVar1S4S90P017P014P019N042: std_logic_vector(   0 downto 0);
        signal cVar1S5S90P017P014P019N042: std_logic_vector(   0 downto 0);
        signal cVar1S6S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S7S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S8S90P017P014P019P042: std_logic_vector(   0 downto 0);
        signal cVar1S9S90P017P014P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S90P017P014P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S90P017P014P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S90P017P014P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S90P017P014P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S90P017P014P047P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S90N017P068P004P025: std_logic_vector(   0 downto 0);
        signal cVar1S16S90N017P068P004N025: std_logic_vector(   0 downto 0);
        signal cVar1S17S90N017P068P004N025: std_logic_vector(   0 downto 0);
        signal cVar1S18S90N017P068P004N025: std_logic_vector(   0 downto 0);
        signal cVar1S19S90N017P068N004P028: std_logic_vector(   0 downto 0);
        signal cVar1S20S90N017P068N004N028: std_logic_vector(   0 downto 0);
        signal cVar1S21S90N017P068N004N028: std_logic_vector(   0 downto 0);
        signal cVar1S22S90N017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S23S90N017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S24S90N017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S25S90N017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S26S90N017P068P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S27S90N017P068P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S28S90N017P068P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S29S90N017P068P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S0S91P017P068P010P004: std_logic_vector(   0 downto 0);
        signal cVar1S1S91P017P068P010P004: std_logic_vector(   0 downto 0);
        signal cVar1S2S91P017P068P010P004: std_logic_vector(   0 downto 0);
        signal cVar1S3S91P017P068P010N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S91P017P068P010N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S91P017P068P010N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S91P017P068P010P021: std_logic_vector(   0 downto 0);
        signal cVar1S7S91P017P068P010P021: std_logic_vector(   0 downto 0);
        signal cVar1S8S91P017P068P010P021: std_logic_vector(   0 downto 0);
        signal cVar1S9S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S10S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S15S91P017P068P064P062: std_logic_vector(   0 downto 0);
        signal cVar1S16S91P017P068P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S17S91P017P068P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S18S91P017P068P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S19S91P017P068P064N019: std_logic_vector(   0 downto 0);
        signal cVar1S20S91P017P044P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S21S91P017P044P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S22S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S23S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S24S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S25S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S26S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S27S91P017N044P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S28S91P017N044P023P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S29S91P017N044P023N065: std_logic_vector(   0 downto 0);
        signal cVar1S0S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S1S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S6S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S7S92P017P059P061P013: std_logic_vector(   0 downto 0);
        signal cVar1S8S92P017P059P061P066: std_logic_vector(   0 downto 0);
        signal cVar1S9S92P017P059P061P066: std_logic_vector(   0 downto 0);
        signal cVar1S10S92P017P059P061N066: std_logic_vector(   0 downto 0);
        signal cVar1S11S92P017P059P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S12S92P017P059P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S92P017P059P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S14S92P017P059N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S15S92P017P059N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S92P017P059N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S92P017P059N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S92P017P059N030P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S92N017P006P027P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S92N017P006P027N048: std_logic_vector(   0 downto 0);
        signal cVar1S21S92N017P006P027N048: std_logic_vector(   0 downto 0);
        signal cVar1S22S92N017P006N027P015: std_logic_vector(   0 downto 0);
        signal cVar1S23S92N017P006N027P015: std_logic_vector(   0 downto 0);
        signal cVar1S24S92N017P006N027N015: std_logic_vector(   0 downto 0);
        signal cVar1S25S92N017P006N027N015: std_logic_vector(   0 downto 0);
        signal cVar1S26S92N017N006P030P028: std_logic_vector(   0 downto 0);
        signal cVar1S27S92N017N006P030P028: std_logic_vector(   0 downto 0);
        signal cVar1S28S92N017N006P030P028: std_logic_vector(   0 downto 0);
        signal cVar1S29S92N017N006P030P028: std_logic_vector(   0 downto 0);
        signal cVar1S30S92N017N006P030P028: std_logic_vector(   0 downto 0);
        signal cVar1S31S92N017N006N030P014: std_logic_vector(   0 downto 0);
        signal cVar1S32S92N017N006N030P014: std_logic_vector(   0 downto 0);
        signal cVar1S33S92N017N006N030P014: std_logic_vector(   0 downto 0);
        signal cVar1S34S92N017N006N030N014: std_logic_vector(   0 downto 0);
        signal cVar1S35S92N017N006N030N014: std_logic_vector(   0 downto 0);
        signal cVar1S0S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S3S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S4S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S5S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S6S93P017P030P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S7S93P017P030P014P021: std_logic_vector(   0 downto 0);
        signal cVar1S8S93P017P030P014P021: std_logic_vector(   0 downto 0);
        signal cVar1S9S93P017P030P014P021: std_logic_vector(   0 downto 0);
        signal cVar1S10S93P017P030P014P021: std_logic_vector(   0 downto 0);
        signal cVar1S11S93P017P030P014P021: std_logic_vector(   0 downto 0);
        signal cVar1S12S93P017P030P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S93P017P030P061N013: std_logic_vector(   0 downto 0);
        signal cVar1S14S93P017P030P061N013: std_logic_vector(   0 downto 0);
        signal cVar1S15S93P017P030N061P032: std_logic_vector(   0 downto 0);
        signal cVar1S16S93P017P030N061P032: std_logic_vector(   0 downto 0);
        signal cVar1S17S93P017P030N061P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S20S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S21S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S22S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S23S93P017P013P003P008: std_logic_vector(   0 downto 0);
        signal cVar1S24S93P017P013P003P053: std_logic_vector(   0 downto 0);
        signal cVar1S25S93P017P013P003P053: std_logic_vector(   0 downto 0);
        signal cVar1S26S93P017N013P003P068: std_logic_vector(   0 downto 0);
        signal cVar1S27S93P017N013P003P068: std_logic_vector(   0 downto 0);
        signal cVar1S28S93P017N013P003P068: std_logic_vector(   0 downto 0);
        signal cVar1S29S93P017N013P003N068: std_logic_vector(   0 downto 0);
        signal cVar1S30S93P017N013P003N068: std_logic_vector(   0 downto 0);
        signal cVar1S31S93P017N013N003P002: std_logic_vector(   0 downto 0);
        signal cVar1S32S93P017N013N003P002: std_logic_vector(   0 downto 0);
        signal cVar1S33S93P017N013N003P002: std_logic_vector(   0 downto 0);
        signal cVar1S34S93P017N013N003P002: std_logic_vector(   0 downto 0);
        signal cVar1S35S93P017N013N003P002: std_logic_vector(   0 downto 0);
        signal cVar1S0S94P013P032P033P007: std_logic_vector(   0 downto 0);
        signal cVar1S1S94P013P032P033P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S94P013P032P033P007: std_logic_vector(   0 downto 0);
        signal cVar1S3S94P013P032P033P007: std_logic_vector(   0 downto 0);
        signal cVar1S4S94P013P032N033P031: std_logic_vector(   0 downto 0);
        signal cVar1S5S94P013P032N033P031: std_logic_vector(   0 downto 0);
        signal cVar1S6S94P013P032N033N031: std_logic_vector(   0 downto 0);
        signal cVar1S7S94P013P032N033N031: std_logic_vector(   0 downto 0);
        signal cVar1S8S94P013P032N033N031: std_logic_vector(   0 downto 0);
        signal cVar1S9S94P013P032P061P067: std_logic_vector(   0 downto 0);
        signal cVar1S10S94P013P032P061P067: std_logic_vector(   0 downto 0);
        signal cVar1S11S94P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S12S94P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S13S94P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S14S94P013P032N061P063: std_logic_vector(   0 downto 0);
        signal cVar1S15S94P013P032N061N063: std_logic_vector(   0 downto 0);
        signal cVar1S16S94P013P032N061N063: std_logic_vector(   0 downto 0);
        signal cVar1S17S94N013P017P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S18S94N013P017P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S19S94N013P017P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S20S94N013P017P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S94N013P017P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S22S94N013P017P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S23S94N013P017P068P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S94N013P017P068P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S94N013P017P068P003: std_logic_vector(   0 downto 0);
        signal cVar1S26S94N013P017P068N003: std_logic_vector(   0 downto 0);
        signal cVar1S27S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S28S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S29S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S30S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S31S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S32S94N013N017P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S33S94N013N017N015P019: std_logic_vector(   0 downto 0);
        signal cVar1S34S94N013N017N015P019: std_logic_vector(   0 downto 0);
        signal cVar1S35S94N013N017N015P019: std_logic_vector(   0 downto 0);
        signal cVar1S36S94N013N017N015N019: std_logic_vector(   0 downto 0);
        signal cVar1S37S94N013N017N015N019: std_logic_vector(   0 downto 0);
        signal cVar1S0S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S1S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S2S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S4S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S5S95P013P032P011P003: std_logic_vector(   0 downto 0);
        signal cVar1S6S95P013P032P011P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S95P013P032P011P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S95P013P032P011P036: std_logic_vector(   0 downto 0);
        signal cVar1S9S95P013P032P011N036: std_logic_vector(   0 downto 0);
        signal cVar1S10S95P013P032P011N036: std_logic_vector(   0 downto 0);
        signal cVar1S11S95P013P032P011N036: std_logic_vector(   0 downto 0);
        signal cVar1S12S95P013P032P011N036: std_logic_vector(   0 downto 0);
        signal cVar1S13S95P013P032P061P067nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S95P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S15S95P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S16S95P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S17S95P013P032P061N067: std_logic_vector(   0 downto 0);
        signal cVar1S18S95P013P032N061P063: std_logic_vector(   0 downto 0);
        signal cVar1S19S95P013P032N061N063: std_logic_vector(   0 downto 0);
        signal cVar1S20S95P013P032N061N063: std_logic_vector(   0 downto 0);
        signal cVar1S21S95N013P019P041P004: std_logic_vector(   0 downto 0);
        signal cVar1S22S95N013P019P041P004: std_logic_vector(   0 downto 0);
        signal cVar1S23S95N013P019P041N004: std_logic_vector(   0 downto 0);
        signal cVar1S24S95N013P019P041N004: std_logic_vector(   0 downto 0);
        signal cVar1S25S95N013P019P041N004: std_logic_vector(   0 downto 0);
        signal cVar1S26S95N013P019N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S27S95N013P019N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S28S95N013P019N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S29S95N013P019N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S30S95N013P019P017P066: std_logic_vector(   0 downto 0);
        signal cVar1S31S95N013P019P017P066: std_logic_vector(   0 downto 0);
        signal cVar1S32S95N013P019P017P066: std_logic_vector(   0 downto 0);
        signal cVar1S33S95N013P019P017P066: std_logic_vector(   0 downto 0);
        signal cVar1S34S95N013P019P017P066: std_logic_vector(   0 downto 0);
        signal cVar1S35S95N013P019N017P048: std_logic_vector(   0 downto 0);
        signal cVar1S36S95N013P019N017P048: std_logic_vector(   0 downto 0);
        signal cVar1S37S95N013P019N017P048: std_logic_vector(   0 downto 0);
        signal cVar1S38S95N013P019N017N048: std_logic_vector(   0 downto 0);
        signal cVar1S39S95N013P019N017N048: std_logic_vector(   0 downto 0);
        signal cVar1S40S95N013P019N017N048: std_logic_vector(   0 downto 0);
        signal cVar1S0S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S1S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S2S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S5S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S6S96P019P012P058P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S8S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S9S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S10S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S12S96P019P012P058P068: std_logic_vector(   0 downto 0);
        signal cVar1S13S96P019P012P043P056: std_logic_vector(   0 downto 0);
        signal cVar1S14S96P019P012P043P056: std_logic_vector(   0 downto 0);
        signal cVar1S15S96P019P012P043P056: std_logic_vector(   0 downto 0);
        signal cVar1S16S96P019P012P043N056: std_logic_vector(   0 downto 0);
        signal cVar1S17S96P019P012P043N056: std_logic_vector(   0 downto 0);
        signal cVar1S18S96P019P012P043N056: std_logic_vector(   0 downto 0);
        signal cVar1S19S96P019P003P057P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S96P019P003P057P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S96P019P003N057P068: std_logic_vector(   0 downto 0);
        signal cVar1S22S96P019P003N057P068: std_logic_vector(   0 downto 0);
        signal cVar1S23S96P019P003N057N068: std_logic_vector(   0 downto 0);
        signal cVar1S24S96P019P003N057N068: std_logic_vector(   0 downto 0);
        signal cVar1S25S96P019P003N057N068: std_logic_vector(   0 downto 0);
        signal cVar1S26S96P019N003P057P025: std_logic_vector(   0 downto 0);
        signal cVar1S27S96P019N003P057P025: std_logic_vector(   0 downto 0);
        signal cVar1S28S96P019N003P057N025: std_logic_vector(   0 downto 0);
        signal cVar1S29S96P019N003P057N025: std_logic_vector(   0 downto 0);
        signal cVar1S30S96P019N003P057N025: std_logic_vector(   0 downto 0);
        signal cVar1S31S96P019N003P057N025: std_logic_vector(   0 downto 0);
        signal cVar1S32S96P019N003P057P066: std_logic_vector(   0 downto 0);
        signal cVar1S33S96P019N003P057P066: std_logic_vector(   0 downto 0);
        signal cVar1S34S96P019N003P057P066: std_logic_vector(   0 downto 0);
        signal cVar1S35S96P019N003P057P066: std_logic_vector(   0 downto 0);
        signal cVar1S36S96P019N003P057P066: std_logic_vector(   0 downto 0);
        signal cVar1S0S97P019P057P069P007: std_logic_vector(   0 downto 0);
        signal cVar1S1S97P019P057P069P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S97P019P057P069N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S97P019P057P069N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S97P019P057P069N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S97P019P057N069P038: std_logic_vector(   0 downto 0);
        signal cVar1S6S97P019P057N069P038: std_logic_vector(   0 downto 0);
        signal cVar1S7S97P019P057N069P038: std_logic_vector(   0 downto 0);
        signal cVar1S8S97P019P057N069P038: std_logic_vector(   0 downto 0);
        signal cVar1S9S97P019P057P003P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S97P019P057P003P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S97P019P057N003P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S97P019P057N003P011: std_logic_vector(   0 downto 0);
        signal cVar1S13S97P019P057N003N011: std_logic_vector(   0 downto 0);
        signal cVar1S14S97P019P057N003N011: std_logic_vector(   0 downto 0);
        signal cVar1S15S97P019P057N003N011: std_logic_vector(   0 downto 0);
        signal cVar1S16S97N019P060P021P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S97N019P060P021P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S97N019P060P021P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S97N019P060P021P055: std_logic_vector(   0 downto 0);
        signal cVar1S20S97N019P060P021P055: std_logic_vector(   0 downto 0);
        signal cVar1S21S97N019P060P021P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S97N019N060P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S23S97N019N060P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S24S97N019N060P068N036: std_logic_vector(   0 downto 0);
        signal cVar1S25S97N019N060P068N036: std_logic_vector(   0 downto 0);
        signal cVar1S26S97N019N060P068N036: std_logic_vector(   0 downto 0);
        signal cVar1S27S97N019N060P068P023: std_logic_vector(   0 downto 0);
        signal cVar1S28S97N019N060P068P023: std_logic_vector(   0 downto 0);
        signal cVar1S29S97N019N060P068P023: std_logic_vector(   0 downto 0);
        signal cVar1S30S97N019N060P068P023: std_logic_vector(   0 downto 0);
        signal cVar1S31S97N019N060P068P023: std_logic_vector(   0 downto 0);
        signal cVar1S0S98P019P060P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S1S98P019P060P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S2S98P019P060P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S98P019P060P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S4S98P019P060P033P003: std_logic_vector(   0 downto 0);
        signal cVar1S5S98P019P060N033P058: std_logic_vector(   0 downto 0);
        signal cVar1S6S98P019P060N033P058: std_logic_vector(   0 downto 0);
        signal cVar1S7S98P019P060N033P058: std_logic_vector(   0 downto 0);
        signal cVar1S8S98P019P060N033P058: std_logic_vector(   0 downto 0);
        signal cVar1S9S98P019P060P021P010: std_logic_vector(   0 downto 0);
        signal cVar1S10S98P019P060P021P010: std_logic_vector(   0 downto 0);
        signal cVar1S11S98P019P060P021P010: std_logic_vector(   0 downto 0);
        signal cVar1S12S98P019P060P021N010: std_logic_vector(   0 downto 0);
        signal cVar1S13S98P019P060P021N010: std_logic_vector(   0 downto 0);
        signal cVar1S14S98P019P060P021P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S98P019P069P013P017: std_logic_vector(   0 downto 0);
        signal cVar1S16S98P019P069P013P017: std_logic_vector(   0 downto 0);
        signal cVar1S17S98P019P069P013P017: std_logic_vector(   0 downto 0);
        signal cVar1S18S98P019P069P013P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S98P019P069N013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S98P019P069N013N022: std_logic_vector(   0 downto 0);
        signal cVar1S21S98P019P069N013N022: std_logic_vector(   0 downto 0);
        signal cVar1S22S98P019P069N013N022: std_logic_vector(   0 downto 0);
        signal cVar1S23S98P019N069P058P063: std_logic_vector(   0 downto 0);
        signal cVar1S24S98P019N069P058P063: std_logic_vector(   0 downto 0);
        signal cVar1S25S98P019N069P058N063: std_logic_vector(   0 downto 0);
        signal cVar1S26S98P019N069P058N063: std_logic_vector(   0 downto 0);
        signal cVar1S27S98P019N069N058P060: std_logic_vector(   0 downto 0);
        signal cVar1S28S98P019N069N058P060: std_logic_vector(   0 downto 0);
        signal cVar1S29S98P019N069N058P060: std_logic_vector(   0 downto 0);
        signal cVar1S30S98P019N069N058P060: std_logic_vector(   0 downto 0);
        signal cVar1S0S99P019P069P006P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S99P019P069P006N027: std_logic_vector(   0 downto 0);
        signal cVar1S2S99P019P069P006N027: std_logic_vector(   0 downto 0);
        signal cVar1S3S99P019P069P006N027: std_logic_vector(   0 downto 0);
        signal cVar1S4S99P019P069N006P047: std_logic_vector(   0 downto 0);
        signal cVar1S5S99P019P069N006P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S99P019P069N006P047: std_logic_vector(   0 downto 0);
        signal cVar1S7S99P019P069N006P047: std_logic_vector(   0 downto 0);
        signal cVar1S8S99P019N069P060P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S99P019N069P060P016: std_logic_vector(   0 downto 0);
        signal cVar1S10S99P019N069P060P016: std_logic_vector(   0 downto 0);
        signal cVar1S11S99P019N069P060P016: std_logic_vector(   0 downto 0);
        signal cVar1S12S99P019N069P060N016: std_logic_vector(   0 downto 0);
        signal cVar1S13S99P019N069P060N016: std_logic_vector(   0 downto 0);
        signal cVar1S14S99P019N069P060N016: std_logic_vector(   0 downto 0);
        signal cVar1S15S99P019N069P060N016: std_logic_vector(   0 downto 0);
        signal cVar1S16S99P019N069P060P058: std_logic_vector(   0 downto 0);
        signal cVar1S17S99P019N069P060N058: std_logic_vector(   0 downto 0);
        signal cVar1S18S99P019N069P060N058: std_logic_vector(   0 downto 0);
        signal cVar1S19S99N019P033P030P003: std_logic_vector(   0 downto 0);
        signal cVar1S20S99N019P033P030P003: std_logic_vector(   0 downto 0);
        signal cVar1S21S99N019P033P030P003: std_logic_vector(   0 downto 0);
        signal cVar1S22S99N019P033P030P003: std_logic_vector(   0 downto 0);
        signal cVar1S23S99N019P033P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S24S99N019P033P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S25S99N019P033P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S26S99N019P033P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S27S99N019N033P036P027: std_logic_vector(   0 downto 0);
        signal cVar1S28S99N019N033P036P027: std_logic_vector(   0 downto 0);
        signal cVar1S29S99N019N033P036P027: std_logic_vector(   0 downto 0);
        signal cVar1S30S99N019N033P036N027: std_logic_vector(   0 downto 0);
        signal cVar1S31S99N019N033P036N027: std_logic_vector(   0 downto 0);
        signal cVar1S32S99N019N033P036N027: std_logic_vector(   0 downto 0);
        signal cVar1S33S99N019N033P036P021: std_logic_vector(   0 downto 0);
        signal cVar1S34S99N019N033P036P021: std_logic_vector(   0 downto 0);
        signal cVar1S35S99N019N033P036P021: std_logic_vector(   0 downto 0);
        signal cVar1S36S99N019N033P036P021: std_logic_vector(   0 downto 0);
        signal cVar1S0S100P036P012P019P014: std_logic_vector(   0 downto 0);
        signal cVar1S1S100P036P012P019P014: std_logic_vector(   0 downto 0);
        signal cVar1S2S100P036P012P019P014: std_logic_vector(   0 downto 0);
        signal cVar1S3S100P036P012P019N014: std_logic_vector(   0 downto 0);
        signal cVar1S4S100P036P012P019N014: std_logic_vector(   0 downto 0);
        signal cVar1S5S100P036P012P019N014: std_logic_vector(   0 downto 0);
        signal cVar1S6S100P036P012P019N014: std_logic_vector(   0 downto 0);
        signal cVar1S7S100P036P012P019P016: std_logic_vector(   0 downto 0);
        signal cVar1S8S100P036P012P019P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S100P036P012P019P016: std_logic_vector(   0 downto 0);
        signal cVar1S10S100P036P012P019P016: std_logic_vector(   0 downto 0);
        signal cVar1S11S100P036P012P019N016: std_logic_vector(   0 downto 0);
        signal cVar1S12S100P036P012P019N016: std_logic_vector(   0 downto 0);
        signal cVar1S13S100P036P012P019N016: std_logic_vector(   0 downto 0);
        signal cVar1S14S100P036P012P018P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S100P036P012P018P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S100P036P012P018P066: std_logic_vector(   0 downto 0);
        signal cVar1S17S100P036P012P018P066: std_logic_vector(   0 downto 0);
        signal cVar1S18S100P036P012P018N066: std_logic_vector(   0 downto 0);
        signal cVar1S19S100P036P012P018N066: std_logic_vector(   0 downto 0);
        signal cVar1S20S100P036P012P018N066: std_logic_vector(   0 downto 0);
        signal cVar1S21S100P036P012N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S22S100P036P012N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S23S100P036P012N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S24S100P036P012N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S25S100P036P006P053P033: std_logic_vector(   0 downto 0);
        signal cVar1S26S100P036P006P053P033: std_logic_vector(   0 downto 0);
        signal cVar1S27S100P036P006P053P033: std_logic_vector(   0 downto 0);
        signal cVar1S28S100P036P006P053P033: std_logic_vector(   0 downto 0);
        signal cVar1S29S100P036N006P008P026: std_logic_vector(   0 downto 0);
        signal cVar1S30S100P036N006P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S31S100P036N006P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S32S100P036N006P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S33S100P036N006N008P047: std_logic_vector(   0 downto 0);
        signal cVar1S34S100P036N006N008P047: std_logic_vector(   0 downto 0);
        signal cVar1S35S100P036N006N008P047: std_logic_vector(   0 downto 0);
        signal cVar1S36S100P036N006N008P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S1S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S2S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S3S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S4S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S5S101P036P005P023P029: std_logic_vector(   0 downto 0);
        signal cVar1S6S101P036P005P023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S101P036P005P023N004: std_logic_vector(   0 downto 0);
        signal cVar1S8S101P036P005P069P013: std_logic_vector(   0 downto 0);
        signal cVar1S9S101P036P005P069P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S101P036P005N069P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S101P036P005N069N032: std_logic_vector(   0 downto 0);
        signal cVar1S12S101N036P014P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S13S101N036P014P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S14S101N036P014P061P069: std_logic_vector(   0 downto 0);
        signal cVar1S15S101N036P014P061N069: std_logic_vector(   0 downto 0);
        signal cVar1S16S101N036P014P061N069: std_logic_vector(   0 downto 0);
        signal cVar1S17S101N036P014P061N069: std_logic_vector(   0 downto 0);
        signal cVar1S18S101N036P014N061P069: std_logic_vector(   0 downto 0);
        signal cVar1S19S101N036P014N061P069: std_logic_vector(   0 downto 0);
        signal cVar1S20S101N036P014N061P069: std_logic_vector(   0 downto 0);
        signal cVar1S21S101N036P014N061P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S101N036P014N061P069: std_logic_vector(   0 downto 0);
        signal cVar1S23S101N036N014P012P023: std_logic_vector(   0 downto 0);
        signal cVar1S24S101N036N014P012P023: std_logic_vector(   0 downto 0);
        signal cVar1S25S101N036N014P012P023: std_logic_vector(   0 downto 0);
        signal cVar1S26S101N036N014P012P023: std_logic_vector(   0 downto 0);
        signal cVar1S27S101N036N014P012P023: std_logic_vector(   0 downto 0);
        signal cVar1S28S101N036N014N012P015: std_logic_vector(   0 downto 0);
        signal cVar1S29S101N036N014N012P015: std_logic_vector(   0 downto 0);
        signal cVar1S30S101N036N014N012P015: std_logic_vector(   0 downto 0);
        signal cVar1S31S101N036N014N012P015: std_logic_vector(   0 downto 0);
        signal cVar1S0S102P036P016P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S1S102P036P016P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S2S102P036P016P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S102P036P016P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S102P036P016N030P028: std_logic_vector(   0 downto 0);
        signal cVar1S5S102P036P016N030P028: std_logic_vector(   0 downto 0);
        signal cVar1S6S102P036P016N030P028: std_logic_vector(   0 downto 0);
        signal cVar1S7S102P036P016N030P028: std_logic_vector(   0 downto 0);
        signal cVar1S8S102P036P016N030N028: std_logic_vector(   0 downto 0);
        signal cVar1S9S102P036P016N030N028: std_logic_vector(   0 downto 0);
        signal cVar1S10S102P036P016N030N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S102P036P016P014P039: std_logic_vector(   0 downto 0);
        signal cVar1S12S102P036P016P014P039: std_logic_vector(   0 downto 0);
        signal cVar1S13S102P036P016P014P039: std_logic_vector(   0 downto 0);
        signal cVar1S14S102P036P016P014P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S102P036P016N014P037: std_logic_vector(   0 downto 0);
        signal cVar1S16S102P036P016N014P037: std_logic_vector(   0 downto 0);
        signal cVar1S17S102P036P016N014P037: std_logic_vector(   0 downto 0);
        signal cVar1S18S102P036P016N014N037: std_logic_vector(   0 downto 0);
        signal cVar1S19S102P036P016N014N037: std_logic_vector(   0 downto 0);
        signal cVar1S20S102P036P016N014N037: std_logic_vector(   0 downto 0);
        signal cVar1S21S102P036P000P069P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S102P036P000N069P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S102P036P000N069P013: std_logic_vector(   0 downto 0);
        signal cVar1S24S102P036N000P030P037: std_logic_vector(   0 downto 0);
        signal cVar1S25S102P036N000P030P037: std_logic_vector(   0 downto 0);
        signal cVar1S26S102P036N000P030P037: std_logic_vector(   0 downto 0);
        signal cVar1S27S102P036N000N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S28S102P036N000N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S29S102P036N000N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S30S102P036N000N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S31S102P036N000N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S0S103P036P001P023P043: std_logic_vector(   0 downto 0);
        signal cVar1S1S103P036P001P023P043: std_logic_vector(   0 downto 0);
        signal cVar1S2S103P036P001P023N043: std_logic_vector(   0 downto 0);
        signal cVar1S3S103P036P001P023N043: std_logic_vector(   0 downto 0);
        signal cVar1S4S103P036P001P023N043: std_logic_vector(   0 downto 0);
        signal cVar1S5S103P036P001P023P042: std_logic_vector(   0 downto 0);
        signal cVar1S6S103P036P001P034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S103P036P001N034P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S103P036P001N034N033: std_logic_vector(   0 downto 0);
        signal cVar1S9S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S10S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S11S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S12S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S13S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S14S103N036P011P040P010: std_logic_vector(   0 downto 0);
        signal cVar1S15S103N036P011P040P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S103N036P011P040N038: std_logic_vector(   0 downto 0);
        signal cVar1S17S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S20S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S21S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S22S103N036N011P016P055: std_logic_vector(   0 downto 0);
        signal cVar1S23S103N036N011N016P013: std_logic_vector(   0 downto 0);
        signal cVar1S24S103N036N011N016P013: std_logic_vector(   0 downto 0);
        signal cVar1S25S103N036N011N016P013: std_logic_vector(   0 downto 0);
        signal cVar1S26S103N036N011N016P013: std_logic_vector(   0 downto 0);
        signal cVar1S27S103N036N011N016N013: std_logic_vector(   0 downto 0);
        signal cVar1S28S103N036N011N016N013: std_logic_vector(   0 downto 0);
        signal cVar1S29S103N036N011N016N013: std_logic_vector(   0 downto 0);
        signal cVar1S0S104P036P051P026P048: std_logic_vector(   0 downto 0);
        signal cVar1S1S104P036P051P026P048: std_logic_vector(   0 downto 0);
        signal cVar1S2S104P036P051N026P028: std_logic_vector(   0 downto 0);
        signal cVar1S3S104P036P051N026P028: std_logic_vector(   0 downto 0);
        signal cVar1S4S104P036P051N026P028: std_logic_vector(   0 downto 0);
        signal cVar1S5S104P036P051N026N028: std_logic_vector(   0 downto 0);
        signal cVar1S6S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S7S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S8S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S9S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S10S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S11S104P036N051P053P009: std_logic_vector(   0 downto 0);
        signal cVar1S12S104P036N051P053P026: std_logic_vector(   0 downto 0);
        signal cVar1S13S104P036N051P053P026: std_logic_vector(   0 downto 0);
        signal cVar1S14S104P036N051P053P026: std_logic_vector(   0 downto 0);
        signal cVar1S15S104P036P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S104P036P043N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S104P036P043N022N024: std_logic_vector(   0 downto 0);
        signal cVar1S18S104P036P043N022N024: std_logic_vector(   0 downto 0);
        signal cVar1S19S104P036N043P045P038: std_logic_vector(   0 downto 0);
        signal cVar1S20S104P036N043P045P038: std_logic_vector(   0 downto 0);
        signal cVar1S21S104P036N043P045P038: std_logic_vector(   0 downto 0);
        signal cVar1S22S104P036N043P045P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S104P036N043P045N016: std_logic_vector(   0 downto 0);
        signal cVar1S0S105P013P061P016P030: std_logic_vector(   0 downto 0);
        signal cVar1S1S105P013P061P016N030: std_logic_vector(   0 downto 0);
        signal cVar1S2S105P013P061P016N030: std_logic_vector(   0 downto 0);
        signal cVar1S3S105P013P061P016P033: std_logic_vector(   0 downto 0);
        signal cVar1S4S105P013P061P016N033: std_logic_vector(   0 downto 0);
        signal cVar1S5S105P013P061P016N033: std_logic_vector(   0 downto 0);
        signal cVar1S6S105P013P061P016N033: std_logic_vector(   0 downto 0);
        signal cVar1S7S105P013N061P032P051: std_logic_vector(   0 downto 0);
        signal cVar1S8S105P013N061P032P051: std_logic_vector(   0 downto 0);
        signal cVar1S9S105P013N061P032P051: std_logic_vector(   0 downto 0);
        signal cVar1S10S105P013N061P032P051: std_logic_vector(   0 downto 0);
        signal cVar1S11S105P013N061P032N051: std_logic_vector(   0 downto 0);
        signal cVar1S12S105P013N061P032N051: std_logic_vector(   0 downto 0);
        signal cVar1S13S105P013N061P032N051: std_logic_vector(   0 downto 0);
        signal cVar1S14S105P013N061P032P063: std_logic_vector(   0 downto 0);
        signal cVar1S15S105P013N061P032N063: std_logic_vector(   0 downto 0);
        signal cVar1S16S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S17S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S18S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S19S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S20S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S21S105N013P036P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S22S105N013P036P002P068: std_logic_vector(   0 downto 0);
        signal cVar1S23S105N013N036P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S24S105N013N036P028P055: std_logic_vector(   0 downto 0);
        signal cVar1S25S105N013N036P028N055: std_logic_vector(   0 downto 0);
        signal cVar1S26S105N013N036P028N055: std_logic_vector(   0 downto 0);
        signal cVar1S27S105N013N036N028P026: std_logic_vector(   0 downto 0);
        signal cVar1S28S105N013N036N028N026: std_logic_vector(   0 downto 0);
        signal cVar1S29S105N013N036N028N026: std_logic_vector(   0 downto 0);
        signal cVar1S30S105N013N036N028N026: std_logic_vector(   0 downto 0);
        signal cVar1S0S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S1S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S2S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S3S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S4S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S5S106P036P064P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S6S106P036P064P002P012: std_logic_vector(   0 downto 0);
        signal cVar1S7S106P036P064P002P012: std_logic_vector(   0 downto 0);
        signal cVar1S8S106P036N064P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S9S106P036N064P062P015: std_logic_vector(   0 downto 0);
        signal cVar1S10S106P036N064P062N015: std_logic_vector(   0 downto 0);
        signal cVar1S11S106P036N064P062N015: std_logic_vector(   0 downto 0);
        signal cVar1S12S106P036N064P062N015: std_logic_vector(   0 downto 0);
        signal cVar1S13S106P036N064P062N015: std_logic_vector(   0 downto 0);
        signal cVar1S14S106P036N064P062P042: std_logic_vector(   0 downto 0);
        signal cVar1S15S106P036N064P062P042: std_logic_vector(   0 downto 0);
        signal cVar1S16S106P036N064P062P042: std_logic_vector(   0 downto 0);
        signal cVar1S17S106P036N064P062P042: std_logic_vector(   0 downto 0);
        signal cVar1S18S106P036P005P013P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S106P036P005P013P008: std_logic_vector(   0 downto 0);
        signal cVar1S20S106P036P005P013P008: std_logic_vector(   0 downto 0);
        signal cVar1S21S106P036P005P013P008: std_logic_vector(   0 downto 0);
        signal cVar1S22S106P036P005P013P008: std_logic_vector(   0 downto 0);
        signal cVar1S23S106P036P005N013P061: std_logic_vector(   0 downto 0);
        signal cVar1S24S106P036P005N013P061: std_logic_vector(   0 downto 0);
        signal cVar1S25S106P036P005N013P061: std_logic_vector(   0 downto 0);
        signal cVar1S26S106P036P005N013P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S106P036P005N013P061: std_logic_vector(   0 downto 0);
        signal cVar1S28S106P036P005P031P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S29S106P036P005P031N020: std_logic_vector(   0 downto 0);
        signal cVar1S30S106P036P005P031N020: std_logic_vector(   0 downto 0);
        signal cVar1S31S106P036P005P031N020: std_logic_vector(   0 downto 0);
        signal cVar1S0S107P036P005P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S1S107P036P005P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S2S107P036P005P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S3S107P036P005P019P047: std_logic_vector(   0 downto 0);
        signal cVar1S4S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S5S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S6S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S7S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S8S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S107P036P005N019P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S107P036P005P031P069: std_logic_vector(   0 downto 0);
        signal cVar1S11S107P036P005P031P069: std_logic_vector(   0 downto 0);
        signal cVar1S12S107P036P005P031N069: std_logic_vector(   0 downto 0);
        signal cVar1S13S107P036P005P031N069: std_logic_vector(   0 downto 0);
        signal cVar1S14S107N036P064P019P059: std_logic_vector(   0 downto 0);
        signal cVar1S15S107N036P064P019P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S107N036P064P019N059: std_logic_vector(   0 downto 0);
        signal cVar1S17S107N036P064P019N059: std_logic_vector(   0 downto 0);
        signal cVar1S18S107N036P064P019N059: std_logic_vector(   0 downto 0);
        signal cVar1S19S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S20S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S21S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S22S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S23S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S24S107N036P064N019P056: std_logic_vector(   0 downto 0);
        signal cVar1S25S107N036N064P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S26S107N036N064P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S27S107N036N064P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S28S107N036N064P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S29S107N036N064P051P057: std_logic_vector(   0 downto 0);
        signal cVar1S30S107N036N064N051P053: std_logic_vector(   0 downto 0);
        signal cVar1S31S107N036N064N051P053: std_logic_vector(   0 downto 0);
        signal cVar1S32S107N036N064N051P053: std_logic_vector(   0 downto 0);
        signal cVar1S33S107N036N064N051P053: std_logic_vector(   0 downto 0);
        signal cVar1S0S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S1S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S2S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S3S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S4S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S5S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S6S108P064P012P031P054: std_logic_vector(   0 downto 0);
        signal cVar1S7S108P064P012P031P005: std_logic_vector(   0 downto 0);
        signal cVar1S8S108P064P012P031P005: std_logic_vector(   0 downto 0);
        signal cVar1S9S108P064P012P031P005: std_logic_vector(   0 downto 0);
        signal cVar1S10S108P064P012P031P005: std_logic_vector(   0 downto 0);
        signal cVar1S11S108P064P012P030P032: std_logic_vector(   0 downto 0);
        signal cVar1S12S108P064P012P030P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S108P064P012P030P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S108P064P012P030P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S108P064P012P030P032: std_logic_vector(   0 downto 0);
        signal cVar1S16S108P064P012N030P054: std_logic_vector(   0 downto 0);
        signal cVar1S17S108P064P012N030P054: std_logic_vector(   0 downto 0);
        signal cVar1S18S108P064P012N030N054: std_logic_vector(   0 downto 0);
        signal cVar1S19S108P064P012N030N054: std_logic_vector(   0 downto 0);
        signal cVar1S20S108P064P068P062P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S108P064P068P062P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S108P064P068P062P066: std_logic_vector(   0 downto 0);
        signal cVar1S23S108P064P068P062N066: std_logic_vector(   0 downto 0);
        signal cVar1S24S108P064P068P062N066: std_logic_vector(   0 downto 0);
        signal cVar1S25S108P064P068P062N066: std_logic_vector(   0 downto 0);
        signal cVar1S26S108P064P068P062P045: std_logic_vector(   0 downto 0);
        signal cVar1S27S108P064P068P062P045: std_logic_vector(   0 downto 0);
        signal cVar1S28S108P064P068P062N045: std_logic_vector(   0 downto 0);
        signal cVar1S29S108P064P068P062N045: std_logic_vector(   0 downto 0);
        signal cVar1S30S108P064P068P012P035: std_logic_vector(   0 downto 0);
        signal cVar1S31S108P064P068P012P035: std_logic_vector(   0 downto 0);
        signal cVar1S32S108P064P068P012P035: std_logic_vector(   0 downto 0);
        signal cVar1S33S108P064P068P012N035: std_logic_vector(   0 downto 0);
        signal cVar1S34S108P064P068P012N035: std_logic_vector(   0 downto 0);
        signal cVar1S35S108P064P068N012P019: std_logic_vector(   0 downto 0);
        signal cVar1S36S108P064P068N012P019: std_logic_vector(   0 downto 0);
        signal cVar1S37S108P064P068N012N019: std_logic_vector(   0 downto 0);
        signal cVar1S38S108P064P068N012N019: std_logic_vector(   0 downto 0);
        signal cVar1S39S108P064P068N012N019: std_logic_vector(   0 downto 0);
        signal cVar1S0S109P064P068P055P056: std_logic_vector(   0 downto 0);
        signal cVar1S1S109P064P068P055P056: std_logic_vector(   0 downto 0);
        signal cVar1S2S109P064P068P055P056: std_logic_vector(   0 downto 0);
        signal cVar1S3S109P064P068P055P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S109P064P068P055P056: std_logic_vector(   0 downto 0);
        signal cVar1S5S109P064P068P055P060: std_logic_vector(   0 downto 0);
        signal cVar1S6S109P064P068P055P060: std_logic_vector(   0 downto 0);
        signal cVar1S7S109P064P068P055P060: std_logic_vector(   0 downto 0);
        signal cVar1S8S109P064P068P051P019: std_logic_vector(   0 downto 0);
        signal cVar1S9S109P064P068P051N019: std_logic_vector(   0 downto 0);
        signal cVar1S10S109P064P068P051N019: std_logic_vector(   0 downto 0);
        signal cVar1S11S109P064P068P051N019: std_logic_vector(   0 downto 0);
        signal cVar1S12S109P064P068P051P017nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S109N064P054P040P015: std_logic_vector(   0 downto 0);
        signal cVar1S14S109N064P054P040P015: std_logic_vector(   0 downto 0);
        signal cVar1S15S109N064P054P040P015: std_logic_vector(   0 downto 0);
        signal cVar1S16S109N064P054P040P015: std_logic_vector(   0 downto 0);
        signal cVar1S17S109N064P054P040N015: std_logic_vector(   0 downto 0);
        signal cVar1S18S109N064P054P040N015: std_logic_vector(   0 downto 0);
        signal cVar1S19S109N064P054P040N015: std_logic_vector(   0 downto 0);
        signal cVar1S20S109N064N054P022P043: std_logic_vector(   0 downto 0);
        signal cVar1S21S109N064N054P022P043: std_logic_vector(   0 downto 0);
        signal cVar1S22S109N064N054P022P043: std_logic_vector(   0 downto 0);
        signal cVar1S23S109N064N054P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S24S109N064N054P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S25S109N064N054P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S26S109N064N054N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S27S109N064N054N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S28S109N064N054N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S29S109N064N054N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S0S110P064P056P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S1S110P064P056P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S110P064P056P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S110P064P056P052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S110P064P056P052N009: std_logic_vector(   0 downto 0);
        signal cVar1S5S110P064P056P052N009: std_logic_vector(   0 downto 0);
        signal cVar1S6S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S7S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S8S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S9S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S10S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S11S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S12S110P064N056P026P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S110P064N056P026P050: std_logic_vector(   0 downto 0);
        signal cVar1S14S110P064N056P026P050: std_logic_vector(   0 downto 0);
        signal cVar1S15S110P064N056P026P050: std_logic_vector(   0 downto 0);
        signal cVar1S16S110P064N056P026N050: std_logic_vector(   0 downto 0);
        signal cVar1S17S110P064N056P026N050: std_logic_vector(   0 downto 0);
        signal cVar1S18S110P064N056P026N050: std_logic_vector(   0 downto 0);
        signal cVar1S19S110P064P013P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S20S110P064P013P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S21S110P064P013P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S22S110P064P013P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S23S110P064P013P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S24S110P064N013P033P022: std_logic_vector(   0 downto 0);
        signal cVar1S25S110P064N013P033P022: std_logic_vector(   0 downto 0);
        signal cVar1S26S110P064N013P033P050: std_logic_vector(   0 downto 0);
        signal cVar1S27S110P064N013P033P050: std_logic_vector(   0 downto 0);
        signal cVar1S0S111P064P033P041P018: std_logic_vector(   0 downto 0);
        signal cVar1S1S111P064P033P041P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S111P064P033P041P018: std_logic_vector(   0 downto 0);
        signal cVar1S3S111P064P033P041P018: std_logic_vector(   0 downto 0);
        signal cVar1S4S111P064P033P041P018: std_logic_vector(   0 downto 0);
        signal cVar1S5S111P064P033P041P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S111P064P033P048P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S111P064P033P048P050: std_logic_vector(   0 downto 0);
        signal cVar1S8S111P064P033P048P050: std_logic_vector(   0 downto 0);
        signal cVar1S9S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S111N064P016P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S15S111N064P016P047P034: std_logic_vector(   0 downto 0);
        signal cVar1S16S111N064P016P047N034: std_logic_vector(   0 downto 0);
        signal cVar1S17S111N064P016P047N034: std_logic_vector(   0 downto 0);
        signal cVar1S18S111N064N016P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S19S111N064N016P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S111N064N016P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S111N064N016P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S22S111N064N016P018N015: std_logic_vector(   0 downto 0);
        signal cVar1S23S111N064N016P018N015: std_logic_vector(   0 downto 0);
        signal cVar1S24S111N064N016P018N015: std_logic_vector(   0 downto 0);
        signal cVar1S25S111N064N016N018P059: std_logic_vector(   0 downto 0);
        signal cVar1S26S111N064N016N018N059: std_logic_vector(   0 downto 0);
        signal cVar1S27S111N064N016N018N059: std_logic_vector(   0 downto 0);
        signal cVar1S0S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S1S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S2S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S3S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S4S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S5S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S6S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S7S112P018P016P027P066: std_logic_vector(   0 downto 0);
        signal cVar1S8S112P018P016P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S9S112P018P016P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S10S112P018P016P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S11S112P018P016P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S12S112P018P016P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S13S112P018P016P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S14S112P018P016P059P065: std_logic_vector(   0 downto 0);
        signal cVar1S15S112P018P016P059P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S112P018P016P059P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S112P018P016N059P066: std_logic_vector(   0 downto 0);
        signal cVar1S18S112P018P016N059P066: std_logic_vector(   0 downto 0);
        signal cVar1S19S112P018P016N059P066: std_logic_vector(   0 downto 0);
        signal cVar1S20S112P018P016N059P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S112P018P016N059P066: std_logic_vector(   0 downto 0);
        signal cVar1S22S112N018P054P040P065: std_logic_vector(   0 downto 0);
        signal cVar1S23S112N018P054P040P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S112N018P054P040P065: std_logic_vector(   0 downto 0);
        signal cVar1S25S112N018P054P040P065: std_logic_vector(   0 downto 0);
        signal cVar1S26S112N018P054P040P065: std_logic_vector(   0 downto 0);
        signal cVar1S27S112N018N054P014P055: std_logic_vector(   0 downto 0);
        signal cVar1S28S112N018N054P014P055: std_logic_vector(   0 downto 0);
        signal cVar1S29S112N018N054P014N055: std_logic_vector(   0 downto 0);
        signal cVar1S30S112N018N054P014N055: std_logic_vector(   0 downto 0);
        signal cVar1S31S112N018N054P014N055: std_logic_vector(   0 downto 0);
        signal cVar1S32S112N018N054P014N055: std_logic_vector(   0 downto 0);
        signal cVar1S33S112N018N054P014P031: std_logic_vector(   0 downto 0);
        signal cVar1S34S112N018N054P014P031: std_logic_vector(   0 downto 0);
        signal cVar1S35S112N018N054P014P031: std_logic_vector(   0 downto 0);
        signal cVar1S36S112N018N054P014P031: std_logic_vector(   0 downto 0);
        signal cVar1S37S112N018N054P014P031: std_logic_vector(   0 downto 0);
        signal cVar1S0S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S1S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S2S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S5S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S6S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S113P014P018P056P011: std_logic_vector(   0 downto 0);
        signal cVar1S8S113P014P018P056P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S113P014P018P056P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S113P014P018P056N017: std_logic_vector(   0 downto 0);
        signal cVar1S11S113P014P018P056N017: std_logic_vector(   0 downto 0);
        signal cVar1S12S113P014P018P056N017: std_logic_vector(   0 downto 0);
        signal cVar1S13S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S14S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S15S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S16S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S17S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S18S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S19S113P014P018P067P050: std_logic_vector(   0 downto 0);
        signal cVar1S20S113P014P018N067P012: std_logic_vector(   0 downto 0);
        signal cVar1S21S113P014P018N067P012: std_logic_vector(   0 downto 0);
        signal cVar1S22S113P014P018N067P012: std_logic_vector(   0 downto 0);
        signal cVar1S23S113P014P018N067P012: std_logic_vector(   0 downto 0);
        signal cVar1S24S113P014P018N067N012: std_logic_vector(   0 downto 0);
        signal cVar1S25S113P014P018N067N012: std_logic_vector(   0 downto 0);
        signal cVar1S26S113P014P018N067N012: std_logic_vector(   0 downto 0);
        signal cVar1S27S113P014P018N067N012: std_logic_vector(   0 downto 0);
        signal cVar1S28S113P014P018P022P023: std_logic_vector(   0 downto 0);
        signal cVar1S29S113P014P018P022N023: std_logic_vector(   0 downto 0);
        signal cVar1S30S113P014P018P022N023: std_logic_vector(   0 downto 0);
        signal cVar1S31S113P014P018P022N023: std_logic_vector(   0 downto 0);
        signal cVar1S32S113P014P018P022N023: std_logic_vector(   0 downto 0);
        signal cVar1S33S113P014P018P022P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S34S113P014P018P022N037: std_logic_vector(   0 downto 0);
        signal cVar1S35S113P014N018P036P035: std_logic_vector(   0 downto 0);
        signal cVar1S36S113P014N018P036P035: std_logic_vector(   0 downto 0);
        signal cVar1S37S113P014N018P036P035: std_logic_vector(   0 downto 0);
        signal cVar1S38S113P014N018P036P035: std_logic_vector(   0 downto 0);
        signal cVar1S39S113P014N018P036N035: std_logic_vector(   0 downto 0);
        signal cVar1S40S113P014N018P036N035: std_logic_vector(   0 downto 0);
        signal cVar1S41S113P014N018P036N035: std_logic_vector(   0 downto 0);
        signal cVar1S42S113P014N018P036N035: std_logic_vector(   0 downto 0);
        signal cVar1S43S113P014N018P036P053: std_logic_vector(   0 downto 0);
        signal cVar1S44S113P014N018P036P053: std_logic_vector(   0 downto 0);
        signal cVar1S0S114P018P064P007P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S114P018P064P007N032: std_logic_vector(   0 downto 0);
        signal cVar1S2S114P018P064P007N032: std_logic_vector(   0 downto 0);
        signal cVar1S3S114P018P064P007N032: std_logic_vector(   0 downto 0);
        signal cVar1S4S114P018P064P007N032: std_logic_vector(   0 downto 0);
        signal cVar1S5S114P018P064P007P059: std_logic_vector(   0 downto 0);
        signal cVar1S6S114P018P064P007P059: std_logic_vector(   0 downto 0);
        signal cVar1S7S114P018P064P007P059: std_logic_vector(   0 downto 0);
        signal cVar1S8S114P018N064P050P034: std_logic_vector(   0 downto 0);
        signal cVar1S9S114P018N064P050P034: std_logic_vector(   0 downto 0);
        signal cVar1S10S114P018N064P050N034: std_logic_vector(   0 downto 0);
        signal cVar1S11S114P018N064P050N034: std_logic_vector(   0 downto 0);
        signal cVar1S12S114P018N064P050N034: std_logic_vector(   0 downto 0);
        signal cVar1S13S114P018N064P050N034: std_logic_vector(   0 downto 0);
        signal cVar1S14S114P018N064P050P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S114P018N064P050P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S114P018N064P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S17S114P018N064P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S18S114P018N064P050N008: std_logic_vector(   0 downto 0);
        signal cVar1S19S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S22S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S23S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S24S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S25S114N018P014P035P015: std_logic_vector(   0 downto 0);
        signal cVar1S26S114N018P014P035P024: std_logic_vector(   0 downto 0);
        signal cVar1S27S114N018P014P035P024: std_logic_vector(   0 downto 0);
        signal cVar1S28S114N018P014P035P024: std_logic_vector(   0 downto 0);
        signal cVar1S29S114N018N014P010P030: std_logic_vector(   0 downto 0);
        signal cVar1S30S114N018N014P010P030: std_logic_vector(   0 downto 0);
        signal cVar1S31S114N018N014P010P030: std_logic_vector(   0 downto 0);
        signal cVar1S32S114N018N014P010N030: std_logic_vector(   0 downto 0);
        signal cVar1S33S114N018N014P010N030: std_logic_vector(   0 downto 0);
        signal cVar1S34S114N018N014P010N030: std_logic_vector(   0 downto 0);
        signal cVar1S35S114N018N014N010P011: std_logic_vector(   0 downto 0);
        signal cVar1S36S114N018N014N010P011: std_logic_vector(   0 downto 0);
        signal cVar1S37S114N018N014N010N011: std_logic_vector(   0 downto 0);
        signal cVar1S38S114N018N014N010N011: std_logic_vector(   0 downto 0);
        signal cVar1S0S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S1S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S2S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S3S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S4S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S5S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S6S115P018P014P069P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S8S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S10S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S11S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S12S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S13S115P018P014N069P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S16S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S17S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S18S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S19S115P018P014P007P064: std_logic_vector(   0 downto 0);
        signal cVar1S20S115P018P014P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S115P018P014P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S115P018P014P007P037: std_logic_vector(   0 downto 0);
        signal cVar1S23S115P018P014P007N037: std_logic_vector(   0 downto 0);
        signal cVar1S24S115P018P014P007N037: std_logic_vector(   0 downto 0);
        signal cVar1S25S115P018P014P007N037: std_logic_vector(   0 downto 0);
        signal cVar1S26S115P018P062P066P042: std_logic_vector(   0 downto 0);
        signal cVar1S27S115P018P062P066P042: std_logic_vector(   0 downto 0);
        signal cVar1S28S115P018P062P066P042: std_logic_vector(   0 downto 0);
        signal cVar1S29S115P018P062P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S30S115P018P062P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S31S115P018P062P066N068: std_logic_vector(   0 downto 0);
        signal cVar1S32S115P018P062P066N068: std_logic_vector(   0 downto 0);
        signal cVar1S33S115P018N062P007P047: std_logic_vector(   0 downto 0);
        signal cVar1S34S115P018N062P007P047: std_logic_vector(   0 downto 0);
        signal cVar1S35S115P018N062P007N047: std_logic_vector(   0 downto 0);
        signal cVar1S36S115P018N062P007N047: std_logic_vector(   0 downto 0);
        signal cVar1S37S115P018N062P007N047: std_logic_vector(   0 downto 0);
        signal cVar1S38S115P018N062N007P034: std_logic_vector(   0 downto 0);
        signal cVar1S39S115P018N062N007P034: std_logic_vector(   0 downto 0);
        signal cVar1S40S115P018N062N007P034: std_logic_vector(   0 downto 0);
        signal cVar1S41S115P018N062N007N034: std_logic_vector(   0 downto 0);
        signal cVar1S42S115P018N062N007N034: std_logic_vector(   0 downto 0);
        signal cVar1S0S116P018P063P049P059: std_logic_vector(   0 downto 0);
        signal cVar1S1S116P018P063P049P059: std_logic_vector(   0 downto 0);
        signal cVar1S2S116P018P063P049P059: std_logic_vector(   0 downto 0);
        signal cVar1S3S116P018P063N049P066: std_logic_vector(   0 downto 0);
        signal cVar1S4S116P018P063N049P066: std_logic_vector(   0 downto 0);
        signal cVar1S5S116P018P063N049P066: std_logic_vector(   0 downto 0);
        signal cVar1S6S116P018P063N049N066: std_logic_vector(   0 downto 0);
        signal cVar1S7S116P018P063N049N066: std_logic_vector(   0 downto 0);
        signal cVar1S8S116P018P063N049N066: std_logic_vector(   0 downto 0);
        signal cVar1S9S116P018P063N049N066: std_logic_vector(   0 downto 0);
        signal cVar1S10S116P018P063P031P056: std_logic_vector(   0 downto 0);
        signal cVar1S11S116P018P063P031P056: std_logic_vector(   0 downto 0);
        signal cVar1S12S116P018P063P031N056: std_logic_vector(   0 downto 0);
        signal cVar1S13S116P018P063N031P033: std_logic_vector(   0 downto 0);
        signal cVar1S14S116P018P063N031P033: std_logic_vector(   0 downto 0);
        signal cVar1S15S116P018P063N031P033: std_logic_vector(   0 downto 0);
        signal cVar1S16S116P018P063N031P033: std_logic_vector(   0 downto 0);
        signal cVar1S17S116P018P063N031N033: std_logic_vector(   0 downto 0);
        signal cVar1S18S116P018P063N031N033: std_logic_vector(   0 downto 0);
        signal cVar1S19S116P018P063N031N033: std_logic_vector(   0 downto 0);
        signal cVar1S20S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S21S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S24S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S25S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S116N018P069P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S27S116N018P069N064P065: std_logic_vector(   0 downto 0);
        signal cVar1S28S116N018P069N064P065: std_logic_vector(   0 downto 0);
        signal cVar1S29S116N018P069N064P065: std_logic_vector(   0 downto 0);
        signal cVar1S30S116N018P069N064P065: std_logic_vector(   0 downto 0);
        signal cVar1S31S116N018P069N064P065: std_logic_vector(   0 downto 0);
        signal cVar1S32S116N018N069P056P012: std_logic_vector(   0 downto 0);
        signal cVar1S33S116N018N069P056P012: std_logic_vector(   0 downto 0);
        signal cVar1S34S116N018N069P056P012: std_logic_vector(   0 downto 0);
        signal cVar1S35S116N018N069P056N012: std_logic_vector(   0 downto 0);
        signal cVar1S36S116N018N069N056P013: std_logic_vector(   0 downto 0);
        signal cVar1S37S116N018N069N056P013: std_logic_vector(   0 downto 0);
        signal cVar1S38S116N018N069N056P013: std_logic_vector(   0 downto 0);
        signal cVar1S39S116N018N069N056P013: std_logic_vector(   0 downto 0);
        signal cVar1S40S116N018N069N056N013: std_logic_vector(   0 downto 0);
        signal cVar1S41S116N018N069N056N013: std_logic_vector(   0 downto 0);
        signal cVar1S0S117P066P069P063P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S117P066P069P063P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S117P066P069P063N067: std_logic_vector(   0 downto 0);
        signal cVar1S3S117P066P069P063N067: std_logic_vector(   0 downto 0);
        signal cVar1S4S117P066P069P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S5S117P066P069P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S6S117P066P069P063P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S117P066N069P068P047: std_logic_vector(   0 downto 0);
        signal cVar1S8S117P066N069P068P047: std_logic_vector(   0 downto 0);
        signal cVar1S9S117P066N069P068P047: std_logic_vector(   0 downto 0);
        signal cVar1S10S117P066N069P068N047: std_logic_vector(   0 downto 0);
        signal cVar1S11S117P066N069P068N047: std_logic_vector(   0 downto 0);
        signal cVar1S12S117P066N069P068N047: std_logic_vector(   0 downto 0);
        signal cVar1S13S117P066N069P068N047: std_logic_vector(   0 downto 0);
        signal cVar1S14S117P066N069P068P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S117P066N069P068P064: std_logic_vector(   0 downto 0);
        signal cVar1S16S117P066N069P068N064: std_logic_vector(   0 downto 0);
        signal cVar1S17S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S18S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S117P066P018P006P047: std_logic_vector(   0 downto 0);
        signal cVar1S23S117P066P018P006P024: std_logic_vector(   0 downto 0);
        signal cVar1S24S117P066P018P006P024: std_logic_vector(   0 downto 0);
        signal cVar1S25S117P066P018P006N024: std_logic_vector(   0 downto 0);
        signal cVar1S26S117P066P018P006N024: std_logic_vector(   0 downto 0);
        signal cVar1S27S117P066P018P049P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S117P066P018P049N051: std_logic_vector(   0 downto 0);
        signal cVar1S29S117P066P018P049N051: std_logic_vector(   0 downto 0);
        signal cVar1S30S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S31S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S32S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S33S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S34S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S35S117P066P018N049P067: std_logic_vector(   0 downto 0);
        signal cVar1S0S118P035P033P002P048: std_logic_vector(   0 downto 0);
        signal cVar1S1S118P035P033P002N048: std_logic_vector(   0 downto 0);
        signal cVar1S2S118P035P033P002N048: std_logic_vector(   0 downto 0);
        signal cVar1S3S118P035P033P002N048: std_logic_vector(   0 downto 0);
        signal cVar1S4S118P035P033P002P018: std_logic_vector(   0 downto 0);
        signal cVar1S5S118P035P033P002N018: std_logic_vector(   0 downto 0);
        signal cVar1S6S118P035P033P002N018: std_logic_vector(   0 downto 0);
        signal cVar1S7S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S8S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S9S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S10S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S11S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S12S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S13S118P035N033P019P069: std_logic_vector(   0 downto 0);
        signal cVar1S14S118P035N033P019P018: std_logic_vector(   0 downto 0);
        signal cVar1S15S118P035N033P019P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S118P035N033P019P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S118P035N033P019N018: std_logic_vector(   0 downto 0);
        signal cVar1S18S118P035N033P019N018: std_logic_vector(   0 downto 0);
        signal cVar1S19S118P035N033P019N018: std_logic_vector(   0 downto 0);
        signal cVar1S20S118P035N033P019N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S118P035P046P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S22S118P035P046P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S23S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S24S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S25S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S26S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S27S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S28S118P035N046P022P034: std_logic_vector(   0 downto 0);
        signal cVar1S29S118P035N046P022P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S118P035N046P022N065: std_logic_vector(   0 downto 0);
        signal cVar1S31S118P035N046P022N065: std_logic_vector(   0 downto 0);
        signal cVar1S0S119P065P027P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S119P065P027P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S119P065P027P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S119P065P027P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S119P065P027P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S5S119P065P027P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S6S119P065N027P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S7S119P065N027P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S8S119P065N027P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S119P065N027P037N016: std_logic_vector(   0 downto 0);
        signal cVar1S10S119P065N027P037N016: std_logic_vector(   0 downto 0);
        signal cVar1S11S119P065N027P037N016: std_logic_vector(   0 downto 0);
        signal cVar1S12S119P065N027P037P008: std_logic_vector(   0 downto 0);
        signal cVar1S13S119P065N027P037P008: std_logic_vector(   0 downto 0);
        signal cVar1S14S119P065N027P037P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S119P065N027P037P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S119P065N027P037N008: std_logic_vector(   0 downto 0);
        signal cVar1S17S119P065N027P037N008: std_logic_vector(   0 downto 0);
        signal cVar1S18S119P065P008P064P069: std_logic_vector(   0 downto 0);
        signal cVar1S19S119P065P008P064P069: std_logic_vector(   0 downto 0);
        signal cVar1S20S119P065P008P064P069: std_logic_vector(   0 downto 0);
        signal cVar1S21S119P065P008P064P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S119P065P008P064P069: std_logic_vector(   0 downto 0);
        signal cVar1S23S119P065P008P064P014: std_logic_vector(   0 downto 0);
        signal cVar1S24S119P065P008P064P014: std_logic_vector(   0 downto 0);
        signal cVar1S25S119P065P008P064P014: std_logic_vector(   0 downto 0);
        signal cVar1S26S119P065P008P064N014: std_logic_vector(   0 downto 0);
        signal cVar1S27S119P065P008P064N014: std_logic_vector(   0 downto 0);
        signal cVar1S28S119P065P008P064N014: std_logic_vector(   0 downto 0);
        signal cVar1S29S119P065P008P064N014: std_logic_vector(   0 downto 0);
        signal cVar1S30S119P065P008P011P014: std_logic_vector(   0 downto 0);
        signal cVar1S31S119P065P008P011P014: std_logic_vector(   0 downto 0);
        signal cVar1S32S119P065P008P011P014: std_logic_vector(   0 downto 0);
        signal cVar1S33S119P065P008N011P056nsss: std_logic_vector(   0 downto 0);
        signal cVar1S34S119P065P008N011N056: std_logic_vector(   0 downto 0);
        signal cVar1S35S119P065P008N011N056: std_logic_vector(   0 downto 0);
        signal cVar1S0S120P037P001P032P018: std_logic_vector(   0 downto 0);
        signal cVar1S1S120P037P001P032P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S120P037P001P032P018: std_logic_vector(   0 downto 0);
        signal cVar1S3S120P037P001P032P018: std_logic_vector(   0 downto 0);
        signal cVar1S4S120P037P001P032N018: std_logic_vector(   0 downto 0);
        signal cVar1S5S120P037P001P032N018: std_logic_vector(   0 downto 0);
        signal cVar1S6S120P037P001N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S120P037P001N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S120P037P001N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S120P037P001N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S120P037P001N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S11S120P037P001N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S12S120P037P001N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S13S120P037P001P036P019: std_logic_vector(   0 downto 0);
        signal cVar1S14S120P037P001P036P019: std_logic_vector(   0 downto 0);
        signal cVar1S15S120P037P001P036P019: std_logic_vector(   0 downto 0);
        signal cVar1S16S120P037P001P036N019: std_logic_vector(   0 downto 0);
        signal cVar1S17S120P037P001P036P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S120N037P036P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S120N037P036P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S20S120N037P036P065P017: std_logic_vector(   0 downto 0);
        signal cVar1S21S120N037P036P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S22S120N037P036P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S23S120N037P036P065N017: std_logic_vector(   0 downto 0);
        signal cVar1S24S120N037P036P065P016: std_logic_vector(   0 downto 0);
        signal cVar1S25S120N037P036P065P016: std_logic_vector(   0 downto 0);
        signal cVar1S26S120N037P036P065P016: std_logic_vector(   0 downto 0);
        signal cVar1S27S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S28S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S29S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S30S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S31S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S32S120N037N036P034P050: std_logic_vector(   0 downto 0);
        signal cVar1S33S120N037N036N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S34S120N037N036N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S35S120N037N036N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S36S120N037N036N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S37S120N037N036N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S0S121P065P052P034P009: std_logic_vector(   0 downto 0);
        signal cVar1S1S121P065P052P034P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S121P065P052P034P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S121P065P052P034N009: std_logic_vector(   0 downto 0);
        signal cVar1S4S121P065P052P034N009: std_logic_vector(   0 downto 0);
        signal cVar1S5S121P065P052P034P011: std_logic_vector(   0 downto 0);
        signal cVar1S6S121P065P052P034N011: std_logic_vector(   0 downto 0);
        signal cVar1S7S121P065N052P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S8S121P065N052P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S9S121P065N052P050P046: std_logic_vector(   0 downto 0);
        signal cVar1S10S121P065N052P050N046: std_logic_vector(   0 downto 0);
        signal cVar1S11S121P065N052P050N046: std_logic_vector(   0 downto 0);
        signal cVar1S12S121P065N052P050N046: std_logic_vector(   0 downto 0);
        signal cVar1S13S121P065N052P050P060: std_logic_vector(   0 downto 0);
        signal cVar1S14S121P065N052P050P060: std_logic_vector(   0 downto 0);
        signal cVar1S15S121P065N052P050P060: std_logic_vector(   0 downto 0);
        signal cVar1S16S121P065N052P050N060: std_logic_vector(   0 downto 0);
        signal cVar1S17S121P065N052P050N060: std_logic_vector(   0 downto 0);
        signal cVar1S18S121P065N052P050N060: std_logic_vector(   0 downto 0);
        signal cVar1S19S121P065P036P024P030: std_logic_vector(   0 downto 0);
        signal cVar1S20S121P065P036P024N030: std_logic_vector(   0 downto 0);
        signal cVar1S21S121P065P036P024N030: std_logic_vector(   0 downto 0);
        signal cVar1S22S121P065P036P024N030: std_logic_vector(   0 downto 0);
        signal cVar1S23S121P065P036P024N030: std_logic_vector(   0 downto 0);
        signal cVar1S24S121P065P036P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S25S121P065N036P008P041: std_logic_vector(   0 downto 0);
        signal cVar1S26S121P065N036P008P041: std_logic_vector(   0 downto 0);
        signal cVar1S27S121P065N036P008P041: std_logic_vector(   0 downto 0);
        signal cVar1S28S121P065N036P008P041: std_logic_vector(   0 downto 0);
        signal cVar1S29S121P065N036P008P037: std_logic_vector(   0 downto 0);
        signal cVar1S30S121P065N036P008P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S121P065N036P008N037: std_logic_vector(   0 downto 0);
        signal cVar1S32S121P065N036P008N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S122P052P009P056nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S122P052P009N056P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S122P052P009N056N010: std_logic_vector(   0 downto 0);
        signal cVar1S3S122P052P009N056N010: std_logic_vector(   0 downto 0);
        signal cVar1S4S122P052N009P056P046: std_logic_vector(   0 downto 0);
        signal cVar1S5S122P052N009P056P046: std_logic_vector(   0 downto 0);
        signal cVar1S6S122P052N009P056P046: std_logic_vector(   0 downto 0);
        signal cVar1S7S122P052N009P056P046: std_logic_vector(   0 downto 0);
        signal cVar1S8S122P052N009P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S122P052N009P056N015: std_logic_vector(   0 downto 0);
        signal cVar1S10S122N052P046P050P042: std_logic_vector(   0 downto 0);
        signal cVar1S11S122N052P046P050P042: std_logic_vector(   0 downto 0);
        signal cVar1S12S122N052P046P050P042: std_logic_vector(   0 downto 0);
        signal cVar1S13S122N052P046P050P042: std_logic_vector(   0 downto 0);
        signal cVar1S14S122N052P046P050P042: std_logic_vector(   0 downto 0);
        signal cVar1S15S122N052P046P050P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S122N052N046P065P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S122N052N046P065P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S122N052N046P065P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S122N052N046P065P008: std_logic_vector(   0 downto 0);
        signal cVar1S20S122N052N046P065P008: std_logic_vector(   0 downto 0);
        signal cVar1S21S122N052N046N065P049: std_logic_vector(   0 downto 0);
        signal cVar1S22S122N052N046N065P049: std_logic_vector(   0 downto 0);
        signal cVar1S23S122N052N046N065N049: std_logic_vector(   0 downto 0);
        signal cVar1S0S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S1S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S2S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S3S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S4S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S5S123P017P036P016P021: std_logic_vector(   0 downto 0);
        signal cVar1S6S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S7S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S8S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S9S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S10S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S123P017P036N016P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S123P017P036P056P052: std_logic_vector(   0 downto 0);
        signal cVar1S13S123P017P036P056P052: std_logic_vector(   0 downto 0);
        signal cVar1S14S123P017P036P056P052: std_logic_vector(   0 downto 0);
        signal cVar1S15S123P017P036N056P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S123P017P036N056P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S123P017P036N056N065: std_logic_vector(   0 downto 0);
        signal cVar1S18S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S19S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S20S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S21S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S24S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S25S123P017P036P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S123P017P036P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S27S123P017P036P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S28S123P017P036P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S29S123P017P036P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S30S123P017P036P065N063: std_logic_vector(   0 downto 0);
        signal cVar1S31S123P017N036P060P069: std_logic_vector(   0 downto 0);
        signal cVar1S32S123P017N036P060P069: std_logic_vector(   0 downto 0);
        signal cVar1S33S123P017N036P060P069: std_logic_vector(   0 downto 0);
        signal cVar1S34S123P017N036P060N069: std_logic_vector(   0 downto 0);
        signal cVar1S35S123P017N036P060N069: std_logic_vector(   0 downto 0);
        signal cVar1S36S123P017N036P060N069: std_logic_vector(   0 downto 0);
        signal cVar1S37S123P017N036N060P037: std_logic_vector(   0 downto 0);
        signal cVar1S38S123P017N036N060P037: std_logic_vector(   0 downto 0);
        signal cVar1S39S123P017N036N060P037: std_logic_vector(   0 downto 0);
        signal cVar1S40S123P017N036N060P037: std_logic_vector(   0 downto 0);
        signal cVar1S41S123P017N036N060N037: std_logic_vector(   0 downto 0);
        signal cVar1S42S123P017N036N060N037: std_logic_vector(   0 downto 0);
        signal cVar1S43S123P017N036N060N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S124P036P065P032P019: std_logic_vector(   0 downto 0);
        signal cVar1S1S124P036P065P032P019: std_logic_vector(   0 downto 0);
        signal cVar1S2S124P036P065P032P019: std_logic_vector(   0 downto 0);
        signal cVar1S3S124P036P065P032P019: std_logic_vector(   0 downto 0);
        signal cVar1S4S124P036P065P032P019: std_logic_vector(   0 downto 0);
        signal cVar1S5S124P036P065P032P055: std_logic_vector(   0 downto 0);
        signal cVar1S6S124P036P065P032P055: std_logic_vector(   0 downto 0);
        signal cVar1S7S124P036P065P024P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S124P036P065P024P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S124P036P065P024P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S124P036P065P024P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S124P036P065P024N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S124P036P065P024N063: std_logic_vector(   0 downto 0);
        signal cVar1S13S124P036P065P024N063: std_logic_vector(   0 downto 0);
        signal cVar1S14S124P036P065P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S15S124N036P017P034P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S124N036P017P034N043: std_logic_vector(   0 downto 0);
        signal cVar1S17S124N036P017P034N043: std_logic_vector(   0 downto 0);
        signal cVar1S18S124N036P017P034N043: std_logic_vector(   0 downto 0);
        signal cVar1S19S124N036P017P034N043: std_logic_vector(   0 downto 0);
        signal cVar1S20S124N036P017N034P002: std_logic_vector(   0 downto 0);
        signal cVar1S21S124N036P017N034P002: std_logic_vector(   0 downto 0);
        signal cVar1S22S124N036P017N034P002: std_logic_vector(   0 downto 0);
        signal cVar1S23S124N036P017N034P002: std_logic_vector(   0 downto 0);
        signal cVar1S24S124N036N017P032P031: std_logic_vector(   0 downto 0);
        signal cVar1S25S124N036N017P032P031: std_logic_vector(   0 downto 0);
        signal cVar1S26S124N036N017P032P031: std_logic_vector(   0 downto 0);
        signal cVar1S27S124N036N017P032P031: std_logic_vector(   0 downto 0);
        signal cVar1S28S124N036N017N032P046: std_logic_vector(   0 downto 0);
        signal cVar1S29S124N036N017N032P046: std_logic_vector(   0 downto 0);
        signal cVar1S30S124N036N017N032N046: std_logic_vector(   0 downto 0);
        signal cVar1S31S124N036N017N032N046: std_logic_vector(   0 downto 0);
        signal cVar1S0S125P032P064P050P022: std_logic_vector(   0 downto 0);
        signal cVar1S1S125P032P064P050P022: std_logic_vector(   0 downto 0);
        signal cVar1S2S125P032P064P050P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S125P032P064P050P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S125P032P064P050P022: std_logic_vector(   0 downto 0);
        signal cVar1S5S125P032P064P050P027: std_logic_vector(   0 downto 0);
        signal cVar1S6S125P032P064P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S7S125P032P064P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S8S125P032P064P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S125P032N064P037P068: std_logic_vector(   0 downto 0);
        signal cVar1S10S125P032N064P037P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S125P032N064P037P068: std_logic_vector(   0 downto 0);
        signal cVar1S12S125P032N064P037N068: std_logic_vector(   0 downto 0);
        signal cVar1S13S125P032N064P037N068: std_logic_vector(   0 downto 0);
        signal cVar1S14S125P032N064P037N068: std_logic_vector(   0 downto 0);
        signal cVar1S15S125P032N064P037P056: std_logic_vector(   0 downto 0);
        signal cVar1S16S125P032N064P037P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S125P032N064P037P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S125P032N064P037P056: std_logic_vector(   0 downto 0);
        signal cVar1S19S125P032N064P037N056: std_logic_vector(   0 downto 0);
        signal cVar1S20S125P032N064P037N056: std_logic_vector(   0 downto 0);
        signal cVar1S21S125P032N064P037N056: std_logic_vector(   0 downto 0);
        signal cVar1S22S125P032P037P063P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S125P032P037P063P016: std_logic_vector(   0 downto 0);
        signal cVar1S24S125P032P037P063P016: std_logic_vector(   0 downto 0);
        signal cVar1S25S125P032P037N063P012: std_logic_vector(   0 downto 0);
        signal cVar1S26S125P032P037N063P012: std_logic_vector(   0 downto 0);
        signal cVar1S27S125P032P037N063N012: std_logic_vector(   0 downto 0);
        signal cVar1S28S125P032P037N063N012: std_logic_vector(   0 downto 0);
        signal cVar1S29S125P032N037P031P068: std_logic_vector(   0 downto 0);
        signal cVar1S30S125P032N037P031P068: std_logic_vector(   0 downto 0);
        signal cVar1S31S125P032N037P031P068: std_logic_vector(   0 downto 0);
        signal cVar1S32S125P032N037P031N068: std_logic_vector(   0 downto 0);
        signal cVar1S33S125P032N037P031N068: std_logic_vector(   0 downto 0);
        signal cVar1S34S125P032N037P031P012: std_logic_vector(   0 downto 0);
        signal cVar1S35S125P032N037P031P012: std_logic_vector(   0 downto 0);
        signal cVar1S36S125P032N037P031P012: std_logic_vector(   0 downto 0);
        signal cVar1S0S126P069P018P026P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S126P069P018P026N064: std_logic_vector(   0 downto 0);
        signal cVar1S2S126P069P018P026N064: std_logic_vector(   0 downto 0);
        signal cVar1S3S126P069P018N026P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S126P069P018N026N031: std_logic_vector(   0 downto 0);
        signal cVar1S5S126P069P018N026N031: std_logic_vector(   0 downto 0);
        signal cVar1S6S126P069P018N026N031: std_logic_vector(   0 downto 0);
        signal cVar1S7S126P069P018N026N031: std_logic_vector(   0 downto 0);
        signal cVar1S8S126P069P018P068P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S126P069P018P068P067: std_logic_vector(   0 downto 0);
        signal cVar1S10S126P069P018P068P067: std_logic_vector(   0 downto 0);
        signal cVar1S11S126P069P018P068N067: std_logic_vector(   0 downto 0);
        signal cVar1S12S126P069P018P068N067: std_logic_vector(   0 downto 0);
        signal cVar1S13S126P069P018P068P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S126P069P018P068N040: std_logic_vector(   0 downto 0);
        signal cVar1S15S126P069P018P068N040: std_logic_vector(   0 downto 0);
        signal cVar1S16S126P069P018P068N040: std_logic_vector(   0 downto 0);
        signal cVar1S17S126N069P018P049P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S126N069P018P049P032: std_logic_vector(   0 downto 0);
        signal cVar1S19S126N069P018P049P032: std_logic_vector(   0 downto 0);
        signal cVar1S20S126N069P018N049P032: std_logic_vector(   0 downto 0);
        signal cVar1S21S126N069P018N049N032: std_logic_vector(   0 downto 0);
        signal cVar1S22S126N069P018N049N032: std_logic_vector(   0 downto 0);
        signal cVar1S23S126N069P018N049N032: std_logic_vector(   0 downto 0);
        signal cVar1S24S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S25S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S26S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S27S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S28S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S29S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S30S126N069N018P066P064: std_logic_vector(   0 downto 0);
        signal cVar1S31S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S32S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S33S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S34S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S35S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S36S126N069N018P066P006: std_logic_vector(   0 downto 0);
        signal cVar1S0S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S1S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S2S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S3S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S4S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S5S127P064P069P034P016: std_logic_vector(   0 downto 0);
        signal cVar1S6S127P064P069P034P008: std_logic_vector(   0 downto 0);
        signal cVar1S7S127P064P069P034P008: std_logic_vector(   0 downto 0);
        signal cVar1S8S127P064P069P034P008: std_logic_vector(   0 downto 0);
        signal cVar1S9S127P064P069P034P008: std_logic_vector(   0 downto 0);
        signal cVar1S10S127P064P069P034P008: std_logic_vector(   0 downto 0);
        signal cVar1S11S127P064P069P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S12S127P064P069P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S13S127P064P069P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S14S127P064P069P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S15S127P064P069N037P016: std_logic_vector(   0 downto 0);
        signal cVar1S16S127P064P069N037P016: std_logic_vector(   0 downto 0);
        signal cVar1S17S127P064P069N037P016: std_logic_vector(   0 downto 0);
        signal cVar1S18S127P064P069N037P016: std_logic_vector(   0 downto 0);
        signal cVar1S19S127P064P069N037N016: std_logic_vector(   0 downto 0);
        signal cVar1S20S127P064P069N037N016: std_logic_vector(   0 downto 0);
        signal cVar1S21S127P064P069N037N016: std_logic_vector(   0 downto 0);
        signal cVar1S22S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S23S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S24S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S25S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S26S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S27S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S28S127P064P018P054P035: std_logic_vector(   0 downto 0);
        signal cVar1S29S127P064P018P054P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S127P064P018P054N065: std_logic_vector(   0 downto 0);
        signal cVar1S31S127P064P018P054N065: std_logic_vector(   0 downto 0);
        signal cVar1S32S127P064N018P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S33S127P064N018P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S34S127P064N018P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S35S127P064N018P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S36S127P064N018P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S37S127P064N018P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S38S127P064N018P050N027: std_logic_vector(   0 downto 0);
        signal cVar2S0S0P062P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S0P062P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S0N062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S0P058P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S0P058N033P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S0N058P068P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S0N058N068P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S0P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S0N036P065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S0P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S0N062P068P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S0N062N068P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S0P018P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S0P018N062P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S0N018P016P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S0P068P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S0N068P067P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S0P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S0P068P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S0P068N066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S0N068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S0N068N064P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S0P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S0P064N016P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S0N064P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S0N064N068P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S0P034P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S0P034N062P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S0P015P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S0P015N032P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S0N015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S0N015N066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S0P013P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S0P013N030P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S0N013P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S0N013N068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S0P051P028P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S0N051P047P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S1P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S1P062P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S1P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S1N029P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S1P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S1P066P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S1P008P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S1N008psss: std_logic_vector(   0 downto 0);
        signal cVar2S9S1P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S1P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S1P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S1P062P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S1P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S1P030P012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S1P030N012P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S1N030P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S1N030N028P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S1P033P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S1P033P069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S1N033P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S1N033N035P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S1P035P058P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S1P035N058P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S1N035P014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S1P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S1N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S1N006N008P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S1P064P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S1P064N051P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S1N064N068P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S2P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S2P043N022P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S2N043P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S2N043P047P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S2P064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S2P064N015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S2P064P059P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S2P064P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S2P064N019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S2P028P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S2N028P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S2P018P019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S2P018P019psss: std_logic_vector(   0 downto 0);
        signal cVar2S13S2P018P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S2P018P069P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S2P018P069psss: std_logic_vector(   0 downto 0);
        signal cVar2S16S2N018P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S2P006P014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S2P060P069P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S2P060P069psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S2P060P058P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S2P064P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S2N064P060P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S2P066P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S2P064P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S2P064N014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S2P064P017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S2P064P017P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S2P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S2N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S2N026N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S2P050P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S2P050N052P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S2N050P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S2N050N046P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S2P064P037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S2P064N037P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S2N064P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S2N064N059P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S3P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S3N024P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S3P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S3N024P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S3N024N023P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S3P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S3P065P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S3P065N016P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S3P014P017P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S3P062P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S3P062P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S3P018P069P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S3P018P069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S3P018P069P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S3P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S3P065P069P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S3N065P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S3N065N061P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S3P065P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S3P065P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S3P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S3N009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S3N009N011P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S3P039P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S3P039N041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S3N039P047P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S4P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S4P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S4N017P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S4P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S4P011P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S4P011N024P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S4P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S4P034P014P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S4P034P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S4P016P010P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S4N016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S4P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S4P011P033P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S4P011P007P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S4P012P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S4P012P030P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S4N012P064P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S4N012N064psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S4P014P035P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S4P069P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S4P069N063P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S4P069P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S4P069N029P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S4P033P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S4N033P035P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S4N033N035P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S5P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S5N008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S5N008N019P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S5P053P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S5P053P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S5P053P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S5P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S5P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S5N038P012P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S5N038N012P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S5P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S5P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S5P036N066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S5N036P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S5N036N018P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S5P056P019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S5P056P019P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S5N056P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S5N056N019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S5P016P013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S5P016P030P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S5P016N030P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S5P065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S5P065N018P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S5P065P011P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S5P029P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S5P029N010P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S5N029P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S5N029N064P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S6P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S6P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S6N018P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S6P033P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S6N033P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S6P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S6P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S6P058P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S6N058P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S6N058N045P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S6P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S6P019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S6P019P069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S6P012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S6P012N011P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S6N012P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S6N012N028P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S6P066P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S6P066N058P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S6P066P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S6P061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S6P061N059P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S6N061P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S6N061N050P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S7P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S7P010N052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S7N010P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S7N010N025P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S7P025P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S7P025N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S7N025P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S7N025N006P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S7P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S7N021P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S7N021N023P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S7P069P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S7N069P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S7N069N031P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S7P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S7N041P020P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S7P051P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S7P051N008P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S7P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S7P064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S7P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S7N017P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S7P017P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S7P017P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S7P016N017P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S7P016P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S8P044P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S8P044P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S8P044N005P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S8P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S8P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S8P068P066P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S8N068P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S8P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S8N004P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S8N004N017P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S8P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S8N049P051P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S8N049N051P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S8P057P049P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S8N057P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S8N057N025P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S8P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S8N016P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S8P001P010P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S8P044P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S8N044P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S9P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S9P066P069P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S9P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S9P066N018P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S9P058P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S9P058P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S9N058P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S9N058N057P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S9P006P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S9P006N065P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S9P068P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S9P059P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S9N059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S9P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S9P064P017P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S9N064P061P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S9N064P061P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S9P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S9N022P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S9P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S9N068P041P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S9N068N041P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S9P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S9N025P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S9N025N022P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S9P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S9N021P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S9N021N023P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S9P003P033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S9P003N033psss: std_logic_vector(   0 downto 0);
        signal cVar2S34S9P003P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S9P003N039P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S10P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S10P066P069P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S10P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S10P066N069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S10P033P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S10P033N047P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S10P006P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S10P006N065P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S10P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S10N059P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S10N059N016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S10P059P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S10N059P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S10P061P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S10P061P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S10P061N068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S10P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S10P036N017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S10N036P044P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S10N036P044P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S10P036P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S10P036N042P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S10P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S10N045P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S10P022P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S10P022N007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S10N022P024P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S10N022N024P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S10P058P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S10P058N014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S10N058P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S10P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S10P044N023P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S10N044P047P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S10N044N047P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S11P069P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S11P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S11P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S11N010P048P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S11P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S11N049P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S11P024P001P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S11P041P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S11P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S11N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S11N022N023P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S11P066P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S11P035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S11P035P066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S11P068P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S11N068P054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S11N068N054P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S11P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S11N038P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S11P013P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S11P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S12P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S12P062P018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S12P062N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S12P063P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S12N063P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S12N063N055P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S12P014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S12P014P034P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S12P014P056P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S12P014N056P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S12P034P017P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S12P034N017psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S12N034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S12N034N037P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S12P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S12P013P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S12P013P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S12P013N059P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S12P064P033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S12P064P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S12P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S12N055P069P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S12P036P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S12N036P053P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S12P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S12N054P012P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S12N054P012P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S12P064P003P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S12P064P032P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S12P064N032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S12P055P012P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S12P055P012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S12P064P034P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S12P005P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S12P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S12P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S12P010P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S12P010P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S12P065P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S13P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S13P012P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S13P031P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S13P031P028P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S13P031P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S13P048P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S13N048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S13N048N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S13P030P012P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S13P030N012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S13N030psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S13P001P065P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S13P001P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S13P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S13N055P019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S13N055N019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S13P049P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S13P049P003P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S13P009P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S13P009P026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S13P009N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S13P069P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S13P069N062P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S13P069P058P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S13P032P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S13N032P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S13P065P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S13P065N015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S13N065P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S13P065P037P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S13P065N037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S13P065P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S13P065N014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S13P030P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S13P030N015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S13N030P055P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S14P011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S14P011P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S14N011P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S14N011P064P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S14P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S14N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S14N018N037P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S14P008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S14P008P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S14P069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S14P013P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S14N013P034P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S14P029N062P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S14P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S14P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S14P062P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S14P062N052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S14P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S14P050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S14P050N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S14P052P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S14P052N008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S14P000P034P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S14P000P034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S14P025P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S14N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S14N025N027P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S14P012P052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S14P012P052P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S14P012P031P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S14P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S14P040N021P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S14N040P032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S15P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S15N021P035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S15N021N035P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S15P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S15P046P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S15P008P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S15N008P049P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S15P009P013P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S15P009P013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S15N009P068P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S15P008P067P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S15P008N067P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S15P008P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S15P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S15N069P019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S15N069N019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S15P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S15N018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S15P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S15P047N026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S15N047P058P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S15P047P031P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S15P047N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S15P047P007P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S15P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S15N018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S15P028P018P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S15N028P069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S16P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S16P068P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S16P069P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S16P069N005P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S16P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S16P068P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S16P068psss: std_logic_vector(   0 downto 0);
        signal cVar2S9S16P049P044P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S16P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S16P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S16P011P013P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S16N011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S16N011N018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S16P014P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S16P014N061P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S16P014P058P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S16P014N058P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S16P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S16P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S16N005P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S16P013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S16P013N022P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S16P033P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S16P033P054P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S16P033P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S16P033N069P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S16P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S16P044N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S16N044P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S16N044N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S17P059P063P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S17P059N063psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S17N059P058P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S17P033P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S17P033N018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S17P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S17P036N018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S17N036P013P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S17P036P012P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S17P017P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S17P017P054P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S17P017P018P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S17P017P018P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S17P017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S17P017P068P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S17N017P026P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S17N017N026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S17P014P064P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S17P014P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S17P014N064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S17P010P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S17P010N033P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S17N010P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S17N010N039P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S17P068P067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S17P068N067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S17N068P014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S17N068N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S17P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S17P017P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S17P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S17P005P053P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S18P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S18P012P014P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S18N012P064P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S18N012N064P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S18P053P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S18P053P050P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S18N053P036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S18N053N036psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S18P036P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S18N036P019P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S18P064P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S18N064P032P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S18P068P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S18P068P036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S18N068P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S18N068N045P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S18P033P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S18N033P002P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S18P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S18N069P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S18P018P055P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S18P018P055P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S18N018P017P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S18P018P055P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S18P018P066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S18P018P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S18P066P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S18P066P010P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S18N066P059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S18P014P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S18P014P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S18P015P016P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S18P015N016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S18P017P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S19P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S19P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S19P056P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S19P056P062P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S19N056P055P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S19P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S19N056P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S19P069P062P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S19P069N062psss: std_logic_vector(   0 downto 0);
        signal cVar2S9S19P069P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S19P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S19P037N018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S19P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S19N014P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S19P011P069P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S19N011P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S19P010P054P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S19P010P054P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S19P010P014P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S19P010P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S19P035P009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S19P035P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S19P059P010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S19P035P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S19N035P016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S19P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S19N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S19N022N024P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S19P008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S19P008N009P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S19N008P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S19P051P026P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S19P051N026P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S19N051P028P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S19P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S19P039N020P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S19N039P030P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S20P006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S20P006P019P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S20P006P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S20P005P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S20P005P015P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S20P003P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S20P003P068psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S20P003P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S20P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S20N014P019P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S20N014N019P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S20P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S20P066P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S20P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S20N007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S20N007N009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S20P010P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S20P010N046P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S20P010P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S20P015P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S20P015P059P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S20P015P061P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S20P015N061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S20P015P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S20P015N061P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S20N015P016P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S20N015N016P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S20P050P042P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S20P050N042P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S20P050P008P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S20P064P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S20P064P067P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S20P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S20N030P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S20P050P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S21P035P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S21P035P046P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S21P035psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S21P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S21P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S21N016P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S21P046P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S21N046P061P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S21N046N061P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S21P037P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S21P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S21P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S21P011P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S21N011P055P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S21N011P055psss: std_logic_vector(   0 downto 0);
        signal cVar2S17S21P014P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S21P014N040P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S21P014P012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S21P014N012P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S21P034P012P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S21P034N012P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S21P034P007P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S21P067P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S21P067N056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S21P067P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S21P017P014P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S21P017N014psss: std_logic_vector(   0 downto 0);
        signal cVar2S29S21N017P015P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S21N017N015P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S21P028P062P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S21P028P062P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S21N028P029P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S22P045P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S22P045P019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S22P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S22N043P046P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S22N043N046P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S22P037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S22P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S22N007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S22N007N005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S22P036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S22N036psss: std_logic_vector(   0 downto 0);
        signal cVar2S13S22P066P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S22P066P037P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S22P031P012P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S22P031N012P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S22N031P069P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S22N031N069P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S22P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S22P036P037P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S22N036P019P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S22N036P019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S22P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S22N003P033P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S22P017P046P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S22P017P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S22P017P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S22P062P018P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S22P062N018P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S22P062P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S23P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S23P016N018P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S23P002P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S23P002N061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S23P002P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S23P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S23P020P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S23P020N040psss: std_logic_vector(   0 downto 0);
        signal cVar2S10S23P020P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S23P044P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S23P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S23N026P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S23N026N014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S23P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S23N004P003P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S23P009P047P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S23P009P047P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S23P027P000P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S23N027P017P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S23N027N017P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S24P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S24P046P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S24P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S24P016N018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S24P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S24N045P037P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S24N045N037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S24P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S24P059N015P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S24N059P006P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S24P018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S24P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S24N062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S24N062N012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S24P023P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S24P023N018P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S24N023P002P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S24P020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S24P020N005P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S24N020P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S24P021P026P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S24P021P019P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S24P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S24P048P013P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S24N048N069P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S25P017P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S25P017N056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S25N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S25N017N018P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S25P018P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S25P062P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S25N062P005P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S25P054P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S25P054N014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S25P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S25N055P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S25P059P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S25P059N013P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S25N059P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S25N059P013P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S25P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S25P015N068P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S25N015P049P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S25N015N049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S25P028P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S25P028P051P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S25N028P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S25N028N032P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S25P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S25P016P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S25P016N019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S25P029P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S25N029P037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S25N029N037P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S26P028P051P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S26P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S26N069P063P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S26P047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S26P065P035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S26P065N035P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S26N065P067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S26N065N067P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S26P002P065P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S26P002N065P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S26P002P012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S26P034P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S26P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S26N037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S26P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S26N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S26N024N025P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S26P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S26P016P014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S26P018P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S26P018N069P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S26N018P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S26P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S26N057P056P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S26N057N056P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S26P064P054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S26P064P054P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S26N064P010P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S26N064N010P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S26P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S26N013P014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S26N013N014P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S26P063P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S26P063N055P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S26N063P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S26P047P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S26N047P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S26N047N046P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S26P023P042P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S26P023N042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S26N023P053P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S27P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S27N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S27N003N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S27P018P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S27P018N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S27P003P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S27P003N039P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S27P017P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S27N017P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S27N017N008P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S27P010P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S27P035P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S27P035P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S27P035P016P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S27P059P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S27P059P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S27P059P061P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S27P059N061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S27P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S27P053P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S27N053P069P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S28P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S28P036P069P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S28P059P058P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S28P059P058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S28N059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S28P034P010P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S28P034N010psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S28P034P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S28P034N064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S28P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S28P003P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S28P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S28P010P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S28P010N066P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S28P002P007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S28P002N007psss: std_logic_vector(   0 downto 0);
        signal cVar2S17S28P002P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S28P035P068P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S28P031P057P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S28P031P019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S28P031N019P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S28P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S28P039N020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S28N039P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S29P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S29N004P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S29N004N019P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S29P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S29N062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S29N062N012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S29P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S29N036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S29P046P035P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S29P063P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S29P063P062P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S29N063P064P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S29N063N064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S29P050P016P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S29P050P016P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S29P050P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S29P051P012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S29P014P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S29P015P036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S30P009P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S30N009P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S30N009P062P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S30P006P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S30P006N026P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S30P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S30P009P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S30N009P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S30P029P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S30P029P051P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S30N029P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S30N029N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S30P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S30P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S30P035N017P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S30P035P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S30P053P049P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S30N053P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S30N053N057P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S30P065P067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S30P065P067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S30P065P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S30P065N036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S30P024P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S30P024P049P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S30N024P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S30P064P028P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S30P064P028P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S30P037P029P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S30N037P061P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S30N037N061P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S30P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S30P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S30N069P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S30P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S30P010P019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S30N010P017P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S30N010N017P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S31P019P017P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S31P019N017P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S31P019P059P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S31P019P059P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S31P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S31P066N019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S31P067P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S31P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S31P017P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S31P017P015P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S31P017N015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S31P062P035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S31P062N035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S31N062P055P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S31N062N055P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S31P034P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S31P034P015P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S31P034P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S31P034N068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S31P067P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S31N067P058P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S31P051P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S31P051P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S31P051P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S31P051N019P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S31P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S31P056P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S31P056N069P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S31P067P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S31P067N049P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S31N067P066P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S31N067N066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S31P037P005P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S31N037P059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S31N037N059P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S31P015P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S31P015N047P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S31P015P016P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S31P015P016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S31P016P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S31P016N068P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S31N016P048P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S43S31N016N048P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S32P023P019P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S32P023P019P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S32P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S32P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S32P034P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S32P034P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S32P034N059P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S32P003P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S32N003P008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S32P017P062P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S32P017P062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S32N017P018P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S32P019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S32P033P064P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S32P033P064P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S32N033P054P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S32P035P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S32P035N032P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S32N035P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S32N035N017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S32P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S32P019P067P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S32P019N067psss: std_logic_vector(   0 downto 0);
        signal cVar2S24S32P019P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S32P019P067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S32P056P038P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S32P056N038P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S32P056P069P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S32P014P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S32N014P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S32N014N015P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S32P018P061P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S33P053P008P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S33P053P008P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S33P035P045P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S33P035P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S33P027P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S33N027P025P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S33N027N025P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S33P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S33P066P062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S33P010P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S33P010N015P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S33N010P053P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S33N010N053P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S33P010P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S33P010N016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S33P010P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S33P023P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S33P023N044P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S33N023P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S33N023N050P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S33P019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S33P019P013P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S33N019P007P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S33P035P062P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S33P035N062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S33P035P016P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S33P018P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S33P015P003P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S33N015P019P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S33P016P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S34P041P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S34N041P063P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S34N041N063psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S34P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S34N010P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S34P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S34P061P013P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S34P013P035P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S34P013P035P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S34N013P015P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S34N013N015P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S34P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S34N066P015P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S34N066P015P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S34P017P058P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S34P017P058P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S34N017P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S34P016P060P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S34N016P012P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S34N016P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S34P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S34P066N069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S34P066P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S34P066N011P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S34P035P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S34P035P012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S34P035P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S34P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S34N014P069P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S34P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S34N059P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S34N059N037P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S34P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S34P036N015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S34N036P019P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S34N036N019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S34P066P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S34P066P060P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S34P066P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S34P061P068P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S34P061N068P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S34N061P060P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S34P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S43S34P050P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S44S34N050P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S35P016P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S35P016N057P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S35P033P058P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S35P033P058P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S35N033P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S35N033P056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S35P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S35P018P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S35P018P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S35N018P068P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S35P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S35P056P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S35P056P052P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S35P056P054P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S35P064P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S35P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S35P033P055P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S35P033P055P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S35P033P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S35P033N017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S35P018P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S35P018N015P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S35P035P036P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S35P035P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S35P049P009P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S35N049N067P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S36P035P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S36P035P019P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S36N035P025P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S36N035P025P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S36P052P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S36P017P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S36P017N061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S36N017P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S36P034P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S36P012P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S36P012N060P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S36N012P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S36N012N040P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S36P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S36P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S36P058P066P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S36P058P066P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S36P058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S36P058P018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S36P062P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S36P062N018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S36P062P060P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S36P035P034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S36P035P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S36P014P010P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S36N014P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S36P052P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S36P052N026P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S36P052P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S36P026P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S36P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S36N043P035P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S36P068P066P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S36N068P069P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S37P066P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S37P066N036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S37N066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S37P011P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S37N011P062P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S37N011N062P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S37P044P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S37P052P060P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S37P014P034P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S37P014P034P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S37P014P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S37P014N047P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S37P058P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S37P058N014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S37P058P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S37P019P010P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S37P019P010P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S37P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S37P012P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S37P012P033P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S37N012P014P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S37N012N014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S37P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S37P066P069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S37P066P036P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S37P066N036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S37P018P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S37P018N057P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S37N018P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S37P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S37P017N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S37N017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S37N017N068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S37P058P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S38P024P029P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S38P024P029P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S38P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S38N062P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S38P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S38N064P003P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S38P062P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S38P062P058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S38P062P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S38P062P067P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S38P011P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S38P011P010P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S38P011P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S38P011N027P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S38P007P011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S38P061P015P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S38P061P015P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S38P061P017P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S38P015P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S38P015N061P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S38N015P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S38P056P057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S38P056P057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S38N056P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S38N056N018P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S38P066P007P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S38P020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S38P020N005P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S38N020P013P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S38P011P060P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S38P011N060psss: std_logic_vector(   0 downto 0);
        signal cVar2S31S38N011P024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S38P064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S38P064P015P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S38P064P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S38P054P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S38P054P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S38P065P063P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S38N065P035P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S39P019P059P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S39P019N059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S39P019P068P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S39P019N068P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S39P068P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S39P068P065P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S39N068P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S39N068N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S39P056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S39P056P057P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S39N056P054P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S39P015P035P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S39P015N035P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S39P037P018P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S39P037N018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S39P037P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S39P037P036P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S39P046P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S39N046P015P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S39P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S39P067P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S39N067P019P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S39P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S39N057P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S39N057N036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S39P009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S39P009N069P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S39P009P018P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S39P037P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S39P037N069P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S39N037P061P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S39P014P015P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S39P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S39N034P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S39N034N018P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S39P026P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S39P026N057P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S39P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S39N026P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S39P067P054P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S39P067P055P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S40P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S40P058P012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S40P058N012P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S40P019P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S40N019P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S40P068P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S40P068N063P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S40P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S40P068P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S40P068N017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S40N068P060P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S40N068N060P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S40P057P006P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S40P030P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S40P030P059P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S40P030P011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S40P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S40N011P056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S40N011P056P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S40P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S40P033P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S40P054P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S40N054P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S40N054N011P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S40P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S40N013P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S40P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S40N045P064P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S40N045P064P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S40P058P013P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S40P058P013P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S40P058P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S40P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S40P062N035P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S40N062P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S40N062N059P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S41P065P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S41P065P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S41P044P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S41P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S41N015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S41P033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S41N033P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S41N033N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S41P067P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S41P067P006P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S41P067P046P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S41P013P031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S41P013N031P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S41N013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S41N013N068P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S41P048P063P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S41P048N063P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S41P046P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S41P046N008P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S41N046P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S41N046P069P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S41P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S41P056P033P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S41P056N033P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S41N056P068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S41N056N068P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S41P069P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S41P069N010P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S42P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S42P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S42N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S42N021N020P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S42P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S42N044P048P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S42P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S42P057P035P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S42P058P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S42N058P052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S42N058N052P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S42P057P019P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S42P057N019P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S42N057P069P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S42N057N069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S42P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S42P032P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S42P032P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S42P032P037P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S42P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S42N014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S42P016P037P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S42P016N037P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S42N016P066P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S42P033P063P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S42P033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S42P019P063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S42P019P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S42P019N009P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S42P060P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S42P060N057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S42P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S42P060N017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S42P062P036P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S42N062P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S43P043P019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S43P043P019P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S43N043P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S43N043P024P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S43P024P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S43P024P049P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S43N024P064P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S43P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S43P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S43N018P017P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S43P022P015P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S43P022P015P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S43P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S43P064P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S43N064P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S43P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S43P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S43N019P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S43N019N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S43P042P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S43P042N017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S43N042P021P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S43P023P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S43P023N057P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S43P066P052P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S43P066N052P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S43P066P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S43P052P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S43P052P035P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S43P052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S43P052N010P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S43P024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S43P024N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S44P026P029P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S44P054P035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S44P054P035P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S44P054P012P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S44P054N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S44P042P047P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S44P042P047P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S44P038P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S44P038N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S44N038P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S44N038N044P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S44P033P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S44P033N014P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S44P033P009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S44P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S44P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S44P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S44N035P037P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S44P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S44N037P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S44N037N017P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S44P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S44P015P059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S44P003P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S44P003P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S45P062P066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S45P062N066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S45P062psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S45P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S45N024P066P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S45P019P034P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S45P019P034P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S45N019P029P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S45N019N029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S45P017P045P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S45N017P019P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S45N017N019P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S45P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S45N008P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S45P027P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S45N027P009P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S45N027P009P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S45P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S45N062P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S45P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S45P008P065P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S45P010P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S45P010N060P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S45N010P005P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S45P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S45P010P012P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S45P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S45N066P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S45P065P059P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S45N065P046P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S45P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S46P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S46N058P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S46N058N007P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S46N069N037P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S46P034P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S46P034P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S46P034P014P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S46P034P014P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S46P019P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S46P019N050P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S46P046P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S46N046P017P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S46N046N017P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S46P067P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S46N067P064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S46N067N064P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S46P005P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S46P005N037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S46P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S46P056P037P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S46P056P037P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S46P056P065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S46P056P065P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S46P064P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S46P064P062P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S46P062P015P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S46P062P015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S46P062P068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S46P015P066P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S46P015P066P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S46N015P019P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S46N015N019P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S47P048P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S47P048P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S47P048N018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S47P027P048P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S47P027N048P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S47N027P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S47N027N051P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S47P047P013P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S47P047N013P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S47P047P035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S47P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S47P046N025P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S47P001P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S47P001N036P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S47P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S47P065N014P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S47N065P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S47P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S47N055P010P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S47P018P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S47P018N036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S47P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S47P018P012P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S47P018N012P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S47N018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S47P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S47P032N061P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S47N032P059P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S47P018P032P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S47N018P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S47P064P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S47P064P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S47P037P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S47N037P013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S48P012P063P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S48P012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S48P069P041P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S48P069N041P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S48N069P046P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S48P066P059P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S48P066P059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S48P066P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S48P066N059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S48P030P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S48P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S48N030P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S48N030P053P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S48P008P065P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S48N008P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S48P002P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S48P002P006P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S48P002P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S48P025P007P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S48P025N007P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S48N025P048P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S48N025P048P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S48P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S48N016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S48P041P033P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S48P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S48N061P033P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S49P028P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S49P028N019P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S49N028psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S49P015P032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S49P015N032P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S49N015P007P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S49P066P005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S49P066P056P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S49P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S49N020P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S49N020N016P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S49P050P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S49N050P055P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S49P015P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S49P015N054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S49N015P009P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S49N015N009P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S49P067P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S49P067N068P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S49N067P002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S49P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S49N016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S49N016N019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S49P065P022P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S49P065P032P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S49P014P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S49P014N065P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S49N014P068P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S49P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S50P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S50N002P004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S50N002N004P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S50P023P042P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S50P023N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S50N023P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S50N023P044P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S50P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S50P028N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S50N028P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S50N028N063P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S50P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S50N007P047P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S50P056P008P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S50N056P031P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S50N056P031P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S50P009P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S50P054P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S50P050P026P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S50P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S50N012P016P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S50N012N016P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S50P037P066P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S50P037N066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S50P000P010P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S50N000P008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S50P005P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S50P005N054P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S50P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S50P037N018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S50N037P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S50N037P012P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S50P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S51P068P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S51P068P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S51P061P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S51P061N064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S51P061P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S51P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S51P014P037P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S51P006P051P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S51P006N051P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S51P006P067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S51P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S51P018P014P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S51N018P007P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S51N018N007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S51P046P042P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S51N046P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S51N046N040P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S51P062P017P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S51P062N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S51P062P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S51P030P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S51P030P055P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S51N030P034P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S51N030N034P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S51P011P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S51P011P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S51P057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S51P057N013P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S51P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S51P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S51N028P012P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S52P049P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S52P049P056P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S52P003P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S52N003P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S52N003N046P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S52P013P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S52P013P030P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S52P013P003P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S52P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S52N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S52P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S52P014P015P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S52N014P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S52N014N007P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S52P004P036P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S52N004P005P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S52P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S52N033P032P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S52P064P012P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S52P064P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S52P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S52N009P024P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S52N009N024P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S52P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S52P051P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S52N051P033P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S53P029P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S53P029P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S53N029P019P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S53N029N019psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S53P018P010P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S53N018P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S53N018N054P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S53P019P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S53P019N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S53P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S53P019P018P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S53P066P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S53P066P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S53N066P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S53N066N053P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S53P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S53N033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S53N033N061P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S53P058P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S53P058P069P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S53P058P034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S53P062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S53P062N061P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S53P062P013P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S53P062N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S53P014P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S53P054P060P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S53P054N060P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S53P054P035P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S53P054N035P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S53P026P005P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S53P033P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S53P033N065P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S53P062P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S53N062P061P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S53P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S53N008P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S53N008N069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S54P036P044P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S54N036P004P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S54N036P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S54P024P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S54P024N023P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S54P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S54N069P040P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S54P032P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S54P032P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S54P048P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S54P020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S54P020N005P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S54N020P008P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S54P051P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S54N051P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S54P000P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S54N000P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S54N000P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S54P013P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S54P013N062P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S54N013P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S54P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S54N059P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S54N059N063P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S54P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S54P036P007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S54P036P007P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S54P036P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S54P012P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S54P012N066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S54N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S54N012N010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S54P034P006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S54N034P063P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S54P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S54N025P004P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S55P041P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S55P041P065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S55N041P003P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S55N041P003P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S55P067P010P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S55P035P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S55N035P058P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S55P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S55P067P035P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S55P067N035P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S55P067P062P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S55P067N062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S55P063P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S55P063P034P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S55P019P015P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S55P019P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S55N019P065P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S55P046P055P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S55P046N055P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S55P046P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S55P010P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S55P010N065P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S55N010P029P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S55P047P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S55P047P018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S55P054P000P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S55P054P035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S55P054N035P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S55P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S55N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S56P060P040P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S56N060P058P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S56N060P058P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S56P062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S56N062P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S56P037P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S56P037P065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S56P037P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S56P066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S56P066N013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S56P020P055P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S56P062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S56N062P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S56P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S56P060P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S56P056P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S56P056N066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S56P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S56N059P018P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S56P060P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S56P060N013P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S56P060P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S56P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S56P051P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S56P051P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S56N051P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S56N051N036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S56P049P026P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S56P049N026P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S57P020P005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S57P020N005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S57N020P019P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S57N020N019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S57P028P055P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S57N028P029P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S57P005P020P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S57P005P062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S57P005N062P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S57P054P060P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S57P054N060P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S57P054P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S57P054N014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S57P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S57N026P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S57P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S57N067P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S57N067N055P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S57P016P059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S57N016P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S57P068P035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S57P068N035P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S57P005P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S57P005N035P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S57P005P009P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S57P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S57P012P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S58P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S58N005P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S58N005N023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S58P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S58P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S58N002P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S58P015P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S58P015P036P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S58N015P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S58P035P034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S58P035P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S58N035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S58N035N013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S58P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S58P064P016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S58N064P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S58P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S58P030P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S58N030P015P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S58N030N015P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S58P035P014P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S58P035N014P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S58N035P014P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S58N035P014P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S58P013P069P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S58P013P069psss: std_logic_vector(   0 downto 0);
        signal cVar2S26S58P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S58P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S58P019P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S58P019P033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S58P019P069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S58P018P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S58N018P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S58P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S58P045P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S58P037P015P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S58N037P047P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S58N037N047P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S59P066P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S59P066N068P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S59P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S59P034P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S59P034P017P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S59P012P067P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S59P012P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S59N012P031P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S59N012P031P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S59P010P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S59P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S59P019P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S59P019P035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S59P019P034P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S59P019N034P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S59P055P061P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S59P067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S59P010P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S59P051P058P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S59P041P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S59P041P016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S59N041P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S59P008P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S59P008N019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S59N008P011P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S60P007P035P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S60P007N035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S60P007P057P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S60P012P048P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S60N012P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S60N012N004P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S60P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S60N015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S60P067P062P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S60P067N062P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S60N067P058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S60P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S60P014N016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S60P014P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S60P067P065P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S60P067P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S60P067P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S60P012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S60N012P059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S60P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S60N007P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S60P014P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S60P014N024P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S60P014P023P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S60P036P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S60P036N064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S60P069P034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S60P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S60P067P036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S60N067P051P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S60P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S60N010P031P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S60N010N031P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S60P033P060P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S60P033N060P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S60N033P055P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S61P065P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S61P065P055P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S61P065P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S61P065N030P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S61P067P064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S61P067N064psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S61N067P033P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S61N067P033P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S61P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S61N046P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S61P064P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S61P064P037P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S61P064N037P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S61P059P062P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S61P059N062P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S61P059P018P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S61P012P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S61P012P032P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S61P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S61P062P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S61N062P049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S61N062N049P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S61P067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S61P067N017P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S61N067P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S61P037P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S61P037N034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S61N037P069P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S61N037N069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S61P007P053P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S61P066P045P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S61P066P052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S61P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S61P067P066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S62P016P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S62P016N065P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S62N016P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S62N016N025P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S62P016P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S62P045P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S62N045P015P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S62N045N015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S62P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S62N039P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S62P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S62P033P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S62P033P015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S62P033P058P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S62P015P032P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S62P015P032P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S62N015P032P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S62N015N032P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S62P036P034P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S62P036P034P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S62P036P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S62P058P061P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S62P058P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S62N058P055P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S62P063P064P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S62P063P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S62P063N029P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S62P012P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S62P012P048P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S62N012P008P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S62P060P069P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S62P060P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S62P060N011P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S62P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S62P067N065P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S62N067P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S63P028P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S63P028P017P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S63P028P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S63P019P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S63N019P013P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S63P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S63P068P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S63P068N029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S63P040P030P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S63P040P030P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S63P034P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S63P034P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S63P034P069P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S63P017P069P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S63N017P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S63N017N045P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S63P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S63P025P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S63P025N062P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S63N025P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S63N025N065P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S63P010P055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S63P010P055P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S63P010P024P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S63P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S63P030P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S63P030N013P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S63P030P009P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S63P034P008P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S63P034P008P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S63N034P025P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S64P030P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S64P030P067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S64P062P047P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S64P062N047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S64P062P006P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S64P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S64P060P062P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S64P032P060P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S64P032N060P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S64P065P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S64P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S64P013P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S64N013P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S64N013N056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S64P011P060P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S64P011N060P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S64N011N014P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S64P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S64N060P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S64P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S65P037P024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S65P019P037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S65P019P037P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S65N019P007P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S65P003P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S65P003N065P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S65N003P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S65P012P056P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S65P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S65N011P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S65P036P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S65P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S65N034P069P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S65P007P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S65P007N016P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S65N007P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S65P036P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S65P036N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S65P036psss: std_logic_vector(   0 downto 0);
        signal cVar2S22S65P004P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S65N004P037P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S65P039P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S65P039N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S65N039P021P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S65P037P069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S66P058P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S66P058N022P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S66P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S66P007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S66P007N005P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S66P007P013P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S66P026P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S66P039P048P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S66P039P048P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S66P039P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S66P032P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S66P032N019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S66N032psss: std_logic_vector(   0 downto 0);
        signal cVar2S15S66P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S66N011P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S66P052P059P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S66P052P059P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S66P052P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S66P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S66P068P018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S66N068P036P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S66P036P037P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S66P036P037P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S66P036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S66P036N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S66P017P051P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S66P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S66N043P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S66P050P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S66P050P011P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S66P050P027P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S66P050N027P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S67P028P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S67P028P034P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S67P028P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S67P028P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S67P035P009P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S67N035P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S67N035N020P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S67P035P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S67P035N012P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S67P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S67P010N019P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S67N010P027P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S67P033P019P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S67P033P019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S67N033P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S67N033N057P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S67P009P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S67P009N068P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S67P010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S67P010N032P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S67P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S67N068P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S67P007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S67P007N005P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S67P007P013P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S67P026P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S67P026P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S67P039P023P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S67P039P023P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S67P039P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S68P062P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S68P062P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S68P062N019P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S68P018P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S68P018N060P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S68P018P023P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S68P018N023P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S68P066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S68P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S68N034P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S68P051P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S68P051N066P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S68P051P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S68P004P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S68P067P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S68P067N049P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S68N067psss: std_logic_vector(   0 downto 0);
        signal cVar2S18S68P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S68P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S68P023N005P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S68P010P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S68P001P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S68P001N068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S68N001P066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S68N001P066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S68P062P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S68P062P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S68P062N015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S68P005P042P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S68P005P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S68P044P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S68N044P023P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S68N044P023P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S69P063P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S69P063N065P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S69P063P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S69P063N005P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S69P065P019P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S69N065P035P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S69N065N035P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S69P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S69N059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S69P009P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S69P009P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S69N009P036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S69N009N036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S69P012P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S69P012N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S69N012P026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S69P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S69P040N002P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S69N040P038P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S69P025P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S69P025N068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S69N025P039P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S69P068P066P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S69P068P016P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S69P051P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S69P051P064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S69N051P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S69P030P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S69P030N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S69N030P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S69N030N032P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S69P068P051P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S69P051P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S69P051N026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S69P051P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S69P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S69N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S69N024N025P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S69P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S69N016P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S69P042P067P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S69P042N067P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S69P042P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S43S69P042N021P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S70P020P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S70P020N047P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S70P047P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S70P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S70P047N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S70P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S70P023P040P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S70P023N040P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S70P039P069P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S70P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S70N001P018P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S70N001N018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S70P020P052P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S70P020P052P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S70P020P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S70P069P012P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S70N069P029P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S70N069N029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S70P048P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S70P048N037P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S70P048P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S70P020P032P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S70P020P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S70N020P065P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S70P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S70N042P037P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S71P016P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S71P016P060P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S71P016P055P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S71P016P055P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S71P019P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S71N019P063P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S71P033P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S71P033N021P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S71P014P007P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S71P014P007P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S71N014P016P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S71N014N016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S71P013P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S71P013N019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S71P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S71P028P019P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S71P028P019P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S71N028P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S71N028N013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S71P034P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S71P034N006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S71P034P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S71P055P004P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S71P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S71N034P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S71N034N012P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S71P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S71P042P013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S71P042P013P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S71P009P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S71N009P000P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S71P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S71P018P047P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S72P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S72P013P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S72N013P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S72N013N006P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S72P054P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S72P054P018P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S72N054P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S72N054N060P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S72P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S72P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S72P006P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S72P006P017P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S72P012P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S72P012P010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S72P020P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S72N020P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S72N020P016P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S72P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S72N031P053P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S72P059P057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S72P059N057P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S72P059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S72P039P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S72P039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S72P039N003P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S72P016P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S72P016P033P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S73P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S73P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S73N065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S73N065N068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S73P018P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S73P018P005P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S73N018P059P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S73N018P059P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S73P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S73N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S73N011N009P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S73P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S73N066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S73P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S73N009P067P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S73N009P067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S73P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S73N048P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S73N048N051P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S73P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S73N002P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S73N002N000P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S73P028P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S73P028N043P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S73N028P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S73N028N067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S73P013P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S73N013P047P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S73P066P064P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S73N066P019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S73P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S74P049P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S74P049N058P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S74N049P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S74N049N050P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S74P055P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S74P055N015P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S74N055P057P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S74P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S74N010P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S74N010N008P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S74P026P037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S74P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S74N028P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S74N028N051P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S74P057P011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S74P057P066P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S74P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S74P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S74N006P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S74P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S74P010N052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S74N010P054P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S74P011P026P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S74P011P010P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S74P018P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S74P018N066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S75P037P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S75P037N048P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S75P045P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S75P045P014P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S75P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S75P056P031P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S75P056N031P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S75P056P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S75P056N032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S75P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S75N011P067P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S75P007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S75N007P016P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S75P065P037P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S75P065N037P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S75N065P030P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S75N065N030P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S75P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S75P009P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S75N009P014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S75N009N014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S75P017P068P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S75P017P068P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S75P017P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S75P017P063P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S75P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S75P019N012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S75P019P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S75P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S75N035P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S75N035P067P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S75P055P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S75P055P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S75P055N068P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S76P033P065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S76P033N065P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S76N033P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S76P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S76P052N029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S76N052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S76P026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S76P026N018P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S76P010P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S76P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S76P037P035P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S76P037N035P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S76P066P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S76N066P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S76P036P008P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S76P036P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S76P001P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S76P001N068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S76N001P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S76P032P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S76P032P037P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S76N032P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S76P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S76N025P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S76P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S76P031P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S76P031N030P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S76P035P053P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S76P035P053P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S76P035P033P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S76P015P011P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S76P015N011P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S76N015P010P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S76N015N010P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S77P064P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S77P064P018P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S77P064P000P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S77P064P000P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S77P051P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S77P051N018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S77P014P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S77P014P030P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S77N014P011P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S77N014P011P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S77P013P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S77P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S77N011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S77N011N015P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S77P000P047P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S77P015P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S77P015N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S77N015P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S77N015N001P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S77P069P060P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S77P060P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S77P060N067P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S77P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S77P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S77P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S77N037P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S77P007P006P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S77P007P006P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S77P007P057P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S78P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S78N015P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S78N015N029P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S78P034P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S78P034P067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S78P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S78P034N012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S78P062P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S78P062N020P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S78N062P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S78P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S78P013P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S78P013P015P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S78P026P009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S78P026P009P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S78P056P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S78P018P007P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S78P018P063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S78P017P056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S78P017N056P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S78N017P065P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S78P051P057P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S78P051N057P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S78P051P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S78P058P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S78P028P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S78P028N011P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S78N028P047P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S78P014P019P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S78P014N019P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S78N014P045P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S78N014N045P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S78P013P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S79P046P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S79N046P057P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S79N046N057psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S79P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S79N056P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S79P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S79N009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S79N009P050P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S79P058P034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S79P019P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S79P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S79N050P029P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S79P015P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S79P015P003P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S79P015P055P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S79P015N055P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S79P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S79N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S79N029N027P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S79P065P069P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S79N065P037P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S79P029P017P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S79P032P059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S79P032P059P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S79P032P059P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S79P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S79N057P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S79P015P059P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S79P015P063P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S80P032P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S80P032P010P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S80P032P061P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S80P014P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S80P014N031P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S80P014P031P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S80P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S80N016P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S80P012P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S80P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S80N044P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S80N044P011P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S80P031P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S80N031P032P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S80P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S80P061P031P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S80P061P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S80P032P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S80N032P058P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S80N032P058P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S80P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S80P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S80P016N068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S80P026P047P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S80P026P053P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S80P034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S80P034P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S80N034P062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S80N034P062P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S80P053P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S80P040P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S80P040N062P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S80N040P055P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S80N040N055P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S80P060P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S80P060N069P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S80N060P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S81P029P030P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S81N029P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S81N029P054P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S81P013P065P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S81N013P052P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S81N013P052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S81P069P061P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S81N069P062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S81P069P026P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S81P069P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S81P027P045P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S81P027P045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S81P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S81N010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S81P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S81N030P015P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S81N030P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S81P012P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S81P012N058P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S81P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S81N027P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S81N027N017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S81P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S81N017P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S81N017N067P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S81P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S81N033P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S81N033N065P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S81P036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S81N036P062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S81P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S81N021P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S81N021P066P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S81P047P007P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S81P047P007P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S81P047P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S81P047N026P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S82P044P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S82N044P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S82N044P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S82P035P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S82P035P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S82P035N007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S82P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S82P067P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S82P067N029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S82N067P019P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S82P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S82P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S82P018P068P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S82P013P011P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S82P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S82P019P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S82N019P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S82N019P069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S82P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S82N005P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S82P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S82P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S82P056P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S82P056P052P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S82P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S82P000P044P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S83P006P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S83N006P060P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S83N006N060P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S83P024P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S83P024P049P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S83P024P002P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S83P003P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S83P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S83P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S83N029P067P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S83N029P067P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S83P062P067P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S83P062N067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S83P062P066P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S83P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S83P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S83P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S83N069P010P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S83P063P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S83P063N005P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S83N063P064P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S83P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S84P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S84P035P067P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S84P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S84N001P036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S84N001P036P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S84P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S84P068P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S84P068P036P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S84P068P037P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S84P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S84P030N057P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S84N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S84P065P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S84P065N058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S84N065P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S84N065N036P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S84P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S84P067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S84P067N037P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S84P059P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S84N059P034P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S84P046P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S84P046P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S84P049P046P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S84N049P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S84N049N046P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S84P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S84N069P018P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S84P012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S84P012P069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S84P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S84P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S84P005P051P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S84P005P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S84P005N039P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S84P059P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S84N059P046P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S84N059N046P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S85P021P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S85P021N058P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S85P021P010P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S85P065P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S85P065N011P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S85N065P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S85N065N012P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S85P017P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S85P017P004P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S85N017P069P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S85N017P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S85P014P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S85P014N010P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S85N014P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S85P007P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S85P007P050P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S85P026P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S85N026P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S85N026N006P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S85P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S85P034P036P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S85P034P036P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S85P034P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S85P013P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S85P013N063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S85N013P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S85P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S85P034P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S85P034N069P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S85N034P068P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S85N034N068P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S85P014P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S85P014P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S85P002P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S85P002N047P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S85P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S85N050P017P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S85N050N017P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S85P052P058P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S85P052P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S85P052N013P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S86P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S86N056P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S86N056N003P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S86P068P013P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S86P068P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S86N068P066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S86P006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S86P006N005P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S86P006P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S86P006N001P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S86P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S86N020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S86P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S86P037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S86P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S86N011P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S86N011N061P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S86P033P057P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S86P033P057P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S86P033P013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S86P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S86P020P005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S86P020P005P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S86P020P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S86P059P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S86N059P012P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S86P063P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S86P039P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S86P039N059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S86P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S86P029N050P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S86P029P026P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S86P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S86P027N050P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S86N027P048P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S86N027P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S86P065P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S86P065N036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S86N065P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S86N065N047P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S87P009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S87P009P008P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S87N009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S87N009N069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S87P009P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S87P009P050P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S87P009N050P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S87N064P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S87P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S87N036P019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S87P035P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S87P035N067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S87N035P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S87P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S87N057P037P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S87N057N037P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S87P042P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S87N042P056P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S87N042N056P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S87P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S87N029P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S87P010P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S87N010P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S87N010N026P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S87P018P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S87P018N056P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S87N018P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S87N018N021P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S87P032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S87N032P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S87N032N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S87P018P037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S87P018P037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S87P018P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S87P018N036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S87P062P037P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S87P062N037P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S87P062P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S88P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S88P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S88P019N015P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S88P058P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S88P058N063P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S88N058P054P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S88P003P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S88P003P015P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S88P003P058P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S88P035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S88P035P069P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S88N035P019P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S88N035N019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S88P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S88N002P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S88N002N042P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S88P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S88N044P004P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S88P048P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S88P048N033P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S88P048N031P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S88P017P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S88P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S88P011P028P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S88P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S88N042P015P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S88N042N015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S88P012P017P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S88P012N017P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S88P012P041P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S88P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S88N036P018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S88P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S89P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S89N034P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S89N034P026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S89P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S89N036P020P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S89N036N020P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S89P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S89N064P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S89N064N066P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S89P064P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S89P064P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S89P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S89N046P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S89N046N033P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S89P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S89N029P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S89N029P046P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S89P023P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S89P023N006P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S89P048P046P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S89P048P062P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S89P027P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S89P027N032P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S89P027P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S89P027N051P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S89P010P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S89P036P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S89P036N056P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S89N036P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S89N036N016P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S89P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S89N036P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S89P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S90P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S90N036P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S90N036N035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S90P000P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S90P000N034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S90N000P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S90P023P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S90P023N027P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S90P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S90P069P060P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S90P069N060P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S90P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S90P066P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S90N066P016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S90P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S90P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S90N040P002P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S90N040P002P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S90P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S90P039P066P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S90N039P020P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S90P051P055P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S90N051P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S90P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S90N032P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S90P062P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S90N062P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S90P015P034P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S90N015N057P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S91P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S91N025P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S91N025P035P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S91P006P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S91P006N027P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S91N006psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S91P000P020P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S91P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S91N015P009P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S91P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S91P058P066P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S91P058N066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S91P060P069P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S91P060P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S91N060P008P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S91N060N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S91P062P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S91N062P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S91P015P034P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S91N015N057P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S91P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S91P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S91P002P038P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S91P002P038P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S91P002P013P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S91P002N013P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S91P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S91N004P019P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S91P010P022P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S92P002P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S92P002P041P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S92P002P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S92P002N040P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S92P058P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S92P058P066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S92N058P002P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S92N058N002P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S92P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S92P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S92P034P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S92P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S92N057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S92P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S92P061P058P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S92P061P058P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S92N061P062P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S92N061N062P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S92P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S92P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S92N052P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S92P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S92P063P037P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S92P054P010P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S92P054P010P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S92P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S92P061N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S92N061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S92P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S92N053P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S92P021P036P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S92P021N036P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S92P021P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S92P041P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S92P041N005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S93P006P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S93P006N013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S93N006P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S93N006P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S93P054P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S93N054P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S93N054N050P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S93P037P051P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S93P037N051P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S93N037P068P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S93N037P068P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S93P013P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S93P016P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S93P016N055P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S93P031P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S93P031P035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S93P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S93P057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S93P057N031P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S93N057P033P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S93N057N033P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S93P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S93N052P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S93P026P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S93P026N050P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S93P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S93N008P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S93N008N005P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S93P008P035P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S93P008P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S93P068P022P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S93P068P022P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S93P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S93N040P037P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S93N040N037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S94P043P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S94P043N061P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S94P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S94P015N068P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S94P065P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S94P065P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S94P037P057P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S94P037N057P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S94N037P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S94P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S94N066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S94P015P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S94P015P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S94P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S94P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S94P014P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S94N014P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S94P008P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S94N008P048P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S94N008P048P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S94P058P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S94P058N066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S94P058P061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S94P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S94N069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S94N069P018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S94P022P016P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S94P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S94P031P054P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S94P031N054P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S94P034P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S94N034P004P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S94N034N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S94P061P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S94P061N000P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S94P061P067P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S94P000P037P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S94P000P033P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S95P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S95P025N046P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S95N025P051P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S95N025N051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S95P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S95N057P019P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S95P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S95N002P033P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S95N002N033P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S95P000P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S95P000N037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S95N000P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S95N000N052P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S95P015P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S95P015N033P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S95P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S95P015N011P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S95P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S95P014P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S95P014N058P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S95P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S95N022P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S95P066P040P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S95P066P040P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S95P066P014P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S95P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S95N012P023P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S95P033P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S95P033N026P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S95P027P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S95P027P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S95N027P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S95N027P002P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S95P000P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S95P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S95N049P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S95N049N010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S95P001P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S95P001P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S95N001P028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S96P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S96N014P060P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S96N014P060P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S96P022P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S96P022N015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S96N022P049P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S96N022N049P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S96P018P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S96P018N061P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S96N018P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S96N018N030P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S96P035P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S96P035P017P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S96P062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S96P062N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S96P062P063P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S96P007P031P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S96P007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S96P007N047P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S96P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S96P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S96N059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S96P067P014P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S96P067N014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S96N067P009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S96P050P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S96P050N013P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S96P010P048P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S96P010N048P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S96N010P047P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S96N010P047P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S96P036P054P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S96P036P054P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S96P036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S96P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S96N065P030P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S97P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S97P008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S97P013P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S97P013P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S97N013psss: std_logic_vector(   0 downto 0);
        signal cVar2S5S97P055P058P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S97P055N058psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S97P055P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S97P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S97P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S97P013P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S97P013P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S97P066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S97P066P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S97P066N013P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S97P028P010P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S97P028N010psss: std_logic_vector(   0 downto 0);
        signal cVar2S18S97P028P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S97P064P033P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S97P064P033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S97P038P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S97P038N064P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S97P056P065P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S97P056P065P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S97N056P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S97P017P064P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S97P017P064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S97P017P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S97P017N057P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S97P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S98P018P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S98P018N065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S98N018P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S98N018N059P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S98P066P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S98P051P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S98N051psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S98P030P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S98N030P034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S98P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S98N014P054P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S98N014N054P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S98P033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S98P033N012P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S98P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S98N058P006P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S98P014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S98N014P003P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S98P007P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S98P007N064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S98N007P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S98P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S98N062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S98P007P037P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S98P007P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S98P054P057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S98P054P057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S98N054P031P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S98P026P066P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S99P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S99N044P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S99N044N047P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S99P025P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S99P025N066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S99N025P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S99P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S99P062P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S99P062N057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S99N062P034P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S99N062P034P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S99P001P011P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S99P001P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S99N001P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S99N001N059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S99P020P002P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S99P026P062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S99P026N062P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S99P020P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S99P020P060P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S99P020P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S99P069P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S99P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S99N013P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S99N013N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S99P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S99P025P057P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S99P025N057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S99P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S99P025P004P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S99P025N004P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S99N025P012P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S99P057P017P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S99P057P030P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S99P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S99N015P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S100P064P005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S100P064P005P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S100P064P068P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S100P044P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S100P044N035P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S100N044P038P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S100N044N038psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S100P029P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S100P029N037P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S100N029P034P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S100N029P034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S100P064P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S100P064P060P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S100P064P037P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S100P061P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S100P061P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S100N061P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S100N061N065P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S100P052P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S100P052P050P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S100N052P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S100P058P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S100P058N001P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S100N058P057P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S100P062P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S100P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S100N027P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S100N027N037P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S100P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S100P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S100P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S100P052N029P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S100N052P029P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S100P023P005P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S100P023P005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S100P023P042P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S100P012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S101P000P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S101P000N069P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S101N000P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S101N000P057P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S101P027P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S101P027N060P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S101P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S101P033P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S101P033N003P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S101P058P010P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S101P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S101N015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S101N015N017P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S101P029P062P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S101P029P062P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S101P029P054P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S101P062P033P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S101P062N033P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S101N062P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S101P021P006P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S101P021N006P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S101P018P064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S101P018N064P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S101N018P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S101N018N033P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S101P010P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S101P058P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S101P058N016P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S101P058P061P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S101P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S102P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S102N059P065P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S102N059P065P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S102P009P068P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S102P055P056P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S102P055P056P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S102N055P013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S102N055N013P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S102P011P013P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S102P011P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S102P011P003P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S102P017P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S102P017N063P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S102N017P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S102N017P069P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S102P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S102P030N057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S102N030P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S102P056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S102P056N012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S102N056P044P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S102P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S102N062P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S102P034P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S102P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S102N065P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S102P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S102P008N026P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S102N008P011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S102P058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S102N058P031P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S103P017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S103P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S103P045P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S103P045P038P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S103P045P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S103P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S103P068P037P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S103P007P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S103P007N050P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S103P007P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S103P007N018P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S103P052P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S103N052P063P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S103P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S103P012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S103P012P013P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S103N012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S103N012N017P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S103P010P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S103P010P018P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S103P067P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S103P067P032P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S103P067P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S103P067N059P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S103P031P007P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S103P031N007P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S103P031P010P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S104P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S104N009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S104P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S104N013P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S104N013N034P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S104P057P031P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S104P049P026P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S104P049P026P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S104P049P007P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S104P049N007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S104P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S104N047P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S104P057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S104P057P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S104P057P019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S104P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S104N062P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S104P005P003P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S104P005P031P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S104P040P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S104P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S104P066P012P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S105P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S105P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S105P055P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S105P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S105P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S105N031P032P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S105N031N032P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S105P028P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S105P028P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S105N028P026P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S105N028N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S105P028P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S105P028N057P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S105P028P030P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S105P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S105P014P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S105P051P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S105P051P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S105P003P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S105P003N017P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S105P003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S105P003N005P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S105P004P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S105P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S105N067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S105P050P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S105N050P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S105P021P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S105P031P029P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S105P031P054P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S105P031N054P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S106P008P037P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S106P008N037P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S106N008P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S106N008N019P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S106P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S106N024P026P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S106P010P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S106P010P017P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S106P051P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S106N051P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S106P023P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S106P023N006P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S106N023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S106N023P042P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S106P060P063P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S106P060P063P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S106N060P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S106N060N065P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S106P002P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S106P002N011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S106N002P033P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S106N002N033P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S106P033P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S106P059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S106P059P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S106P058P059P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S106P058N059P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S106P058P014P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S106P069P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S106N069P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S106N069N061P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S107P061P037P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S107P061P037P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S107P061P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S107P049P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S107P012P032P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S107P012P032P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S107P012P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S107P012N056P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S107P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S107N026P009P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S107P033P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S107P033N003P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S107P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S107N032P058P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S107P010P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S107P010P013P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S107P030P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S107N030P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S107N030P017P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S107P003P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S107N003P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S107P035P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S107P035N055P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S107N035P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S107N035N009P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S107P066P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S107N066P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S107N066N024P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S107P053P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S107P053N030P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S107P023P006P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S107P023N006P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S107N023P059P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S107P026P057P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S108P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S108P030P057P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S108P030P029P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S108P029P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S108P029N008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S108N029P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S108N029N061P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S108P054P015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S108P054N015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S108N054P057P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S108P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S108P056P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S108P056P033P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S108P056P010P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S108P061P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S108N061P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S108P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S108P060P059P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S108P060P004P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S108N060P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S108P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S108N061P014P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S108N061P014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S108P069P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S108P069N034P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S108N069P063P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S108P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S108N016P015P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S108P043P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S108P043N008P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S108P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S108N065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S108N065N018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S108P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S108N057P013P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S108P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S108N030P051P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S108P017P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S108P017N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S108N017P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S109P057P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S109P057N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S109N057P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S109N057P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S109P052P067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S109P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S109N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S109N031N029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S109P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S109P009P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S109P009N063P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S109N009P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S109P013P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S109P013N058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S109N013P052P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S109N013N052P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S109P008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S109P008P011P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S109N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S109P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S109N003P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S109N003N007P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S109P042P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S109P042N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S109N042P006P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S109P047P024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S109P047N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S109N047P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S109P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S110P050P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S110P050P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S110P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S110P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S110N015P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S110P016P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S110P016N065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S110N016P063P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S110N016P063P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S110P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S110N024P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S110N024N027P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S110P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S110N036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S110N036P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S110P051P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S110P051N019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S110N051P046P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S110P019P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S110P019N028psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S110P019P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S110P019N068P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S110P009P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S110P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S110P036P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S110P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S110N034P048P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S111P015P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S111N015P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S111N015P058P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S111P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S111N065P011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S111P034P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S111N034P003P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S111N034N003P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S111P020P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S111P020N057P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S111P020P015P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S111P020P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S111P006P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S111N006P001P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S111P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S111P065P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S111P065N018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S111P049P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S111P049N067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S111N049P017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S111N049N017P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S111P004P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S111P004N017P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S111N004P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S111P042P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S111P061P014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S111P061P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S112P009P033P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S112P009P033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S112P009P065P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S112P009N065P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S112P012P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S112P012N009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S112N012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S112N012P069P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S112P066P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S112P066N049P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S112P066P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S112P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S112N063P015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S112N063N015P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S112P024P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S112P024N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S112P069P061P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S112P061P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S112P061N063P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S112P061P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S112P067P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S112P067N051P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S112P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S112N024P035P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S112N024N035P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S112P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S112N037P063P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S112P013P061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S112P013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S112P057P011P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S112P057P011P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S112P057P059P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S112P057N059P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S112P001P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S112P001P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S112N001P065P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S112N001N065P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S112P055P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S113P057P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S113P057P055P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S113P057P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S113P057N012P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S113P055P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S113P055N029P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S113N055P008P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S113N055N008P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S113P052P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S113P052P016P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S113P057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S113P057N013P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S113P057P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S113P030P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S113P030N056P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S113N030P062P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S113N030P062P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S113P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S113N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S113N012N010P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S113P064P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S113P064N032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S113N064P034P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S113N064N034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S113P016P052P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S113P016N052P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S113P016P035P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S113P016N035P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S113P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S113P037P032P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S113P037N032P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S113N037P033P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S113N037N033P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S113P066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S113P034P061P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S113P034P061P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S113P034P016P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S113P034N016P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S113P064P007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S113P064P007P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S113P064P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S113P064N068P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S43S113P030P008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S44S113P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S114P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S114P049P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S114P049N009P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S114N049P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S114N049P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S114P013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S114P013N003P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S114P013P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S114P033P059P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S114N033P028P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S114P007P059P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S114P007N059P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S114N007P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S114N007N035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S114P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S114N029P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S114P013P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S114P013N028P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S114P013P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S114P021P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S114P021P011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S114P021P010P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S114P033P032P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S114P033N032P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S114P033P032P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S114P033P032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S114P034P040P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S114P034P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S114P034N017P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S114P056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S114P056N012P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S114P056P012P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S114P013P060P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S114N013P016P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S114N013P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S114P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S114P007P062P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S114P017P015P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S114P017P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S115P028P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S115P028N019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S115N028P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S115N028N037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S115P016P037P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S115P016P037P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S115N016P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S115P011P013P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S115P011N013P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S115P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S115P011P066P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S115P019P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S115P019N036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S115N019P062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S115P036P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S115P036N030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S115P036P053P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S115P032P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S115P032N069P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S115N032P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S115P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S115N006P016P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S115N006N016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S115P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S115N045P002P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S115N045N002P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S115P007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S115P007N047P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S115P007P059P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S115P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S115N061P037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S115P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S115N005P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S115P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S115N066P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S115P059P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S115N059P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S115N059N028P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S115P033P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S115P033N009P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S115N033P028P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S115P058P032P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S115P058N032P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S116P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S116N026P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S116N026N006P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S116P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S116N046P069P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S116N046P069psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S116P048P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S116P048N028P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S116P048P006P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S116P048N006P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S116P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S116N012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S116P035P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S116P015P036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S116P015N036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S116P015P065P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S116P015N065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S116P002P067P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S116P002N067P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S116P002N015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S116P017P037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S116P017P037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S116P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S116P017P016P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S116P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S116N012P017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S116N012N017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S116P045P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S116P045N047P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S116N045P043P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S116P060P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S116N060P034P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S116P010P034P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S116P010N034P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S116P010P013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S116P005P047P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S116P058P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S116P058N008P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S116N058P008P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S116N058P008P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S116P033P036P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S116P033N036P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S117P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S117N016P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S117P035P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S117N035P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S117P065P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S117N065P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S117P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S117P018P051P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S117N018P049P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S117N018N049P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S117P031P007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S117P031P007P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S117N031P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S117N031N035P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S117P035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S117P035P037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S117P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S117P010P002P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S117P010P002P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S117P010P054P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S117P010N054P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S117P024P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S117N024P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S117P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S117P019P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S117P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S117N069P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S117P068P009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S117P068P009P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S117P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S117P016N069P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S117P016P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S117P016P026P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S117N016P034P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S117N016P034P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S118P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S118P006P061P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S118P006P061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S118P006P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S118P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S118P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S118N011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S118P068P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S118P068P036P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S118P068P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S118P068N018P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S118P066P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S118P066P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S118N066P030P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S118P048P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S118P048N029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S118P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S118P048P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S118P048P066P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S118N048P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S118N048N045P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S118P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S118N063P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S118P006P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S118P006P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S118P006N028P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S118P008P033P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S118P008N033P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S118P008P060P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S118P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S118N013P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S119P001P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S119P001P026P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S119P052P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S119P036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S119N036P050P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S119N036N050P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S119P034P019P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S119N034P069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S119N034N069P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S119P036P068P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S119P036N068P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S119P036P053P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S119P024P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S119P024N047P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S119N024P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S119N024N052P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S119P057P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S119N057P009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S119P060P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S119P060P066P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S119P060P057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S119P059P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S119P059P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S119P035P034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S119P035P034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S119P035P009P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S119P063P067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S119P063P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S119P063P069P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S119P063N069P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S119P063P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S119P063N036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S119P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S119P019P015P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S119N019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S120P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S120P017P019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S120P017P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S120P017N060P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S120P068P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S120P068P036P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S120P018P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S120P018N069psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S120P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S120P018P017P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S120P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S120N052P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S120N052P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S120P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S120P016N068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S120P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S120P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S120P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S120P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S120N027P010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S120N027P010P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S120P056P003P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S120N056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S120N056P012P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S120P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S120N048P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S120P024P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S120P061P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S120P061N019P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S120N061P059P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S120N061P059P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S120P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S120N017P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S120P017P063P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S120P017P061P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S120P017N061P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S120P035P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S120N035P063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S121P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S121N056P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S121N056N008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S121P056P048P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S121P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S121P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S121P015P062P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S121P004P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S121P004N025P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S121N004P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S121P051P009P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S121P051N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S121N051P027P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S121P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S121N067P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S121N067N016P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S121P048P046P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S121N048P067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S121N048N067P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S121P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S121P066P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S121P066P016P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S121P066P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S121P066N013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S121P067P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S121P060P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S121P060N032P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S121N060P032P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S121P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S121P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S121N062P018P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S121P063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S121P063N011P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S122P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S122P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S122N050P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S122P061P048P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S122P061P048P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S122P061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S122P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S122P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S122P004P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S122P004N025P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S122N004P027P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S122N004N027P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S122P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S122P041P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S122P041N036P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S122P041P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S122P011P036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S122N011P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S122P001P018P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S122P001N018P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S122P007P029P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S123P044P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S123P044P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S123N044P058P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S123N044N058psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S123P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S123N004P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S123P065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S123P065P069P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S123P065P069P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S123P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S123N030P015P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S123N030N015P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S123P013P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S123P013P011P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S123P013N011P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S123P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S123P005P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S123P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S123P064P004P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S123P064N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S123P064P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S123P064P067P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S123P018P058P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S123P018P058P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S123P018P058P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S123P018N058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S123P011P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S123P011N069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S123N011P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S123N011N056P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S123P062P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S123P015P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S123P015N034P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S123P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S123P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S123N000P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S123N000P061P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S123P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S123P010N028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S39S123N010P042P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S40S123N010P042P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S41S123P014P034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S42S123P014N034P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S43S123N014P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S124P040P012P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S124P040P012P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S124P040P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S124P042P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S124N042P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S124P003P066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S124P003N066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S124P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S124P017P037P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S124N017P033P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S124N017N033P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S124P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S124N015P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S124N015P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S124P067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S124P009P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S124P009N058P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S124N009P020P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S124N009N020P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S124P010P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S124N010P046P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S124P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S124N040P037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S124P052P005P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S124P052P059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S124P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S124P012P014P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S124P040P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S124P040N025P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S124P025P023P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S124P025P047P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S125P067P069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S125P067N069psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S125P067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S125P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S125P036N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S125P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S125P035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S125P035N037P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S125N035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S125P052P013P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S125P052N013psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S125P052P050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S125P030P031P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S125N030P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S125N030N004P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S125P067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S125P067P066P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S125N067P065P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S125N067N065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S125P016P024P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S125P016P024P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S125N016P007P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S125P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S125N019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S125P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S125P011P009P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S125P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S125P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S125P056P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S125P017P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S125P017N059P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S125N017P003P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S125P008P033P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S125P008N033P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S125P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S125N054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S125P056P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S126P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S126N019P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S126P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S126P067P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S126P067N064P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S126P067P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S126P067N045P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S126P062P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S126P062P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S126P062P063P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S126P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S126N064P019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S126P063P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S126P063N019P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S126N063P033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S126P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S126P014P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S126P014P013P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S126P045P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S126P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S126P043N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S126N043P022P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S126P068P065P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S126P068P058P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S126P068N058P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S126P062P068P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S126P062N068P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S126N062P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S126N062N015P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S126P047P007P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S126P047P019P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S126P024P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S126P024P019P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S126N024P035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S126N024N035P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S127P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S127P000P044P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S127P067P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S127P067P025P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S127P067P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S127P067N066P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S127P036P051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S127P036N051P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S127P036P030P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S127P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S127N026P067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S127P007P000P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S127P007N000psss: std_logic_vector(   0 downto 0);
        signal cVar2S13S127P007P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S127P005P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S127P008P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S127P008N060P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S127N008P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S127N008N052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S127P053P017P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S127P053N017P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S127P053P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S127P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S127P015P063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S127P015N063P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S127P063P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S127P063P067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S127P063P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S127P063N019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S127P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S127N052P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S127P003P015P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S127P003N015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S127N003P043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S127P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S127P035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S38S127N035P069nsss: std_logic_vector(   0 downto 0);
        signal oVar1S0: std_logic_vector(   0 downto 0);
        signal oVar1S1: std_logic_vector(   0 downto 0);
        signal oVar1S2: std_logic_vector(   0 downto 0);
        signal oVar1S3: std_logic_vector(   0 downto 0);
        signal oVar1S4: std_logic_vector(   0 downto 0);
        signal oVar1S5: std_logic_vector(   0 downto 0);
        signal oVar1S6: std_logic_vector(   0 downto 0);
        signal oVar1S7: std_logic_vector(   0 downto 0);
        signal oVar1S8: std_logic_vector(   0 downto 0);
        signal oVar1S9: std_logic_vector(   0 downto 0);
        signal oVar1S10: std_logic_vector(   0 downto 0);
        signal oVar1S11: std_logic_vector(   0 downto 0);
        signal oVar1S12: std_logic_vector(   0 downto 0);
        signal oVar1S13: std_logic_vector(   0 downto 0);
        signal oVar1S14: std_logic_vector(   0 downto 0);
        signal oVar1S15: std_logic_vector(   0 downto 0);
        signal oVar1S16: std_logic_vector(   0 downto 0);
        signal oVar1S17: std_logic_vector(   0 downto 0);
        signal oVar1S19: std_logic_vector(   0 downto 0);
        signal oVar1S20: std_logic_vector(   0 downto 0);
        signal oVar1S21: std_logic_vector(   0 downto 0);
        signal oVar1S22: std_logic_vector(   0 downto 0);
        signal oVar1S23: std_logic_vector(   0 downto 0);
        signal oVar1S24: std_logic_vector(   0 downto 0);
        signal oVar1S25: std_logic_vector(   0 downto 0);
        signal oVar1S26: std_logic_vector(   0 downto 0);
        signal oVar1S27: std_logic_vector(   0 downto 0);
        signal oVar1S28: std_logic_vector(   0 downto 0);
        signal oVar1S29: std_logic_vector(   0 downto 0);
        signal oVar1S30: std_logic_vector(   0 downto 0);
        signal oVar1S31: std_logic_vector(   0 downto 0);
        signal oVar1S32: std_logic_vector(   0 downto 0);
        signal oVar1S33: std_logic_vector(   0 downto 0);
        signal oVar1S34: std_logic_vector(   0 downto 0);
        signal oVar1S35: std_logic_vector(   0 downto 0);
        signal oVar1S36: std_logic_vector(   0 downto 0);
        signal oVar1S38: std_logic_vector(   0 downto 0);
        signal oVar1S39: std_logic_vector(   0 downto 0);
        signal oVar1S40: std_logic_vector(   0 downto 0);
        signal oVar1S41: std_logic_vector(   0 downto 0);
        signal oVar1S42: std_logic_vector(   0 downto 0);
        signal oVar1S43: std_logic_vector(   0 downto 0);
        signal oVar1S44: std_logic_vector(   0 downto 0);
        signal oVar1S45: std_logic_vector(   0 downto 0);
        signal oVar1S46: std_logic_vector(   0 downto 0);
        signal oVar1S47: std_logic_vector(   0 downto 0);
        signal oVar1S48: std_logic_vector(   0 downto 0);
        signal oVar1S49: std_logic_vector(   0 downto 0);
        signal oVar1S50: std_logic_vector(   0 downto 0);
        signal oVar1S51: std_logic_vector(   0 downto 0);
        signal oVar1S52: std_logic_vector(   0 downto 0);
        signal oVar1S53: std_logic_vector(   0 downto 0);
        signal oVar1S54: std_logic_vector(   0 downto 0);
        signal oVar1S55: std_logic_vector(   0 downto 0);
        signal oVar1S56: std_logic_vector(   0 downto 0);
        signal oVar1S57: std_logic_vector(   0 downto 0);
        signal oVar1S58: std_logic_vector(   0 downto 0);
        signal oVar1S59: std_logic_vector(   0 downto 0);
        signal oVar1S60: std_logic_vector(   0 downto 0);
        signal oVar1S61: std_logic_vector(   0 downto 0);
        signal oVar1S62: std_logic_vector(   0 downto 0);
        signal oVar1S63: std_logic_vector(   0 downto 0);
        signal oVar1S64: std_logic_vector(   0 downto 0);
        signal oVar1S65: std_logic_vector(   0 downto 0);
        signal oVar1S66: std_logic_vector(   0 downto 0);
        signal oVar1S67: std_logic_vector(   0 downto 0);
        signal oVar1S68: std_logic_vector(   0 downto 0);
        signal oVar1S69: std_logic_vector(   0 downto 0);
        signal oVar1S70: std_logic_vector(   0 downto 0);
        signal oVar1S71: std_logic_vector(   0 downto 0);
        signal oVar1S72: std_logic_vector(   0 downto 0);
        signal oVar1S73: std_logic_vector(   0 downto 0);
        signal oVar1S74: std_logic_vector(   0 downto 0);
        signal oVar1S75: std_logic_vector(   0 downto 0);
        signal oVar1S76: std_logic_vector(   0 downto 0);
        signal oVar1S77: std_logic_vector(   0 downto 0);
        signal oVar1S78: std_logic_vector(   0 downto 0);
        signal oVar1S79: std_logic_vector(   0 downto 0);
        signal oVar1S80: std_logic_vector(   0 downto 0);
        signal oVar1S81: std_logic_vector(   0 downto 0);
        signal oVar1S82: std_logic_vector(   0 downto 0);
        signal oVar1S83: std_logic_vector(   0 downto 0);
        signal oVar1S84: std_logic_vector(   0 downto 0);
        signal oVar1S85: std_logic_vector(   0 downto 0);
        signal oVar1S87: std_logic_vector(   0 downto 0);
        signal oVar1S88: std_logic_vector(   0 downto 0);
        signal oVar1S89: std_logic_vector(   0 downto 0);
        signal oVar1S90: std_logic_vector(   0 downto 0);
        signal oVar1S91: std_logic_vector(   0 downto 0);
        signal oVar1S92: std_logic_vector(   0 downto 0);
        signal oVar1S93: std_logic_vector(   0 downto 0);
        signal oVar1S94: std_logic_vector(   0 downto 0);
        signal oVar1S95: std_logic_vector(   0 downto 0);
        signal oVar1S97: std_logic_vector(   0 downto 0);
        signal oVar1S98: std_logic_vector(   0 downto 0);
        signal oVar1S99: std_logic_vector(   0 downto 0);
        signal oVar1S100: std_logic_vector(   0 downto 0);
        signal oVar1S101: std_logic_vector(   0 downto 0);
        signal oVar1S102: std_logic_vector(   0 downto 0);
        signal oVar1S104: std_logic_vector(   0 downto 0);
        signal oVar1S105: std_logic_vector(   0 downto 0);
        signal oVar1S106: std_logic_vector(   0 downto 0);
        signal oVar1S107: std_logic_vector(   0 downto 0);
        signal oVar1S108: std_logic_vector(   0 downto 0);
        signal oVar1S109: std_logic_vector(   0 downto 0);
        signal oVar1S110: std_logic_vector(   0 downto 0);
        signal oVar1S111: std_logic_vector(   0 downto 0);
        signal oVar1S112: std_logic_vector(   0 downto 0);
        signal oVar1S113: std_logic_vector(   0 downto 0);
        signal oVar1S114: std_logic_vector(   0 downto 0);
        signal oVar1S115: std_logic_vector(   0 downto 0);
        signal oVar1S116: std_logic_vector(   0 downto 0);
        signal oVar1S117: std_logic_vector(   0 downto 0);
        signal oVar1S118: std_logic_vector(   0 downto 0);
        signal oVar1S119: std_logic_vector(   0 downto 0);
        signal oVar1S120: std_logic_vector(   0 downto 0);
        signal oVar1S121: std_logic_vector(   0 downto 0);
        signal oVar1S122: std_logic_vector(   0 downto 0);
        signal oVar1S123: std_logic_vector(   0 downto 0);
        signal oVar1S124: std_logic_vector(   0 downto 0);
        signal oVar1S125: std_logic_vector(   0 downto 0);
        signal oVar1S126: std_logic_vector(   0 downto 0);
        signal oVar1S127: std_logic_vector(   0 downto 0);
        signal oVar1S128: std_logic_vector(   0 downto 0);
        signal oVar1S129: std_logic_vector(   0 downto 0);
        signal oVar1S130: std_logic_vector(   0 downto 0);
        signal oVar1S131: std_logic_vector(   0 downto 0);
        signal oVar1S132: std_logic_vector(   0 downto 0);
        signal oVar1S133: std_logic_vector(   0 downto 0);
        signal oVar1S134: std_logic_vector(   0 downto 0);
        signal oVar1S135: std_logic_vector(   0 downto 0);
        signal oVar1S136: std_logic_vector(   0 downto 0);
        signal oVar1S137: std_logic_vector(   0 downto 0);
        signal oVar1S138: std_logic_vector(   0 downto 0);
        signal oVar1S139: std_logic_vector(   0 downto 0);
        signal oVar1S140: std_logic_vector(   0 downto 0);
        signal oVar1S141: std_logic_vector(   0 downto 0);
        signal oVar1S142: std_logic_vector(   0 downto 0);
        signal oVar1S143: std_logic_vector(   0 downto 0);
        signal oVar1S144: std_logic_vector(   0 downto 0);
        signal oVar1S145: std_logic_vector(   0 downto 0);
        signal oVar1S146: std_logic_vector(   0 downto 0);
        signal oVar1S147: std_logic_vector(   0 downto 0);
        signal oVar1S148: std_logic_vector(   0 downto 0);
        signal oVar1S150: std_logic_vector(   0 downto 0);
        signal oVar1S151: std_logic_vector(   0 downto 0);
        signal oVar1S152: std_logic_vector(   0 downto 0);
        signal oVar1S153: std_logic_vector(   0 downto 0);
        signal oVar1S154: std_logic_vector(   0 downto 0);
        signal oVar1S155: std_logic_vector(   0 downto 0);
        signal oVar1S156: std_logic_vector(   0 downto 0);
        signal oVar1S157: std_logic_vector(   0 downto 0);
        signal oVar1S158: std_logic_vector(   0 downto 0);
        signal oVar1S159: std_logic_vector(   0 downto 0);
        signal oVar1S160: std_logic_vector(   0 downto 0);
        signal oVar1S161: std_logic_vector(   0 downto 0);
        signal oVar1S162: std_logic_vector(   0 downto 0);
        signal oVar1S163: std_logic_vector(   0 downto 0);
        signal oVar1S164: std_logic_vector(   0 downto 0);
        signal oVar1S165: std_logic_vector(   0 downto 0);
        signal oVar1S166: std_logic_vector(   0 downto 0);
        signal oVar1S167: std_logic_vector(   0 downto 0);
        signal oVar1S168: std_logic_vector(   0 downto 0);
        signal oVar1S169: std_logic_vector(   0 downto 0);
        signal oVar1S170: std_logic_vector(   0 downto 0);
        signal oVar1S171: std_logic_vector(   0 downto 0);
        signal oVar1S172: std_logic_vector(   0 downto 0);
        signal oVar1S173: std_logic_vector(   0 downto 0);
        signal oVar1S174: std_logic_vector(   0 downto 0);
        signal oVar1S175: std_logic_vector(   0 downto 0);
        signal oVar1S176: std_logic_vector(   0 downto 0);
        signal oVar1S177: std_logic_vector(   0 downto 0);
        signal oVar1S178: std_logic_vector(   0 downto 0);
        signal oVar1S179: std_logic_vector(   0 downto 0);
        signal oVar1S180: std_logic_vector(   0 downto 0);
        signal oVar1S181: std_logic_vector(   0 downto 0);
        signal oVar1S182: std_logic_vector(   0 downto 0);
        signal oVar1S183: std_logic_vector(   0 downto 0);
        signal oVar1S184: std_logic_vector(   0 downto 0);
        signal oVar1S185: std_logic_vector(   0 downto 0);
        signal oVar1S186: std_logic_vector(   0 downto 0);
        signal oVar1S187: std_logic_vector(   0 downto 0);
        signal oVar1S188: std_logic_vector(   0 downto 0);
        signal oVar1S189: std_logic_vector(   0 downto 0);
        signal oVar1S190: std_logic_vector(   0 downto 0);
        signal oVar1S191: std_logic_vector(   0 downto 0);
        signal oVar1S192: std_logic_vector(   0 downto 0);
        signal oVar1S193: std_logic_vector(   0 downto 0);
        signal oVar1S194: std_logic_vector(   0 downto 0);
        signal oVar1S195: std_logic_vector(   0 downto 0);
        signal oVar1S196: std_logic_vector(   0 downto 0);
        signal oVar1S197: std_logic_vector(   0 downto 0);
        signal oVar1S198: std_logic_vector(   0 downto 0);
        signal oVar1S199: std_logic_vector(   0 downto 0);
        signal oVar1S200: std_logic_vector(   0 downto 0);
        signal oVar1S201: std_logic_vector(   0 downto 0);
        signal oVar1S202: std_logic_vector(   0 downto 0);
        signal oVar1S203: std_logic_vector(   0 downto 0);
        signal oVar1S204: std_logic_vector(   0 downto 0);
        signal oVar1S205: std_logic_vector(   0 downto 0);
        signal oVar1S206: std_logic_vector(   0 downto 0);
        signal oVar1S207: std_logic_vector(   0 downto 0);
        signal oVar1S208: std_logic_vector(   0 downto 0);
        signal oVar1S209: std_logic_vector(   0 downto 0);
        signal oVar1S210: std_logic_vector(   0 downto 0);
        signal oVar1S211: std_logic_vector(   0 downto 0);
        signal oVar1S212: std_logic_vector(   0 downto 0);
        signal oVar1S213: std_logic_vector(   0 downto 0);
        signal oVar1S214: std_logic_vector(   0 downto 0);
        signal oVar1S215: std_logic_vector(   0 downto 0);
        signal oVar1S216: std_logic_vector(   0 downto 0);
        signal oVar1S217: std_logic_vector(   0 downto 0);
        signal oVar1S218: std_logic_vector(   0 downto 0);
        signal oVar1S219: std_logic_vector(   0 downto 0);
        signal oVar1S220: std_logic_vector(   0 downto 0);
        signal oVar1S221: std_logic_vector(   0 downto 0);
        signal oVar1S222: std_logic_vector(   0 downto 0);
        signal oVar1S223: std_logic_vector(   0 downto 0);
        signal oVar1S224: std_logic_vector(   0 downto 0);
        signal oVar1S225: std_logic_vector(   0 downto 0);
        signal oVar1S226: std_logic_vector(   0 downto 0);
        signal oVar1S227: std_logic_vector(   0 downto 0);
        signal oVar1S228: std_logic_vector(   0 downto 0);
        signal oVar1S229: std_logic_vector(   0 downto 0);
        signal oVar1S230: std_logic_vector(   0 downto 0);
        signal oVar1S231: std_logic_vector(   0 downto 0);
        signal oVar1S232: std_logic_vector(   0 downto 0);
        signal oVar1S233: std_logic_vector(   0 downto 0);
        signal oVar1S234: std_logic_vector(   0 downto 0);
        signal oVar1S235: std_logic_vector(   0 downto 0);
        signal oVar1S236: std_logic_vector(   0 downto 0);
        signal oVar1S237: std_logic_vector(   0 downto 0);
        signal oVar1S238: std_logic_vector(   0 downto 0);
        signal oVar1S239: std_logic_vector(   0 downto 0);
        signal oVar1S240: std_logic_vector(   0 downto 0);
        signal oVar1S241: std_logic_vector(   0 downto 0);
        signal oVar1S242: std_logic_vector(   0 downto 0);
        signal oVar1S244: std_logic_vector(   0 downto 0);
        signal oVar1S245: std_logic_vector(   0 downto 0);
        signal oVar1S246: std_logic_vector(   0 downto 0);
        signal oVar1S247: std_logic_vector(   0 downto 0);
        signal oVar1S248: std_logic_vector(   0 downto 0);
        signal oVar1S249: std_logic_vector(   0 downto 0);
        signal oVar1S250: std_logic_vector(   0 downto 0);
        signal oVar1S251: std_logic_vector(   0 downto 0);
        signal oVar1S252: std_logic_vector(   0 downto 0);
        signal oVar1S253: std_logic_vector(   0 downto 0);
        signal oVar1S254: std_logic_vector(   0 downto 0);
        signal oVar1S255: std_logic_vector(   0 downto 0);
        signal oVar1S256: std_logic_vector(   0 downto 0);
        signal oVar1S257: std_logic_vector(   0 downto 0);
        signal oVar1S258: std_logic_vector(   0 downto 0);
        signal oVar1S259: std_logic_vector(   0 downto 0);
        signal oVar1S260: std_logic_vector(   0 downto 0);
        signal oVar1S261: std_logic_vector(   0 downto 0);
        signal oVar1S262: std_logic_vector(   0 downto 0);
        signal oVar1S263: std_logic_vector(   0 downto 0);
        signal oVar1S264: std_logic_vector(   0 downto 0);
        signal oVar1S265: std_logic_vector(   0 downto 0);
        signal oVar1S266: std_logic_vector(   0 downto 0);
        signal oVar1S267: std_logic_vector(   0 downto 0);
        signal oVar1S268: std_logic_vector(   0 downto 0);
        signal oVar1S269: std_logic_vector(   0 downto 0);
        signal oVar1S270: std_logic_vector(   0 downto 0);
        signal oVar1S271: std_logic_vector(   0 downto 0);
        signal oVar1S272: std_logic_vector(   0 downto 0);
        signal oVar1S273: std_logic_vector(   0 downto 0);
        signal oVar1S274: std_logic_vector(   0 downto 0);
        signal oVar1S275: std_logic_vector(   0 downto 0);
        signal oVar1S276: std_logic_vector(   0 downto 0);
        signal oVar1S277: std_logic_vector(   0 downto 0);
        signal oVar1S279: std_logic_vector(   0 downto 0);
        signal oVar1S280: std_logic_vector(   0 downto 0);
        signal oVar1S281: std_logic_vector(   0 downto 0);
        signal oVar1S282: std_logic_vector(   0 downto 0);
        signal oVar1S283: std_logic_vector(   0 downto 0);
        signal oVar1S284: std_logic_vector(   0 downto 0);
        signal oVar1S285: std_logic_vector(   0 downto 0);
        signal oVar1S286: std_logic_vector(   0 downto 0);
        signal oVar1S287: std_logic_vector(   0 downto 0);
        signal oVar1S288: std_logic_vector(   0 downto 0);
        signal oVar1S289: std_logic_vector(   0 downto 0);
        signal oVar1S290: std_logic_vector(   0 downto 0);
        signal oVar1S291: std_logic_vector(   0 downto 0);
        signal oVar1S292: std_logic_vector(   0 downto 0);
        signal oVar1S293: std_logic_vector(   0 downto 0);
        signal oVar1S294: std_logic_vector(   0 downto 0);
        signal oVar1S295: std_logic_vector(   0 downto 0);
        signal oVar1S297: std_logic_vector(   0 downto 0);
        signal oVar1S298: std_logic_vector(   0 downto 0);
        signal oVar1S299: std_logic_vector(   0 downto 0);
        signal oVar1S300: std_logic_vector(   0 downto 0);
        signal oVar1S301: std_logic_vector(   0 downto 0);
        signal oVar1S302: std_logic_vector(   0 downto 0);
        signal oVar1S303: std_logic_vector(   0 downto 0);
        signal oVar1S304: std_logic_vector(   0 downto 0);
        signal oVar1S305: std_logic_vector(   0 downto 0);
        signal oVar1S306: std_logic_vector(   0 downto 0);
        signal oVar1S307: std_logic_vector(   0 downto 0);
        signal oVar1S308: std_logic_vector(   0 downto 0);
        signal oVar1S309: std_logic_vector(   0 downto 0);
        signal oVar1S310: std_logic_vector(   0 downto 0);
        signal oVar1S311: std_logic_vector(   0 downto 0);
        signal oVar1S312: std_logic_vector(   0 downto 0);
        signal oVar1S313: std_logic_vector(   0 downto 0);
        signal oVar1S314: std_logic_vector(   0 downto 0);
        signal oVar1S315: std_logic_vector(   0 downto 0);
        signal oVar1S317: std_logic_vector(   0 downto 0);
        signal oVar1S318: std_logic_vector(   0 downto 0);
        signal oVar1S319: std_logic_vector(   0 downto 0);
        signal oVar1S320: std_logic_vector(   0 downto 0);
        signal oVar1S321: std_logic_vector(   0 downto 0);
        signal oVar1S322: std_logic_vector(   0 downto 0);
        signal oVar1S323: std_logic_vector(   0 downto 0);
        signal oVar1S324: std_logic_vector(   0 downto 0);
        signal oVar1S325: std_logic_vector(   0 downto 0);
        signal oVar1S326: std_logic_vector(   0 downto 0);
        signal oVar1S327: std_logic_vector(   0 downto 0);
        signal oVar1S328: std_logic_vector(   0 downto 0);
        signal oVar1S329: std_logic_vector(   0 downto 0);
        signal oVar1S330: std_logic_vector(   0 downto 0);
        signal oVar1S331: std_logic_vector(   0 downto 0);
        signal oVar1S332: std_logic_vector(   0 downto 0);
        signal oVar1S333: std_logic_vector(   0 downto 0);
        signal oVar1S334: std_logic_vector(   0 downto 0);
        signal oVar1S335: std_logic_vector(   0 downto 0);
        signal oVar1S336: std_logic_vector(   0 downto 0);
        signal oVar1S337: std_logic_vector(   0 downto 0);
        signal oVar1S338: std_logic_vector(   0 downto 0);
        signal oVar1S339: std_logic_vector(   0 downto 0);
        signal oVar1S340: std_logic_vector(   0 downto 0);
        signal oVar1S341: std_logic_vector(   0 downto 0);
        signal oVar1S342: std_logic_vector(   0 downto 0);
        signal oVar1S343: std_logic_vector(   0 downto 0);
        signal oVar1S344: std_logic_vector(   0 downto 0);
        signal oVar1S345: std_logic_vector(   0 downto 0);
        signal oVar1S346: std_logic_vector(   0 downto 0);
        signal oVar1S347: std_logic_vector(   0 downto 0);
        signal oVar1S348: std_logic_vector(   0 downto 0);
        signal oVar1S349: std_logic_vector(   0 downto 0);
        signal oVar1S350: std_logic_vector(   0 downto 0);
        signal oVar1S351: std_logic_vector(   0 downto 0);
        signal oVar1S352: std_logic_vector(   0 downto 0);
        signal oVar1S353: std_logic_vector(   0 downto 0);
        signal oVar1S354: std_logic_vector(   0 downto 0);
        signal oVar1S355: std_logic_vector(   0 downto 0);
        signal oVar1S356: std_logic_vector(   0 downto 0);
        signal oVar1S357: std_logic_vector(   0 downto 0);
        signal oVar1S358: std_logic_vector(   0 downto 0);
        signal oVar1S359: std_logic_vector(   0 downto 0);
        signal oVar1S360: std_logic_vector(   0 downto 0);
        signal oVar1S361: std_logic_vector(   0 downto 0);
        signal oVar1S362: std_logic_vector(   0 downto 0);
        signal oVar1S363: std_logic_vector(   0 downto 0);
        signal oVar1S364: std_logic_vector(   0 downto 0);
        signal oVar1S365: std_logic_vector(   0 downto 0);
        signal oVar1S366: std_logic_vector(   0 downto 0);
        signal oVar1S367: std_logic_vector(   0 downto 0);
        signal oVar1S368: std_logic_vector(   0 downto 0);
        signal oVar1S369: std_logic_vector(   0 downto 0);
        signal oVar1S370: std_logic_vector(   0 downto 0);
        signal oVar1S371: std_logic_vector(   0 downto 0);
        signal oVar1S372: std_logic_vector(   0 downto 0);
        signal oVar1S373: std_logic_vector(   0 downto 0);
        signal oVar1S374: std_logic_vector(   0 downto 0);
        signal oVar1S375: std_logic_vector(   0 downto 0);
        signal oVar1S376: std_logic_vector(   0 downto 0);
        signal oVar1S377: std_logic_vector(   0 downto 0);
        signal oVar1S378: std_logic_vector(   0 downto 0);
        signal oVar1S379: std_logic_vector(   0 downto 0);
        signal oVar1S380: std_logic_vector(   0 downto 0);
        signal oVar1S381: std_logic_vector(   0 downto 0);
        signal oVar1S382: std_logic_vector(   0 downto 0);
        signal oVar1S383: std_logic_vector(   0 downto 0);
        signal oVar1S384: std_logic_vector(   0 downto 0);
        signal oVar1S385: std_logic_vector(   0 downto 0);
        signal oVar1S386: std_logic_vector(   0 downto 0);
        signal oVar1S387: std_logic_vector(   0 downto 0);
        signal oVar1S388: std_logic_vector(   0 downto 0);
        signal oVar1S389: std_logic_vector(   0 downto 0);
        signal oVar1S390: std_logic_vector(   0 downto 0);
        signal oVar1S391: std_logic_vector(   0 downto 0);
        signal oVar1S392: std_logic_vector(   0 downto 0);
        signal oVar1S393: std_logic_vector(   0 downto 0);
        signal oVar1S394: std_logic_vector(   0 downto 0);
        signal oVar1S395: std_logic_vector(   0 downto 0);
        signal oVar1S396: std_logic_vector(   0 downto 0);
        signal oVar1S397: std_logic_vector(   0 downto 0);
        signal oVar1S398: std_logic_vector(   0 downto 0);
        signal oVar1S399: std_logic_vector(   0 downto 0);
        signal oVar1S400: std_logic_vector(   0 downto 0);
        signal oVar1S401: std_logic_vector(   0 downto 0);
        signal oVar1S402: std_logic_vector(   0 downto 0);
        signal oVar1S403: std_logic_vector(   0 downto 0);
        signal oVar1S404: std_logic_vector(   0 downto 0);
        signal oVar1S405: std_logic_vector(   0 downto 0);
        signal oVar1S406: std_logic_vector(   0 downto 0);
        signal oVar1S407: std_logic_vector(   0 downto 0);
        signal oVar1S408: std_logic_vector(   0 downto 0);
        signal oVar1S409: std_logic_vector(   0 downto 0);
        signal oVar1S410: std_logic_vector(   0 downto 0);
        signal oVar1S411: std_logic_vector(   0 downto 0);
        signal oVar1S412: std_logic_vector(   0 downto 0);
        signal oVar1S413: std_logic_vector(   0 downto 0);
        signal oVar1S414: std_logic_vector(   0 downto 0);
        signal oVar1S415: std_logic_vector(   0 downto 0);
        signal oVar1S416: std_logic_vector(   0 downto 0);
        signal oVar1S417: std_logic_vector(   0 downto 0);
        signal oVar1S418: std_logic_vector(   0 downto 0);
        signal oVar1S419: std_logic_vector(   0 downto 0);
        signal oVar1S420: std_logic_vector(   0 downto 0);
        signal oVar1S421: std_logic_vector(   0 downto 0);
        signal oVar1S422: std_logic_vector(   0 downto 0);
        signal oVar1S423: std_logic_vector(   0 downto 0);
        signal oVar1S424: std_logic_vector(   0 downto 0);
        signal oVar1S425: std_logic_vector(   0 downto 0);
        signal oVar1S426: std_logic_vector(   0 downto 0);
        signal oVar1S427: std_logic_vector(   0 downto 0);
        signal oVar1S428: std_logic_vector(   0 downto 0);
        signal oVar1S429: std_logic_vector(   0 downto 0);
        signal oVar1S430: std_logic_vector(   0 downto 0);
        signal oVar1S431: std_logic_vector(   0 downto 0);
        signal oVar1S432: std_logic_vector(   0 downto 0);
        signal oVar1S434: std_logic_vector(   0 downto 0);
        signal oVar1S435: std_logic_vector(   0 downto 0);
        signal oVar1S436: std_logic_vector(   0 downto 0);
        signal oVar1S437: std_logic_vector(   0 downto 0);
        signal oVar1S438: std_logic_vector(   0 downto 0);
        signal oVar1S439: std_logic_vector(   0 downto 0);
        signal oVar1S440: std_logic_vector(   0 downto 0);
        signal oVar1S441: std_logic_vector(   0 downto 0);
        signal oVar1S442: std_logic_vector(   0 downto 0);
        signal oVar1S443: std_logic_vector(   0 downto 0);
        signal oVar1S444: std_logic_vector(   0 downto 0);
        signal oVar1S445: std_logic_vector(   0 downto 0);
        signal oVar1S446: std_logic_vector(   0 downto 0);
        signal oVar1S447: std_logic_vector(   0 downto 0);
        signal oVar1S448: std_logic_vector(   0 downto 0);
        signal oVar1S449: std_logic_vector(   0 downto 0);
        signal oVar1S450: std_logic_vector(   0 downto 0);
        signal oVar1S451: std_logic_vector(   0 downto 0);
        signal oVar1S452: std_logic_vector(   0 downto 0);
        signal oVar1S453: std_logic_vector(   0 downto 0);
        signal oVar1S454: std_logic_vector(   0 downto 0);
        signal oVar1S455: std_logic_vector(   0 downto 0);
        signal oVar1S456: std_logic_vector(   0 downto 0);
        signal oVar1S457: std_logic_vector(   0 downto 0);
        signal oVar1S458: std_logic_vector(   0 downto 0);
        signal oVar1S460: std_logic_vector(   0 downto 0);
        signal oVar1S461: std_logic_vector(   0 downto 0);
        signal oVar1S462: std_logic_vector(   0 downto 0);
        signal oVar1S463: std_logic_vector(   0 downto 0);
        signal oVar1S464: std_logic_vector(   0 downto 0);
        signal oVar1S465: std_logic_vector(   0 downto 0);
        signal oVar1S466: std_logic_vector(   0 downto 0);
        signal oVar1S468: std_logic_vector(   0 downto 0);
        signal oVar1S469: std_logic_vector(   0 downto 0);
        signal oVar1S470: std_logic_vector(   0 downto 0);
        signal oVar1S471: std_logic_vector(   0 downto 0);
        signal oVar1S472: std_logic_vector(   0 downto 0);
        signal oVar1S473: std_logic_vector(   0 downto 0);
        signal oVar1S474: std_logic_vector(   0 downto 0);
        signal oVar1S475: std_logic_vector(   0 downto 0);
        signal oVar1S476: std_logic_vector(   0 downto 0);
        signal oVar1S477: std_logic_vector(   0 downto 0);
        signal oVar1S478: std_logic_vector(   0 downto 0);
        signal oVar1S479: std_logic_vector(   0 downto 0);
        signal oVar1S480: std_logic_vector(   0 downto 0);
        signal oVar1S481: std_logic_vector(   0 downto 0);
        signal oVar1S482: std_logic_vector(   0 downto 0);
        signal oVar1S483: std_logic_vector(   0 downto 0);
        signal oVar1S484: std_logic_vector(   0 downto 0);
        signal oVar1S485: std_logic_vector(   0 downto 0);
        signal oVar1S486: std_logic_vector(   0 downto 0);
        signal oVar1S488: std_logic_vector(   0 downto 0);
        signal oVar1S489: std_logic_vector(   0 downto 0);
        signal oVar1S490: std_logic_vector(   0 downto 0);
        signal oVar1S491: std_logic_vector(   0 downto 0);
        signal oVar1S492: std_logic_vector(   0 downto 0);
        signal oVar1S493: std_logic_vector(   0 downto 0);
        signal oVar1S494: std_logic_vector(   0 downto 0);
        signal oVar1S495: std_logic_vector(   0 downto 0);
        signal oVar1S497: std_logic_vector(   0 downto 0);
        signal oVar1S498: std_logic_vector(   0 downto 0);
        signal oVar1S499: std_logic_vector(   0 downto 0);
        signal oVar1S500: std_logic_vector(   0 downto 0);
        signal oVar1S501: std_logic_vector(   0 downto 0);
        signal oVar1S502: std_logic_vector(   0 downto 0);
        signal oVar1S503: std_logic_vector(   0 downto 0);
        signal oVar1S504: std_logic_vector(   0 downto 0);
        signal oVar1S505: std_logic_vector(   0 downto 0);
        signal oVar1S506: std_logic_vector(   0 downto 0);
        signal oVar1S507: std_logic_vector(   0 downto 0);
        signal oVar1S508: std_logic_vector(   0 downto 0);
        signal oVar1S509: std_logic_vector(   0 downto 0);
        signal oVar1S510: std_logic_vector(   0 downto 0);
        signal oVar1S511: std_logic_vector(   0 downto 0);
        signal oVar1S512: std_logic_vector(   0 downto 0);
        signal oVar1S513: std_logic_vector(   0 downto 0);
        signal oVar1S514: std_logic_vector(   0 downto 0);
        signal oVar1S515: std_logic_vector(   0 downto 0);
        signal oVar1S516: std_logic_vector(   0 downto 0);
        signal oVar1S517: std_logic_vector(   0 downto 0);
        signal oVar1S518: std_logic_vector(   0 downto 0);
        signal oVar1S519: std_logic_vector(   0 downto 0);
        signal oVar1S520: std_logic_vector(   0 downto 0);
        signal oVar1S521: std_logic_vector(   0 downto 0);
        signal oVar1S522: std_logic_vector(   0 downto 0);
        signal oVar1S523: std_logic_vector(   0 downto 0);
        signal oVar1S524: std_logic_vector(   0 downto 0);
        signal oVar1S525: std_logic_vector(   0 downto 0);
        signal oVar1S526: std_logic_vector(   0 downto 0);
        signal oVar1S527: std_logic_vector(   0 downto 0);
        signal oVar1S528: std_logic_vector(   0 downto 0);
        signal oVar1S529: std_logic_vector(   0 downto 0);
        signal oVar1S530: std_logic_vector(   0 downto 0);
        signal oVar1S531: std_logic_vector(   0 downto 0);
        signal oVar1S532: std_logic_vector(   0 downto 0);
        signal oVar1S533: std_logic_vector(   0 downto 0);
        signal oVar1S534: std_logic_vector(   0 downto 0);
        signal oVar1S535: std_logic_vector(   0 downto 0);
        signal oVar1S536: std_logic_vector(   0 downto 0);
        signal oVar1S537: std_logic_vector(   0 downto 0);
        signal oVar1S538: std_logic_vector(   0 downto 0);
        signal oVar1S539: std_logic_vector(   0 downto 0);
        signal oVar1S540: std_logic_vector(   0 downto 0);
        signal oVar1S541: std_logic_vector(   0 downto 0);
        signal oVar1S542: std_logic_vector(   0 downto 0);
        signal oVar1S543: std_logic_vector(   0 downto 0);
        signal oVar1S544: std_logic_vector(   0 downto 0);
        signal oVar1S545: std_logic_vector(   0 downto 0);
        signal oVar1S546: std_logic_vector(   0 downto 0);
        signal oVar1S547: std_logic_vector(   0 downto 0);
        signal oVar1S548: std_logic_vector(   0 downto 0);
        signal oVar1S549: std_logic_vector(   0 downto 0);
        signal oVar1S550: std_logic_vector(   0 downto 0);
        signal oVar1S551: std_logic_vector(   0 downto 0);
        signal oVar1S552: std_logic_vector(   0 downto 0);
        signal oVar1S553: std_logic_vector(   0 downto 0);
        signal oVar1S554: std_logic_vector(   0 downto 0);
        signal oVar1S555: std_logic_vector(   0 downto 0);
        signal oVar1S556: std_logic_vector(   0 downto 0);
        signal oVar1S557: std_logic_vector(   0 downto 0);
        signal oVar1S558: std_logic_vector(   0 downto 0);
        signal oVar1S559: std_logic_vector(   0 downto 0);
        signal oVar1S560: std_logic_vector(   0 downto 0);
        signal oVar1S561: std_logic_vector(   0 downto 0);
        signal oVar1S562: std_logic_vector(   0 downto 0);
        signal oVar1S563: std_logic_vector(   0 downto 0);
        signal oVar1S564: std_logic_vector(   0 downto 0);
        signal oVar1S565: std_logic_vector(   0 downto 0);
        signal oVar1S566: std_logic_vector(   0 downto 0);
        signal oVar1S568: std_logic_vector(   0 downto 0);
        signal oVar1S569: std_logic_vector(   0 downto 0);
        signal oVar1S570: std_logic_vector(   0 downto 0);
        signal oVar1S571: std_logic_vector(   0 downto 0);
        signal oVar1S572: std_logic_vector(   0 downto 0);
        signal oVar1S573: std_logic_vector(   0 downto 0);
        signal oVar1S574: std_logic_vector(   0 downto 0);
        signal oVar1S575: std_logic_vector(   0 downto 0);
        signal oVar1S576: std_logic_vector(   0 downto 0);
        signal oVar1S577: std_logic_vector(   0 downto 0);
        signal oVar1S578: std_logic_vector(   0 downto 0);
        signal oVar1S579: std_logic_vector(   0 downto 0);
        signal oVar1S580: std_logic_vector(   0 downto 0);
        signal oVar1S582: std_logic_vector(   0 downto 0);
        signal oVar1S583: std_logic_vector(   0 downto 0);
        signal oVar1S584: std_logic_vector(   0 downto 0);
        signal oVar1S585: std_logic_vector(   0 downto 0);
        signal oVar1S586: std_logic_vector(   0 downto 0);
        signal oVar1S587: std_logic_vector(   0 downto 0);
        signal oVar1S588: std_logic_vector(   0 downto 0);
        signal oVar1S589: std_logic_vector(   0 downto 0);
        signal oVar1S590: std_logic_vector(   0 downto 0);
        signal oVar1S591: std_logic_vector(   0 downto 0);
        signal oVar1S592: std_logic_vector(   0 downto 0);
        signal oVar1S593: std_logic_vector(   0 downto 0);
        signal oVar1S594: std_logic_vector(   0 downto 0);
        signal oVar1S595: std_logic_vector(   0 downto 0);
        signal oVar1S596: std_logic_vector(   0 downto 0);
        signal oVar1S597: std_logic_vector(   0 downto 0);
        signal oVar1S598: std_logic_vector(   0 downto 0);
        signal oVar1S600: std_logic_vector(   0 downto 0);
        signal oVar1S601: std_logic_vector(   0 downto 0);
        signal oVar1S602: std_logic_vector(   0 downto 0);
        signal oVar1S603: std_logic_vector(   0 downto 0);
        signal oVar1S604: std_logic_vector(   0 downto 0);
        signal oVar1S605: std_logic_vector(   0 downto 0);
        signal oVar1S606: std_logic_vector(   0 downto 0);
        signal oVar1S607: std_logic_vector(   0 downto 0);
        signal oVar1S608: std_logic_vector(   0 downto 0);
        signal oVar1S609: std_logic_vector(   0 downto 0);
        signal oVar1S610: std_logic_vector(   0 downto 0);
        signal oVar1S611: std_logic_vector(   0 downto 0);
        signal oVar1S612: std_logic_vector(   0 downto 0);
        signal oVar1S613: std_logic_vector(   0 downto 0);
        signal oVar1S614: std_logic_vector(   0 downto 0);
        signal oVar1S615: std_logic_vector(   0 downto 0);
        signal oVar1S616: std_logic_vector(   0 downto 0);
        signal oVar1S617: std_logic_vector(   0 downto 0);
        signal oVar1S618: std_logic_vector(   0 downto 0);
        signal oVar1S619: std_logic_vector(   0 downto 0);
        signal oVar1S621: std_logic_vector(   0 downto 0);
        signal oVar1S622: std_logic_vector(   0 downto 0);
        signal oVar1S623: std_logic_vector(   0 downto 0);
        signal oVar1S624: std_logic_vector(   0 downto 0);
        signal oVar1S625: std_logic_vector(   0 downto 0);
        signal oVar1S626: std_logic_vector(   0 downto 0);
        signal oVar1S627: std_logic_vector(   0 downto 0);
        signal oVar1S629: std_logic_vector(   0 downto 0);
        signal oVar1S630: std_logic_vector(   0 downto 0);
        signal oVar1S631: std_logic_vector(   0 downto 0);
        signal oVar1S632: std_logic_vector(   0 downto 0);
        signal oVar1S633: std_logic_vector(   0 downto 0);
        signal oVar1S634: std_logic_vector(   0 downto 0);
        signal oVar1S635: std_logic_vector(   0 downto 0);
        signal oVar1S636: std_logic_vector(   0 downto 0);
        signal oVar1S637: std_logic_vector(   0 downto 0);
        signal oVar1S638: std_logic_vector(   0 downto 0);
        signal oVar1S639: std_logic_vector(   0 downto 0);
        signal oVar1S640: std_logic_vector(   0 downto 0);
        signal oVar1S641: std_logic_vector(   0 downto 0);
        signal oVar1S642: std_logic_vector(   0 downto 0);
        signal oVar1S643: std_logic_vector(   0 downto 0);
        signal oVar1S644: std_logic_vector(   0 downto 0);
        signal oVar1S646: std_logic_vector(   0 downto 0);
        signal oVar1S647: std_logic_vector(   0 downto 0);
        signal oVar1S648: std_logic_vector(   0 downto 0);
        signal oVar1S649: std_logic_vector(   0 downto 0);
        signal oVar1S650: std_logic_vector(   0 downto 0);
        signal oVar1S651: std_logic_vector(   0 downto 0);
        signal oVar1S652: std_logic_vector(   0 downto 0);
        signal oVar1S653: std_logic_vector(   0 downto 0);
        signal oVar1S654: std_logic_vector(   0 downto 0);
        signal oVar1S655: std_logic_vector(   0 downto 0);
        signal oVar1S656: std_logic_vector(   0 downto 0);
        signal oVar1S657: std_logic_vector(   0 downto 0);
        signal oVar1S658: std_logic_vector(   0 downto 0);
        signal oVar1S659: std_logic_vector(   0 downto 0);
        signal oVar1S660: std_logic_vector(   0 downto 0);
        signal oVar1S662: std_logic_vector(   0 downto 0);
        signal oVar1S663: std_logic_vector(   0 downto 0);
        signal oVar1S664: std_logic_vector(   0 downto 0);
        signal oVar1S665: std_logic_vector(   0 downto 0);
        signal oVar1S666: std_logic_vector(   0 downto 0);
        signal oVar1S667: std_logic_vector(   0 downto 0);
        signal oVar1S668: std_logic_vector(   0 downto 0);
        signal oVar1S669: std_logic_vector(   0 downto 0);
        signal oVar1S670: std_logic_vector(   0 downto 0);
        signal oVar1S671: std_logic_vector(   0 downto 0);
        signal oVar1S672: std_logic_vector(   0 downto 0);
        signal oVar1S673: std_logic_vector(   0 downto 0);
        signal oVar1S674: std_logic_vector(   0 downto 0);
        signal oVar1S675: std_logic_vector(   0 downto 0);
        signal oVar1S676: std_logic_vector(   0 downto 0);
        signal oVar1S677: std_logic_vector(   0 downto 0);
        signal oVar1S678: std_logic_vector(   0 downto 0);
        signal oVar1S679: std_logic_vector(   0 downto 0);
        signal oVar1S680: std_logic_vector(   0 downto 0);
        signal oVar1S681: std_logic_vector(   0 downto 0);
        signal oVar1S682: std_logic_vector(   0 downto 0);
        signal oVar1S683: std_logic_vector(   0 downto 0);
        signal oVar1S684: std_logic_vector(   0 downto 0);
        signal oVar1S685: std_logic_vector(   0 downto 0);
        signal oVar1S686: std_logic_vector(   0 downto 0);
        signal oVar1S687: std_logic_vector(   0 downto 0);
        signal oVar1S688: std_logic_vector(   0 downto 0);
        signal oVar1S689: std_logic_vector(   0 downto 0);
        signal oVar1S690: std_logic_vector(   0 downto 0);
        signal oVar1S691: std_logic_vector(   0 downto 0);
        signal oVar1S692: std_logic_vector(   0 downto 0);
        signal oVar1S693: std_logic_vector(   0 downto 0);
        signal oVar1S694: std_logic_vector(   0 downto 0);
        signal oVar1S695: std_logic_vector(   0 downto 0);
        signal oVar1S696: std_logic_vector(   0 downto 0);
        signal oVar1S697: std_logic_vector(   0 downto 0);
        signal oVar1S698: std_logic_vector(   0 downto 0);
        signal oVar1S699: std_logic_vector(   0 downto 0);
        signal oVar1S700: std_logic_vector(   0 downto 0);
        signal oVar1S701: std_logic_vector(   0 downto 0);
        signal oVar1S702: std_logic_vector(   0 downto 0);
        signal oVar1S703: std_logic_vector(   0 downto 0);
        signal oVar1S704: std_logic_vector(   0 downto 0);
        signal oVar1S705: std_logic_vector(   0 downto 0);
        signal oVar1S706: std_logic_vector(   0 downto 0);
        signal oVar1S707: std_logic_vector(   0 downto 0);
        signal oVar1S708: std_logic_vector(   0 downto 0);
        signal oVar1S709: std_logic_vector(   0 downto 0);
        signal oVar1S710: std_logic_vector(   0 downto 0);
        signal oVar1S711: std_logic_vector(   0 downto 0);
        signal oVar1S712: std_logic_vector(   0 downto 0);
        signal oVar1S713: std_logic_vector(   0 downto 0);
        signal oVar1S714: std_logic_vector(   0 downto 0);
        signal oVar1S715: std_logic_vector(   0 downto 0);
        signal oVar1S716: std_logic_vector(   0 downto 0);
        signal oVar1S717: std_logic_vector(   0 downto 0);
        signal oVar1S718: std_logic_vector(   0 downto 0);
        signal oVar1S719: std_logic_vector(   0 downto 0);
        signal oVar1S720: std_logic_vector(   0 downto 0);
        signal oVar1S721: std_logic_vector(   0 downto 0);
        signal oVar1S722: std_logic_vector(   0 downto 0);
        signal oVar1S723: std_logic_vector(   0 downto 0);
        signal oVar1S724: std_logic_vector(   0 downto 0);
        signal oVar1S725: std_logic_vector(   0 downto 0);
        signal oVar1S726: std_logic_vector(   0 downto 0);
        signal oVar1S727: std_logic_vector(   0 downto 0);
        signal oVar1S728: std_logic_vector(   0 downto 0);
        signal oVar1S729: std_logic_vector(   0 downto 0);
        signal oVar1S730: std_logic_vector(   0 downto 0);
        signal oVar1S731: std_logic_vector(   0 downto 0);
        signal oVar1S732: std_logic_vector(   0 downto 0);
        signal oVar1S733: std_logic_vector(   0 downto 0);
        signal oVar1S734: std_logic_vector(   0 downto 0);
        signal oVar1S735: std_logic_vector(   0 downto 0);
        signal oVar1S736: std_logic_vector(   0 downto 0);
        signal oVar1S737: std_logic_vector(   0 downto 0);
        signal oVar1S739: std_logic_vector(   0 downto 0);
        signal oVar1S740: std_logic_vector(   0 downto 0);
        signal oVar1S741: std_logic_vector(   0 downto 0);
        signal oVar1S742: std_logic_vector(   0 downto 0);
        signal oVar1S743: std_logic_vector(   0 downto 0);
        signal oVar1S744: std_logic_vector(   0 downto 0);
        signal oVar1S745: std_logic_vector(   0 downto 0);
        signal oVar1S746: std_logic_vector(   0 downto 0);
        signal oVar1S747: std_logic_vector(   0 downto 0);
        signal oVar1S748: std_logic_vector(   0 downto 0);
        signal oVar1S749: std_logic_vector(   0 downto 0);
        signal oVar1S750: std_logic_vector(   0 downto 0);
        signal oVar1S751: std_logic_vector(   0 downto 0);
        signal oVar1S752: std_logic_vector(   0 downto 0);
        signal oVar1S753: std_logic_vector(   0 downto 0);
        signal oVar1S754: std_logic_vector(   0 downto 0);
        signal oVar1S755: std_logic_vector(   0 downto 0);
        signal oVar1S756: std_logic_vector(   0 downto 0);
        signal oVar1S757: std_logic_vector(   0 downto 0);
        signal oVar1S758: std_logic_vector(   0 downto 0);
        signal oVar1S759: std_logic_vector(   0 downto 0);
        signal oVar1S760: std_logic_vector(   0 downto 0);
        signal oVar1S761: std_logic_vector(   0 downto 0);
        signal oVar1S762: std_logic_vector(   0 downto 0);
        signal oVar1S763: std_logic_vector(   0 downto 0);
        signal oVar1S764: std_logic_vector(   0 downto 0);
        signal oVar1S765: std_logic_vector(   0 downto 0);
        signal oVar1S766: std_logic_vector(   0 downto 0);
        signal oVar1S767: std_logic_vector(   0 downto 0);
        signal oVar1S768: std_logic_vector(   0 downto 0);
        signal oVar1S769: std_logic_vector(   0 downto 0);
        signal oVar1S770: std_logic_vector(   0 downto 0);
        signal oVar1S771: std_logic_vector(   0 downto 0);
        signal oVar1S772: std_logic_vector(   0 downto 0);
        signal oVar1S773: std_logic_vector(   0 downto 0);
        signal oVar1S774: std_logic_vector(   0 downto 0);
        signal oVar1S775: std_logic_vector(   0 downto 0);
        signal oVar1S776: std_logic_vector(   0 downto 0);
        signal oVar1S777: std_logic_vector(   0 downto 0);
        signal oVar1S778: std_logic_vector(   0 downto 0);
        signal oVar1S779: std_logic_vector(   0 downto 0);
        signal oVar1S780: std_logic_vector(   0 downto 0);
        signal oVar1S782: std_logic_vector(   0 downto 0);
        signal oVar1S783: std_logic_vector(   0 downto 0);
        signal oVar1S784: std_logic_vector(   0 downto 0);
        signal oVar1S785: std_logic_vector(   0 downto 0);
        signal oVar1S786: std_logic_vector(   0 downto 0);
        signal oVar1S787: std_logic_vector(   0 downto 0);
        signal oVar1S788: std_logic_vector(   0 downto 0);
        signal oVar1S789: std_logic_vector(   0 downto 0);
        signal oVar1S790: std_logic_vector(   0 downto 0);
        signal oVar1S791: std_logic_vector(   0 downto 0);
        signal oVar1S792: std_logic_vector(   0 downto 0);
        signal oVar1S793: std_logic_vector(   0 downto 0);
        signal oVar1S794: std_logic_vector(   0 downto 0);
        signal oVar1S795: std_logic_vector(   0 downto 0);
        signal oVar1S796: std_logic_vector(   0 downto 0);
        signal oVar1S797: std_logic_vector(   0 downto 0);
        signal oVar1S798: std_logic_vector(   0 downto 0);
        signal oVar1S799: std_logic_vector(   0 downto 0);
        signal oVar1S800: std_logic_vector(   0 downto 0);
        signal oVar1S801: std_logic_vector(   0 downto 0);
        signal oVar1S802: std_logic_vector(   0 downto 0);
        signal oVar1S803: std_logic_vector(   0 downto 0);
        signal oVar1S804: std_logic_vector(   0 downto 0);
        signal oVar1S805: std_logic_vector(   0 downto 0);
        signal oVar1S806: std_logic_vector(   0 downto 0);
        signal oVar1S807: std_logic_vector(   0 downto 0);
        signal oVar1S808: std_logic_vector(   0 downto 0);
        signal oVar1S809: std_logic_vector(   0 downto 0);
        signal oVar1S810: std_logic_vector(   0 downto 0);
        signal oVar1S811: std_logic_vector(   0 downto 0);
        signal oVar1S812: std_logic_vector(   0 downto 0);
        signal oVar1S813: std_logic_vector(   0 downto 0);
        signal oVar1S814: std_logic_vector(   0 downto 0);
        signal oVar1S815: std_logic_vector(   0 downto 0);
        signal oVar1S816: std_logic_vector(   0 downto 0);
        signal oVar1S817: std_logic_vector(   0 downto 0);
        signal oVar1S818: std_logic_vector(   0 downto 0);
        signal oVar1S819: std_logic_vector(   0 downto 0);
        signal oVar1S820: std_logic_vector(   0 downto 0);
        signal oVar1S821: std_logic_vector(   0 downto 0);
        signal oVar1S822: std_logic_vector(   0 downto 0);
        signal oVar1S823: std_logic_vector(   0 downto 0);
        signal oVar1S824: std_logic_vector(   0 downto 0);
        signal oVar1S826: std_logic_vector(   0 downto 0);
        signal oVar1S827: std_logic_vector(   0 downto 0);
        signal oVar1S828: std_logic_vector(   0 downto 0);
        signal oVar1S829: std_logic_vector(   0 downto 0);
        signal oVar1S830: std_logic_vector(   0 downto 0);
        signal oVar1S831: std_logic_vector(   0 downto 0);
        signal oVar1S832: std_logic_vector(   0 downto 0);
        signal oVar1S833: std_logic_vector(   0 downto 0);
        signal oVar1S834: std_logic_vector(   0 downto 0);
        signal oVar1S836: std_logic_vector(   0 downto 0);
        signal oVar1S837: std_logic_vector(   0 downto 0);
        signal oVar1S838: std_logic_vector(   0 downto 0);
        signal oVar1S839: std_logic_vector(   0 downto 0);
        signal oVar1S840: std_logic_vector(   0 downto 0);
        signal oVar1S841: std_logic_vector(   0 downto 0);
        signal oVar1S842: std_logic_vector(   0 downto 0);
        signal oVar1S843: std_logic_vector(   0 downto 0);
        signal oVar1S844: std_logic_vector(   0 downto 0);
        signal oVar1S845: std_logic_vector(   0 downto 0);
        signal oVar1S846: std_logic_vector(   0 downto 0);
        signal oVar1S847: std_logic_vector(   0 downto 0);
        signal oVar1S848: std_logic_vector(   0 downto 0);
        signal oVar1S849: std_logic_vector(   0 downto 0);
        signal oVar1S850: std_logic_vector(   0 downto 0);
        signal oVar1S851: std_logic_vector(   0 downto 0);
        signal oVar1S852: std_logic_vector(   0 downto 0);
        signal oVar1S853: std_logic_vector(   0 downto 0);
        signal oVar1S854: std_logic_vector(   0 downto 0);
        signal oVar1S855: std_logic_vector(   0 downto 0);
        signal oVar1S856: std_logic_vector(   0 downto 0);
        signal oVar1S857: std_logic_vector(   0 downto 0);
        signal oVar1S858: std_logic_vector(   0 downto 0);
        signal oVar1S859: std_logic_vector(   0 downto 0);
        signal oVar1S860: std_logic_vector(   0 downto 0);
        signal oVar1S861: std_logic_vector(   0 downto 0);
        signal oVar1S862: std_logic_vector(   0 downto 0);
        signal oVar1S863: std_logic_vector(   0 downto 0);
        signal oVar1S864: std_logic_vector(   0 downto 0);
        signal oVar1S865: std_logic_vector(   0 downto 0);
        signal oVar1S866: std_logic_vector(   0 downto 0);
        signal oVar1S867: std_logic_vector(   0 downto 0);
        signal oVar1S868: std_logic_vector(   0 downto 0);
        signal oVar1S869: std_logic_vector(   0 downto 0);
        signal oVar1S870: std_logic_vector(   0 downto 0);
        signal oVar1S871: std_logic_vector(   0 downto 0);
        signal oVar1S872: std_logic_vector(   0 downto 0);
        signal oVar1S873: std_logic_vector(   0 downto 0);
        signal oVar1S874: std_logic_vector(   0 downto 0);
        signal oVar1S876: std_logic_vector(   0 downto 0);
        signal oVar1S877: std_logic_vector(   0 downto 0);
        signal oVar1S878: std_logic_vector(   0 downto 0);
        signal oVar1S879: std_logic_vector(   0 downto 0);
        signal oVar1S880: std_logic_vector(   0 downto 0);
        signal oVar1S881: std_logic_vector(   0 downto 0);
        signal oVar1S882: std_logic_vector(   0 downto 0);
        signal oVar1S883: std_logic_vector(   0 downto 0);
        signal oVar1S884: std_logic_vector(   0 downto 0);
        signal oVar1S885: std_logic_vector(   0 downto 0);
        signal oVar1S886: std_logic_vector(   0 downto 0);
        signal oVar1S887: std_logic_vector(   0 downto 0);
        signal oVar1S888: std_logic_vector(   0 downto 0);
        signal oVar1S889: std_logic_vector(   0 downto 0);
        signal oVar1S890: std_logic_vector(   0 downto 0);
        signal oVar1S891: std_logic_vector(   0 downto 0);
        signal oVar1S892: std_logic_vector(   0 downto 0);
        signal oVar1S893: std_logic_vector(   0 downto 0);
        signal oVar1S894: std_logic_vector(   0 downto 0);
        signal oVar1S895: std_logic_vector(   0 downto 0);
        signal oVar1S896: std_logic_vector(   0 downto 0);
        signal oVar1S897: std_logic_vector(   0 downto 0);
        signal oVar1S898: std_logic_vector(   0 downto 0);
        signal oVar1S899: std_logic_vector(   0 downto 0);
        signal oVar1S900: std_logic_vector(   0 downto 0);
        signal oVar1S901: std_logic_vector(   0 downto 0);
        signal oVar1S902: std_logic_vector(   0 downto 0);
        signal oVar1S903: std_logic_vector(   0 downto 0);
        signal oVar1S904: std_logic_vector(   0 downto 0);
        signal oVar1S905: std_logic_vector(   0 downto 0);
        signal oVar1S906: std_logic_vector(   0 downto 0);
        signal oVar1S907: std_logic_vector(   0 downto 0);
        signal oVar1S908: std_logic_vector(   0 downto 0);
        signal oVar1S909: std_logic_vector(   0 downto 0);
        signal oVar1S910: std_logic_vector(   0 downto 0);
        signal oVar1S911: std_logic_vector(   0 downto 0);
        signal oVar1S913: std_logic_vector(   0 downto 0);
        signal oVar1S914: std_logic_vector(   0 downto 0);
        signal oVar1S915: std_logic_vector(   0 downto 0);
        signal oVar1S916: std_logic_vector(   0 downto 0);
        signal oVar1S917: std_logic_vector(   0 downto 0);
        signal oVar1S918: std_logic_vector(   0 downto 0);
        signal oVar1S919: std_logic_vector(   0 downto 0);
        signal oVar1S920: std_logic_vector(   0 downto 0);
        signal oVar1S922: std_logic_vector(   0 downto 0);
        signal oVar1S923: std_logic_vector(   0 downto 0);
        signal oVar1S924: std_logic_vector(   0 downto 0);
        signal oVar1S925: std_logic_vector(   0 downto 0);
        signal oVar1S926: std_logic_vector(   0 downto 0);
        signal oVar1S927: std_logic_vector(   0 downto 0);
        signal oVar1S928: std_logic_vector(   0 downto 0);
        signal oVar1S929: std_logic_vector(   0 downto 0);
        signal oVar1S930: std_logic_vector(   0 downto 0);
        signal oVar1S931: std_logic_vector(   0 downto 0);
        signal oVar1S932: std_logic_vector(   0 downto 0);
        signal oVar1S933: std_logic_vector(   0 downto 0);
        signal oVar1S934: std_logic_vector(   0 downto 0);
        signal oVar1S935: std_logic_vector(   0 downto 0);
        signal oVar1S937: std_logic_vector(   0 downto 0);
        signal oVar1S938: std_logic_vector(   0 downto 0);
        signal oVar1S939: std_logic_vector(   0 downto 0);
        signal oVar1S940: std_logic_vector(   0 downto 0);
        signal oVar1S941: std_logic_vector(   0 downto 0);
        signal oVar1S942: std_logic_vector(   0 downto 0);
        signal oVar1S943: std_logic_vector(   0 downto 0);
        signal oVar1S944: std_logic_vector(   0 downto 0);
        signal oVar1S945: std_logic_vector(   0 downto 0);
        signal oVar1S946: std_logic_vector(   0 downto 0);
        signal oVar1S947: std_logic_vector(   0 downto 0);
        signal oVar1S948: std_logic_vector(   0 downto 0);
        signal oVar1S949: std_logic_vector(   0 downto 0);
        signal oVar1S950: std_logic_vector(   0 downto 0);
        signal oVar1S951: std_logic_vector(   0 downto 0);
        signal oVar1S952: std_logic_vector(   0 downto 0);
        signal oVar1S954: std_logic_vector(   0 downto 0);
        signal oVar1S955: std_logic_vector(   0 downto 0);
        signal oVar1S956: std_logic_vector(   0 downto 0);
        signal oVar1S957: std_logic_vector(   0 downto 0);
        signal oVar1S958: std_logic_vector(   0 downto 0);
        signal oVar1S959: std_logic_vector(   0 downto 0);
        signal oVar1S960: std_logic_vector(   0 downto 0);
        signal oVar1S961: std_logic_vector(   0 downto 0);
        signal oVar1S962: std_logic_vector(   0 downto 0);
        signal oVar1S963: std_logic_vector(   0 downto 0);
        signal oVar1S964: std_logic_vector(   0 downto 0);
        signal oVar1S965: std_logic_vector(   0 downto 0);
        signal oVar1S966: std_logic_vector(   0 downto 0);
        signal oVar1S967: std_logic_vector(   0 downto 0);
        signal oVar1S968: std_logic_vector(   0 downto 0);
        signal oVar1S969: std_logic_vector(   0 downto 0);
        signal oVar1S970: std_logic_vector(   0 downto 0);
        signal oVar1S971: std_logic_vector(   0 downto 0);
        signal oVar1S972: std_logic_vector(   0 downto 0);
        signal oVar1S974: std_logic_vector(   0 downto 0);
        signal oVar1S975: std_logic_vector(   0 downto 0);
        signal oVar1S976: std_logic_vector(   0 downto 0);
        signal oVar1S977: std_logic_vector(   0 downto 0);
        signal oVar1S978: std_logic_vector(   0 downto 0);
        signal oVar1S979: std_logic_vector(   0 downto 0);
        signal oVar1S980: std_logic_vector(   0 downto 0);
        signal oVar1S981: std_logic_vector(   0 downto 0);
        signal oVar1S982: std_logic_vector(   0 downto 0);
        signal oVar1S983: std_logic_vector(   0 downto 0);
        signal oVar1S984: std_logic_vector(   0 downto 0);
        signal oVar1S985: std_logic_vector(   0 downto 0);
        signal oVar1S986: std_logic_vector(   0 downto 0);
        signal oVar1S987: std_logic_vector(   0 downto 0);
        signal oVar1S988: std_logic_vector(   0 downto 0);
        signal oVar1S990: std_logic_vector(   0 downto 0);
        signal oVar1S991: std_logic_vector(   0 downto 0);
        signal oVar1S992: std_logic_vector(   0 downto 0);
        signal oVar1S993: std_logic_vector(   0 downto 0);
        signal oVar1S994: std_logic_vector(   0 downto 0);
        signal oVar1S995: std_logic_vector(   0 downto 0);
        signal oVar1S996: std_logic_vector(   0 downto 0);
        signal oVar1S998: std_logic_vector(   0 downto 0);
        signal oVar1S999: std_logic_vector(   0 downto 0);
        signal oVar1S1000: std_logic_vector(   0 downto 0);
        signal oVar1S1001: std_logic_vector(   0 downto 0);
        signal oVar1S1002: std_logic_vector(   0 downto 0);
        signal oVar1S1003: std_logic_vector(   0 downto 0);
        signal oVar1S1004: std_logic_vector(   0 downto 0);
        signal oVar1S1005: std_logic_vector(   0 downto 0);
        signal oVar1S1006: std_logic_vector(   0 downto 0);
        signal oVar1S1007: std_logic_vector(   0 downto 0);
        signal oVar1S1008: std_logic_vector(   0 downto 0);
        signal oVar1S1009: std_logic_vector(   0 downto 0);
        signal oVar1S1010: std_logic_vector(   0 downto 0);
        signal oVar1S1011: std_logic_vector(   0 downto 0);
        signal oVar1S1012: std_logic_vector(   0 downto 0);
        signal oVar1S1013: std_logic_vector(   0 downto 0);
        signal oVar1S1014: std_logic_vector(   0 downto 0);
        signal oVar1S1015: std_logic_vector(   0 downto 0);
        signal oVar1S1016: std_logic_vector(   0 downto 0);
        signal oVar1S1017: std_logic_vector(   0 downto 0);
        signal oVar1S1018: std_logic_vector(   0 downto 0);
        signal oVar1S1019: std_logic_vector(   0 downto 0);
        signal oVar1S1020: std_logic_vector(   0 downto 0);
        signal oVar1S1021: std_logic_vector(   0 downto 0);
        signal oVar1S1022: std_logic_vector(   0 downto 0);
        signal oVar1S1023: std_logic_vector(   0 downto 0);
        signal oVar1S1024: std_logic_vector(   0 downto 0);
        signal oVar1S1025: std_logic_vector(   0 downto 0);
        signal oVar1S1026: std_logic_vector(   0 downto 0);
        signal oVar1S1027: std_logic_vector(   0 downto 0);
        signal oVar1S1028: std_logic_vector(   0 downto 0);
        signal oVar1S1029: std_logic_vector(   0 downto 0);
        signal oVar1S1030: std_logic_vector(   0 downto 0);
        signal oVar1S1031: std_logic_vector(   0 downto 0);
        signal oVar1S1032: std_logic_vector(   0 downto 0);
        signal oVar1S1033: std_logic_vector(   0 downto 0);
        signal oVar1S1034: std_logic_vector(   0 downto 0);
        signal oVar1S1035: std_logic_vector(   0 downto 0);
        signal oVar1S1036: std_logic_vector(   0 downto 0);
        signal oVar1S1037: std_logic_vector(   0 downto 0);
        signal oVar1S1038: std_logic_vector(   0 downto 0);
        signal oVar1S1039: std_logic_vector(   0 downto 0);
        signal oVar1S1040: std_logic_vector(   0 downto 0);
        signal oVar1S1041: std_logic_vector(   0 downto 0);
        signal oVar1S1042: std_logic_vector(   0 downto 0);
        signal oVar1S1043: std_logic_vector(   0 downto 0);
        signal oVar1S1044: std_logic_vector(   0 downto 0);
        signal oVar1S1045: std_logic_vector(   0 downto 0);
        signal oVar1S1046: std_logic_vector(   0 downto 0);
        signal oVar1S1047: std_logic_vector(   0 downto 0);
        signal oVar1S1048: std_logic_vector(   0 downto 0);
        signal oVar1S1049: std_logic_vector(   0 downto 0);
        signal oVar1S1050: std_logic_vector(   0 downto 0);
        signal oVar1S1051: std_logic_vector(   0 downto 0);
        signal oVar1S1052: std_logic_vector(   0 downto 0);
        signal oVar1S1053: std_logic_vector(   0 downto 0);
        signal oVar1S1054: std_logic_vector(   0 downto 0);
        signal oVar1S1055: std_logic_vector(   0 downto 0);
        signal oVar1S1056: std_logic_vector(   0 downto 0);
        signal oVar1S1057: std_logic_vector(   0 downto 0);
        signal oVar1S1058: std_logic_vector(   0 downto 0);
        signal oVar1S1059: std_logic_vector(   0 downto 0);
        signal oVar1S1060: std_logic_vector(   0 downto 0);
        signal oVar1S1062: std_logic_vector(   0 downto 0);
        signal oVar1S1063: std_logic_vector(   0 downto 0);
        signal oVar1S1064: std_logic_vector(   0 downto 0);
        signal oVar1S1065: std_logic_vector(   0 downto 0);
        signal oVar1S1066: std_logic_vector(   0 downto 0);
        signal oVar1S1067: std_logic_vector(   0 downto 0);
        signal oVar1S1068: std_logic_vector(   0 downto 0);
        signal oVar1S1069: std_logic_vector(   0 downto 0);
        signal oVar1S1071: std_logic_vector(   0 downto 0);
        signal oVar1S1072: std_logic_vector(   0 downto 0);
        signal oVar1S1073: std_logic_vector(   0 downto 0);
        signal oVar1S1074: std_logic_vector(   0 downto 0);
        signal oVar1S1075: std_logic_vector(   0 downto 0);
        signal oVar1S1076: std_logic_vector(   0 downto 0);
        signal oVar1S1077: std_logic_vector(   0 downto 0);
        signal oVar1S1078: std_logic_vector(   0 downto 0);
        signal oVar1S1079: std_logic_vector(   0 downto 0);
        signal oVar1S1081: std_logic_vector(   0 downto 0);
        signal oVar1S1082: std_logic_vector(   0 downto 0);
        signal oVar1S1083: std_logic_vector(   0 downto 0);
        signal oVar1S1084: std_logic_vector(   0 downto 0);
        signal oVar1S1085: std_logic_vector(   0 downto 0);
        signal oVar1S1086: std_logic_vector(   0 downto 0);
        signal oVar1S1087: std_logic_vector(   0 downto 0);
        signal oVar1S1088: std_logic_vector(   0 downto 0);
        signal oVar1S1089: std_logic_vector(   0 downto 0);
        signal oVar1S1090: std_logic_vector(   0 downto 0);
        signal oVar1S1091: std_logic_vector(   0 downto 0);
        signal oVar1S1092: std_logic_vector(   0 downto 0);
        signal oVar1S1093: std_logic_vector(   0 downto 0);
        signal oVar1S1094: std_logic_vector(   0 downto 0);
        signal oVar1S1095: std_logic_vector(   0 downto 0);
        signal oVar1S1096: std_logic_vector(   0 downto 0);
        signal oVar1S1097: std_logic_vector(   0 downto 0);
        signal oVar1S1098: std_logic_vector(   0 downto 0);
        signal oVar1S1099: std_logic_vector(   0 downto 0);
        signal oVar1S1100: std_logic_vector(   0 downto 0);
        signal oVar1S1101: std_logic_vector(   0 downto 0);
        signal oVar1S1102: std_logic_vector(   0 downto 0);
        signal oVar1S1103: std_logic_vector(   0 downto 0);
        signal oVar1S1104: std_logic_vector(   0 downto 0);
        signal oVar1S1105: std_logic_vector(   0 downto 0);
        signal oVar1S1107: std_logic_vector(   0 downto 0);
        signal oVar1S1108: std_logic_vector(   0 downto 0);
        signal oVar1S1109: std_logic_vector(   0 downto 0);
        signal oVar1S1110: std_logic_vector(   0 downto 0);
        signal oVar1S1111: std_logic_vector(   0 downto 0);
        signal oVar1S1112: std_logic_vector(   0 downto 0);
        signal oVar1S1113: std_logic_vector(   0 downto 0);
        signal oVar1S1114: std_logic_vector(   0 downto 0);
        signal oVar1S1115: std_logic_vector(   0 downto 0);
        signal oVar1S1116: std_logic_vector(   0 downto 0);
        signal oVar1S1117: std_logic_vector(   0 downto 0);
        signal oVar1S1119: std_logic_vector(   0 downto 0);
        signal oVar1S1120: std_logic_vector(   0 downto 0);
        signal oVar1S1121: std_logic_vector(   0 downto 0);
        signal oVar1S1122: std_logic_vector(   0 downto 0);
        signal oVar1S1123: std_logic_vector(   0 downto 0);
        signal oVar1S1124: std_logic_vector(   0 downto 0);
        signal oVar1S1125: std_logic_vector(   0 downto 0);
        signal oVar1S1126: std_logic_vector(   0 downto 0);
        signal oVar1S1128: std_logic_vector(   0 downto 0);
        signal oVar1S1129: std_logic_vector(   0 downto 0);
        signal oVar1S1130: std_logic_vector(   0 downto 0);
        signal oVar1S1131: std_logic_vector(   0 downto 0);
        signal oVar1S1132: std_logic_vector(   0 downto 0);
        signal oVar1S1133: std_logic_vector(   0 downto 0);
        signal oVar1S1134: std_logic_vector(   0 downto 0);
        signal oVar1S1135: std_logic_vector(   0 downto 0);
        signal oVar1S1136: std_logic_vector(   0 downto 0);
        signal oVar1S1137: std_logic_vector(   0 downto 0);
        signal oVar1S1138: std_logic_vector(   0 downto 0);
        signal oVar1S1139: std_logic_vector(   0 downto 0);
        signal oVar1S1140: std_logic_vector(   0 downto 0);
        signal oVar1S1141: std_logic_vector(   0 downto 0);
        signal oVar1S1142: std_logic_vector(   0 downto 0);
        signal oVar1S1143: std_logic_vector(   0 downto 0);
        signal oVar1S1144: std_logic_vector(   0 downto 0);
        signal oVar1S1145: std_logic_vector(   0 downto 0);
        signal oVar1S1146: std_logic_vector(   0 downto 0);
        signal oVar1S1147: std_logic_vector(   0 downto 0);
        signal oVar1S1148: std_logic_vector(   0 downto 0);
        signal oVar1S1149: std_logic_vector(   0 downto 0);
        signal oVar1S1150: std_logic_vector(   0 downto 0);
        signal oVar1S1151: std_logic_vector(   0 downto 0);
        signal oVar1S1152: std_logic_vector(   0 downto 0);
        signal oVar1S1153: std_logic_vector(   0 downto 0);
        signal oVar1S1154: std_logic_vector(   0 downto 0);
        signal oVar1S1155: std_logic_vector(   0 downto 0);
        signal oVar1S1156: std_logic_vector(   0 downto 0);
        signal oVar1S1157: std_logic_vector(   0 downto 0);
        signal oVar2S0: std_logic_vector(   0 downto 0);
        signal oVar2S1: std_logic_vector(   0 downto 0);
        signal oVar2S2: std_logic_vector(   0 downto 0);
        signal oVar2S3: std_logic_vector(   0 downto 0);
        signal oVar2S4: std_logic_vector(   0 downto 0);
        signal oVar2S6: std_logic_vector(   0 downto 0);
        signal oVar2S7: std_logic_vector(   0 downto 0);
        signal oVar2S8: std_logic_vector(   0 downto 0);
        signal oVar2S9: std_logic_vector(   0 downto 0);
        signal oVar2S10: std_logic_vector(   0 downto 0);
        signal oVar2S12: std_logic_vector(   0 downto 0);
        signal oVar2S13: std_logic_vector(   0 downto 0);
        signal oVar2S15: std_logic_vector(   0 downto 0);
        signal oVar2S16: std_logic_vector(   0 downto 0);
        signal oVar2S17: std_logic_vector(   0 downto 0);
        signal oVar2S18: std_logic_vector(   0 downto 0);
        signal oVar2S19: std_logic_vector(   0 downto 0);
        signal oVar2S20: std_logic_vector(   0 downto 0);
        signal oVar2S21: std_logic_vector(   0 downto 0);
        signal oVar2S23: std_logic_vector(   0 downto 0);
        signal oVar2S24: std_logic_vector(   0 downto 0);
        signal oVar2S25: std_logic_vector(   0 downto 0);
        signal oVar2S26: std_logic_vector(   0 downto 0);
        signal oVar2S27: std_logic_vector(   0 downto 0);
        signal oVar2S28: std_logic_vector(   0 downto 0);
        signal oVar2S29: std_logic_vector(   0 downto 0);
        signal oVar2S30: std_logic_vector(   0 downto 0);
        signal oVar2S31: std_logic_vector(   0 downto 0);
        signal oVar2S32: std_logic_vector(   0 downto 0);
        signal oVar2S33: std_logic_vector(   0 downto 0);
        signal oVar2S34: std_logic_vector(   0 downto 0);
        signal oVar2S35: std_logic_vector(   0 downto 0);
        signal oVar2S36: std_logic_vector(   0 downto 0);
        signal oVar2S37: std_logic_vector(   0 downto 0);
        signal oVar2S38: std_logic_vector(   0 downto 0);
        signal oVar2S39: std_logic_vector(   0 downto 0);
        signal oVar2S40: std_logic_vector(   0 downto 0);
        signal oVar2S41: std_logic_vector(   0 downto 0);
        signal oVar2S42: std_logic_vector(   0 downto 0);
        signal oVar2S43: std_logic_vector(   0 downto 0);
        signal oVar2S45: std_logic_vector(   0 downto 0);
        signal oVar2S46: std_logic_vector(   0 downto 0);
        signal oVar2S48: std_logic_vector(   0 downto 0);
        signal oVar2S49: std_logic_vector(   0 downto 0);
        signal oVar2S50: std_logic_vector(   0 downto 0);
        signal oVar2S51: std_logic_vector(   0 downto 0);
        signal oVar2S52: std_logic_vector(   0 downto 0);
        signal oVar2S53: std_logic_vector(   0 downto 0);
        signal oVar2S54: std_logic_vector(   0 downto 0);
        signal oVar2S55: std_logic_vector(   0 downto 0);
        signal oVar2S56: std_logic_vector(   0 downto 0);
        signal oVar2S57: std_logic_vector(   0 downto 0);
        signal oVar2S58: std_logic_vector(   0 downto 0);
        signal oVar2S59: std_logic_vector(   0 downto 0);
        signal oVar2S60: std_logic_vector(   0 downto 0);
        signal oVar2S61: std_logic_vector(   0 downto 0);
        signal oVar2S62: std_logic_vector(   0 downto 0);
        signal oVar2S63: std_logic_vector(   0 downto 0);
        signal oVar2S64: std_logic_vector(   0 downto 0);
        signal oVar2S66: std_logic_vector(   0 downto 0);
        signal oVar2S67: std_logic_vector(   0 downto 0);
        signal oVar2S68: std_logic_vector(   0 downto 0);
        signal oVar2S69: std_logic_vector(   0 downto 0);
        signal oVar2S71: std_logic_vector(   0 downto 0);
        signal oVar2S72: std_logic_vector(   0 downto 0);
        signal oVar2S74: std_logic_vector(   0 downto 0);
        signal oVar2S75: std_logic_vector(   0 downto 0);
        signal oVar2S76: std_logic_vector(   0 downto 0);
        signal oVar2S77: std_logic_vector(   0 downto 0);
        signal oVar2S78: std_logic_vector(   0 downto 0);
        signal oVar2S79: std_logic_vector(   0 downto 0);
        signal oVar2S80: std_logic_vector(   0 downto 0);
        signal oVar2S81: std_logic_vector(   0 downto 0);
        signal oVar2S82: std_logic_vector(   0 downto 0);
        signal oVar2S83: std_logic_vector(   0 downto 0);
        signal oVar2S84: std_logic_vector(   0 downto 0);
        signal oVar2S85: std_logic_vector(   0 downto 0);
        signal oVar2S86: std_logic_vector(   0 downto 0);
        signal oVar2S87: std_logic_vector(   0 downto 0);
        signal oVar2S88: std_logic_vector(   0 downto 0);
        signal oVar2S90: std_logic_vector(   0 downto 0);
        signal oVar2S91: std_logic_vector(   0 downto 0);
        signal oVar2S92: std_logic_vector(   0 downto 0);
        signal oVar2S93: std_logic_vector(   0 downto 0);
        signal oVar2S94: std_logic_vector(   0 downto 0);
        signal oVar2S96: std_logic_vector(   0 downto 0);
        signal oVar2S97: std_logic_vector(   0 downto 0);
        signal oVar2S98: std_logic_vector(   0 downto 0);
        signal oVar2S100: std_logic_vector(   0 downto 0);
        signal oVar2S101: std_logic_vector(   0 downto 0);
        signal oVar2S103: std_logic_vector(   0 downto 0);
        signal oVar2S104: std_logic_vector(   0 downto 0);
        signal oVar2S105: std_logic_vector(   0 downto 0);
        signal oVar2S106: std_logic_vector(   0 downto 0);
        signal oVar2S107: std_logic_vector(   0 downto 0);
        signal oVar2S108: std_logic_vector(   0 downto 0);
        signal oVar2S109: std_logic_vector(   0 downto 0);
        signal oVar2S110: std_logic_vector(   0 downto 0);
        signal oVar2S111: std_logic_vector(   0 downto 0);
        signal oVar2S112: std_logic_vector(   0 downto 0);
        signal oVar2S113: std_logic_vector(   0 downto 0);
        signal oVar2S114: std_logic_vector(   0 downto 0);
        signal oVar2S115: std_logic_vector(   0 downto 0);
        signal oVar2S116: std_logic_vector(   0 downto 0);
        signal oVar2S117: std_logic_vector(   0 downto 0);
        signal oVar2S118: std_logic_vector(   0 downto 0);
        signal oVar2S119: std_logic_vector(   0 downto 0);
        signal oVar2S121: std_logic_vector(   0 downto 0);
        signal oVar2S122: std_logic_vector(   0 downto 0);
        signal oVar2S123: std_logic_vector(   0 downto 0);
        signal oVar2S124: std_logic_vector(   0 downto 0);
        signal oVar2S125: std_logic_vector(   0 downto 0);
        signal oVar2S126: std_logic_vector(   0 downto 0);
        signal oVar2S127: std_logic_vector(   0 downto 0);
        signal oVar2S128: std_logic_vector(   0 downto 0);
        signal oVar2S129: std_logic_vector(   0 downto 0);
        signal oVar2S130: std_logic_vector(   0 downto 0);
        signal oVar2S132: std_logic_vector(   0 downto 0);
        signal oVar2S133: std_logic_vector(   0 downto 0);
        signal oVar2S134: std_logic_vector(   0 downto 0);
        signal oVar2S135: std_logic_vector(   0 downto 0);
        signal oVar2S136: std_logic_vector(   0 downto 0);
        signal oVar2S137: std_logic_vector(   0 downto 0);
        signal oVar2S138: std_logic_vector(   0 downto 0);
        signal oVar2S139: std_logic_vector(   0 downto 0);
        signal oVar2S141: std_logic_vector(   0 downto 0);
        signal oVar2S142: std_logic_vector(   0 downto 0);
        signal oVar2S144: std_logic_vector(   0 downto 0);
        signal oVar2S145: std_logic_vector(   0 downto 0);
        signal oVar2S146: std_logic_vector(   0 downto 0);
        signal oVar2S147: std_logic_vector(   0 downto 0);
        signal oVar2S148: std_logic_vector(   0 downto 0);
        signal oVar2S150: std_logic_vector(   0 downto 0);
        signal oVar2S151: std_logic_vector(   0 downto 0);
        signal oVar2S153: std_logic_vector(   0 downto 0);
        signal oVar2S154: std_logic_vector(   0 downto 0);
        signal oVar2S155: std_logic_vector(   0 downto 0);
        signal oVar2S156: std_logic_vector(   0 downto 0);
        signal oVar2S157: std_logic_vector(   0 downto 0);
        signal oVar2S158: std_logic_vector(   0 downto 0);
        signal oVar2S159: std_logic_vector(   0 downto 0);
        signal oVar2S160: std_logic_vector(   0 downto 0);
        signal oVar2S162: std_logic_vector(   0 downto 0);
        signal oVar2S163: std_logic_vector(   0 downto 0);
        signal oVar2S165: std_logic_vector(   0 downto 0);
        signal oVar2S166: std_logic_vector(   0 downto 0);
        signal oVar2S168: std_logic_vector(   0 downto 0);
        signal oVar2S169: std_logic_vector(   0 downto 0);
        signal oVar2S170: std_logic_vector(   0 downto 0);
        signal oVar2S171: std_logic_vector(   0 downto 0);
        signal oVar2S172: std_logic_vector(   0 downto 0);
        signal oVar2S173: std_logic_vector(   0 downto 0);
        signal oVar2S174: std_logic_vector(   0 downto 0);
        signal oVar2S175: std_logic_vector(   0 downto 0);
        signal oVar2S176: std_logic_vector(   0 downto 0);
        signal oVar2S177: std_logic_vector(   0 downto 0);
        signal oVar2S178: std_logic_vector(   0 downto 0);
        signal oVar2S179: std_logic_vector(   0 downto 0);
        signal oVar2S180: std_logic_vector(   0 downto 0);
        signal oVar2S181: std_logic_vector(   0 downto 0);
        signal oVar2S182: std_logic_vector(   0 downto 0);
        signal oVar2S183: std_logic_vector(   0 downto 0);
        signal oVar2S185: std_logic_vector(   0 downto 0);
        signal oVar2S186: std_logic_vector(   0 downto 0);
        signal oVar2S187: std_logic_vector(   0 downto 0);
        signal oVar2S188: std_logic_vector(   0 downto 0);
        signal oVar2S190: std_logic_vector(   0 downto 0);
        signal oVar2S191: std_logic_vector(   0 downto 0);
        signal oVar2S192: std_logic_vector(   0 downto 0);
        signal oVar2S193: std_logic_vector(   0 downto 0);
        signal oVar2S194: std_logic_vector(   0 downto 0);
        signal oVar2S196: std_logic_vector(   0 downto 0);
        signal oVar2S197: std_logic_vector(   0 downto 0);
        signal oVar2S198: std_logic_vector(   0 downto 0);
        signal oVar2S199: std_logic_vector(   0 downto 0);
        signal oVar2S200: std_logic_vector(   0 downto 0);
        signal oVar2S201: std_logic_vector(   0 downto 0);
        signal oVar2S203: std_logic_vector(   0 downto 0);
        signal oVar2S204: std_logic_vector(   0 downto 0);
        signal oVar2S206: std_logic_vector(   0 downto 0);
        signal oVar2S207: std_logic_vector(   0 downto 0);
        signal oVar2S208: std_logic_vector(   0 downto 0);
        signal oVar2S209: std_logic_vector(   0 downto 0);
        signal oVar2S210: std_logic_vector(   0 downto 0);
        signal oVar2S212: std_logic_vector(   0 downto 0);
        signal oVar2S213: std_logic_vector(   0 downto 0);
        signal oVar2S215: std_logic_vector(   0 downto 0);
        signal oVar2S216: std_logic_vector(   0 downto 0);
        signal oVar2S218: std_logic_vector(   0 downto 0);
        signal oVar2S219: std_logic_vector(   0 downto 0);
        signal oVar2S220: std_logic_vector(   0 downto 0);
        signal oVar2S221: std_logic_vector(   0 downto 0);
        signal oVar2S222: std_logic_vector(   0 downto 0);
        signal oVar2S223: std_logic_vector(   0 downto 0);
        signal oVar2S224: std_logic_vector(   0 downto 0);
        signal oVar2S225: std_logic_vector(   0 downto 0);
        signal oVar2S227: std_logic_vector(   0 downto 0);
        signal oVar2S228: std_logic_vector(   0 downto 0);
        signal oVar2S229: std_logic_vector(   0 downto 0);
        signal oVar2S230: std_logic_vector(   0 downto 0);
        signal oVar2S231: std_logic_vector(   0 downto 0);
        signal oVar2S233: std_logic_vector(   0 downto 0);
        signal oVar2S234: std_logic_vector(   0 downto 0);
        signal oVar2S235: std_logic_vector(   0 downto 0);
        signal oVar2S236: std_logic_vector(   0 downto 0);
        signal oVar2S237: std_logic_vector(   0 downto 0);
        signal oVar2S238: std_logic_vector(   0 downto 0);
        signal oVar2S239: std_logic_vector(   0 downto 0);
        signal oVar2S240: std_logic_vector(   0 downto 0);
        signal oVar2S241: std_logic_vector(   0 downto 0);
        signal oVar2S242: std_logic_vector(   0 downto 0);
        signal oVar2S243: std_logic_vector(   0 downto 0);
        signal oVar2S244: std_logic_vector(   0 downto 0);
        signal oVar2S245: std_logic_vector(   0 downto 0);
        signal oVar2S246: std_logic_vector(   0 downto 0);
        signal oVar2S247: std_logic_vector(   0 downto 0);
        signal oVar2S248: std_logic_vector(   0 downto 0);
        signal oVar2S249: std_logic_vector(   0 downto 0);
        signal oVar2S250: std_logic_vector(   0 downto 0);
        signal oVar2S251: std_logic_vector(   0 downto 0);
        signal oVar2S252: std_logic_vector(   0 downto 0);
        signal oVar2S253: std_logic_vector(   0 downto 0);
        signal oVar2S254: std_logic_vector(   0 downto 0);
        signal oVar2S255: std_logic_vector(   0 downto 0);
        signal oVar2S256: std_logic_vector(   0 downto 0);
        signal oVar2S257: std_logic_vector(   0 downto 0);
        signal oVar2S258: std_logic_vector(   0 downto 0);
        signal oVar2S259: std_logic_vector(   0 downto 0);
        signal oVar2S260: std_logic_vector(   0 downto 0);
        signal oVar2S261: std_logic_vector(   0 downto 0);
        signal oVar2S262: std_logic_vector(   0 downto 0);
        signal oVar2S264: std_logic_vector(   0 downto 0);
        signal oVar2S265: std_logic_vector(   0 downto 0);
        signal oVar2S267: std_logic_vector(   0 downto 0);
        signal oVar2S268: std_logic_vector(   0 downto 0);
        signal oVar2S269: std_logic_vector(   0 downto 0);
        signal oVar2S270: std_logic_vector(   0 downto 0);
        signal oVar2S271: std_logic_vector(   0 downto 0);
        signal oVar2S272: std_logic_vector(   0 downto 0);
        signal oVar2S273: std_logic_vector(   0 downto 0);
        signal oVar2S274: std_logic_vector(   0 downto 0);
        signal oVar2S275: std_logic_vector(   0 downto 0);
        signal oVar2S276: std_logic_vector(   0 downto 0);
        signal oVar2S277: std_logic_vector(   0 downto 0);
        signal oVar2S278: std_logic_vector(   0 downto 0);
        signal oVar2S279: std_logic_vector(   0 downto 0);
        signal oVar2S280: std_logic_vector(   0 downto 0);
        signal oVar2S281: std_logic_vector(   0 downto 0);
        signal oVar2S282: std_logic_vector(   0 downto 0);
        signal oVar2S283: std_logic_vector(   0 downto 0);
        signal oVar2S285: std_logic_vector(   0 downto 0);
        signal oVar2S286: std_logic_vector(   0 downto 0);
        signal oVar2S288: std_logic_vector(   0 downto 0);
        signal oVar2S289: std_logic_vector(   0 downto 0);
        signal oVar2S290: std_logic_vector(   0 downto 0);
        signal oVar2S291: std_logic_vector(   0 downto 0);
        signal oVar2S292: std_logic_vector(   0 downto 0);
        signal oVar2S293: std_logic_vector(   0 downto 0);
        signal oVar2S294: std_logic_vector(   0 downto 0);
        signal oVar2S295: std_logic_vector(   0 downto 0);
        signal oVar2S297: std_logic_vector(   0 downto 0);
        signal oVar2S298: std_logic_vector(   0 downto 0);
        signal oVar2S300: std_logic_vector(   0 downto 0);
        signal oVar2S301: std_logic_vector(   0 downto 0);
        signal oVar2S303: std_logic_vector(   0 downto 0);
        signal oVar2S304: std_logic_vector(   0 downto 0);
        signal oVar2S305: std_logic_vector(   0 downto 0);
        signal oVar2S306: std_logic_vector(   0 downto 0);
        signal oVar2S308: std_logic_vector(   0 downto 0);
        signal oVar2S309: std_logic_vector(   0 downto 0);
        signal oVar2S311: std_logic_vector(   0 downto 0);
        signal oVar2S312: std_logic_vector(   0 downto 0);
        signal oVar2S313: std_logic_vector(   0 downto 0);
        signal oVar2S314: std_logic_vector(   0 downto 0);
        signal oVar2S315: std_logic_vector(   0 downto 0);
        signal oVar2S316: std_logic_vector(   0 downto 0);
        signal oVar2S317: std_logic_vector(   0 downto 0);
        signal oVar2S318: std_logic_vector(   0 downto 0);
        signal oVar2S320: std_logic_vector(   0 downto 0);
        signal oVar2S321: std_logic_vector(   0 downto 0);
        signal oVar2S323: std_logic_vector(   0 downto 0);
        signal oVar2S324: std_logic_vector(   0 downto 0);
        signal oVar2S326: std_logic_vector(   0 downto 0);
        signal oVar2S327: std_logic_vector(   0 downto 0);
        signal oVar2S328: std_logic_vector(   0 downto 0);
        signal oVar2S329: std_logic_vector(   0 downto 0);
        signal oVar2S330: std_logic_vector(   0 downto 0);
        signal oVar2S331: std_logic_vector(   0 downto 0);
        signal oVar2S333: std_logic_vector(   0 downto 0);
        signal oVar2S334: std_logic_vector(   0 downto 0);
        signal oVar2S335: std_logic_vector(   0 downto 0);
        signal oVar2S336: std_logic_vector(   0 downto 0);
        signal oVar2S337: std_logic_vector(   0 downto 0);
        signal oVar2S338: std_logic_vector(   0 downto 0);
        signal oVar2S339: std_logic_vector(   0 downto 0);
        signal oVar2S340: std_logic_vector(   0 downto 0);
        signal oVar2S341: std_logic_vector(   0 downto 0);
        signal oVar2S342: std_logic_vector(   0 downto 0);
        signal oVar2S343: std_logic_vector(   0 downto 0);
        signal oVar2S344: std_logic_vector(   0 downto 0);
        signal oVar2S345: std_logic_vector(   0 downto 0);
        signal oVar2S346: std_logic_vector(   0 downto 0);
        signal oVar2S348: std_logic_vector(   0 downto 0);
        signal oVar2S349: std_logic_vector(   0 downto 0);
        signal oVar2S350: std_logic_vector(   0 downto 0);
        signal oVar2S351: std_logic_vector(   0 downto 0);
        signal oVar2S352: std_logic_vector(   0 downto 0);
        signal oVar2S353: std_logic_vector(   0 downto 0);
        signal oVar2S354: std_logic_vector(   0 downto 0);
        signal oVar2S355: std_logic_vector(   0 downto 0);
        signal oVar2S356: std_logic_vector(   0 downto 0);
        signal oVar2S357: std_logic_vector(   0 downto 0);
        signal oVar2S358: std_logic_vector(   0 downto 0);
        signal oVar2S359: std_logic_vector(   0 downto 0);
        signal oVar2S360: std_logic_vector(   0 downto 0);
        signal oVar2S361: std_logic_vector(   0 downto 0);
        signal oVar2S363: std_logic_vector(   0 downto 0);
        signal oVar2S364: std_logic_vector(   0 downto 0);
        signal oVar2S366: std_logic_vector(   0 downto 0);
        signal oVar2S367: std_logic_vector(   0 downto 0);
        signal oVar2S368: std_logic_vector(   0 downto 0);
        signal oVar2S369: std_logic_vector(   0 downto 0);
        signal oVar2S370: std_logic_vector(   0 downto 0);
        signal oVar2S371: std_logic_vector(   0 downto 0);
        signal oVar2S372: std_logic_vector(   0 downto 0);
        signal oVar2S373: std_logic_vector(   0 downto 0);
        signal oVar2S374: std_logic_vector(   0 downto 0);
        signal oVar3S0: std_logic_vector(   0 downto 0);
        signal oVar3S1: std_logic_vector(   0 downto 0);
        signal oVar3S2: std_logic_vector(   0 downto 0);
        signal oVar3S3: std_logic_vector(   0 downto 0);
        signal oVar3S4: std_logic_vector(   0 downto 0);
        signal oVar3S5: std_logic_vector(   0 downto 0);
        signal oVar3S6: std_logic_vector(   0 downto 0);
        signal oVar3S7: std_logic_vector(   0 downto 0);
        signal oVar3S8: std_logic_vector(   0 downto 0);
        signal oVar3S9: std_logic_vector(   0 downto 0);
        signal oVar3S10: std_logic_vector(   0 downto 0);
        signal oVar3S11: std_logic_vector(   0 downto 0);
        signal oVar3S12: std_logic_vector(   0 downto 0);
        signal oVar3S13: std_logic_vector(   0 downto 0);
        signal oVar3S14: std_logic_vector(   0 downto 0);
        signal oVar3S15: std_logic_vector(   0 downto 0);
        signal oVar3S16: std_logic_vector(   0 downto 0);
        signal oVar3S17: std_logic_vector(   0 downto 0);
        signal oVar3S18: std_logic_vector(   0 downto 0);
        signal oVar3S19: std_logic_vector(   0 downto 0);
        signal oVar3S20: std_logic_vector(   0 downto 0);
        signal oVar3S21: std_logic_vector(   0 downto 0);
        signal oVar3S22: std_logic_vector(   0 downto 0);
        signal oVar3S23: std_logic_vector(   0 downto 0);
        signal oVar3S24: std_logic_vector(   0 downto 0);
        signal oVar3S25: std_logic_vector(   0 downto 0);
        signal oVar3S26: std_logic_vector(   0 downto 0);
        signal oVar3S27: std_logic_vector(   0 downto 0);
        signal oVar3S28: std_logic_vector(   0 downto 0);
        signal oVar3S29: std_logic_vector(   0 downto 0);
        signal oVar3S30: std_logic_vector(   0 downto 0);
        signal oVar3S31: std_logic_vector(   0 downto 0);
        signal oVar3S33: std_logic_vector(   0 downto 0);
        signal oVar3S34: std_logic_vector(   0 downto 0);
        signal oVar3S35: std_logic_vector(   0 downto 0);
        signal oVar3S37: std_logic_vector(   0 downto 0);
        signal oVar3S38: std_logic_vector(   0 downto 0);
        signal oVar3S39: std_logic_vector(   0 downto 0);
        signal oVar3S40: std_logic_vector(   0 downto 0);
        signal oVar3S41: std_logic_vector(   0 downto 0);
        signal oVar3S42: std_logic_vector(   0 downto 0);
        signal oVar3S43: std_logic_vector(   0 downto 0);
        signal oVar3S44: std_logic_vector(   0 downto 0);
        signal oVar3S45: std_logic_vector(   0 downto 0);
        signal oVar3S46: std_logic_vector(   0 downto 0);
        signal oVar3S47: std_logic_vector(   0 downto 0);
        signal oVar3S48: std_logic_vector(   0 downto 0);
        signal oVar3S49: std_logic_vector(   0 downto 0);
        signal oVar3S50: std_logic_vector(   0 downto 0);
        signal oVar3S51: std_logic_vector(   0 downto 0);
        signal oVar3S52: std_logic_vector(   0 downto 0);
        signal oVar3S53: std_logic_vector(   0 downto 0);
        signal oVar3S54: std_logic_vector(   0 downto 0);
        signal oVar3S55: std_logic_vector(   0 downto 0);
        signal oVar3S56: std_logic_vector(   0 downto 0);
        signal oVar3S57: std_logic_vector(   0 downto 0);
        signal oVar3S58: std_logic_vector(   0 downto 0);
        signal oVar3S59: std_logic_vector(   0 downto 0);
        signal oVar3S60: std_logic_vector(   0 downto 0);
        signal oVar3S61: std_logic_vector(   0 downto 0);
        signal oVar3S62: std_logic_vector(   0 downto 0);
        signal oVar3S63: std_logic_vector(   0 downto 0);
        signal oVar3S64: std_logic_vector(   0 downto 0);
        signal oVar3S65: std_logic_vector(   0 downto 0);
        signal oVar3S66: std_logic_vector(   0 downto 0);
        signal oVar3S67: std_logic_vector(   0 downto 0);
        signal oVar3S68: std_logic_vector(   0 downto 0);
        signal oVar3S69: std_logic_vector(   0 downto 0);
        signal oVar3S70: std_logic_vector(   0 downto 0);
        signal oVar3S71: std_logic_vector(   0 downto 0);
        signal oVar3S73: std_logic_vector(   0 downto 0);
        signal oVar3S74: std_logic_vector(   0 downto 0);
        signal oVar3S75: std_logic_vector(   0 downto 0);
        signal oVar3S76: std_logic_vector(   0 downto 0);
        signal oVar3S77: std_logic_vector(   0 downto 0);
        signal oVar3S78: std_logic_vector(   0 downto 0);
        signal oVar3S79: std_logic_vector(   0 downto 0);
        signal oVar3S80: std_logic_vector(   0 downto 0);
        signal oVar3S81: std_logic_vector(   0 downto 0);
        signal oVar3S82: std_logic_vector(   0 downto 0);
        signal oVar3S83: std_logic_vector(   0 downto 0);
        signal oVar3S84: std_logic_vector(   0 downto 0);
        signal oVar3S85: std_logic_vector(   0 downto 0);
        signal oVar3S86: std_logic_vector(   0 downto 0);
        signal oVar3S87: std_logic_vector(   0 downto 0);
        signal oVar3S88: std_logic_vector(   0 downto 0);
        signal oVar3S89: std_logic_vector(   0 downto 0);
        signal oVar3S90: std_logic_vector(   0 downto 0);
        signal oVar3S91: std_logic_vector(   0 downto 0);
        signal oVar3S92: std_logic_vector(   0 downto 0);
        signal oVar3S93: std_logic_vector(   0 downto 0);
        signal oVar3S94: std_logic_vector(   0 downto 0);
        signal oVar3S95: std_logic_vector(   0 downto 0);
        signal oVar3S96: std_logic_vector(   0 downto 0);
        signal oVar3S97: std_logic_vector(   0 downto 0);
        signal oVar3S98: std_logic_vector(   0 downto 0);
        signal oVar3S99: std_logic_vector(   0 downto 0);
        signal oVar3S100: std_logic_vector(   0 downto 0);
        signal oVar3S101: std_logic_vector(   0 downto 0);
        signal oVar3S102: std_logic_vector(   0 downto 0);
        signal oVar3S103: std_logic_vector(   0 downto 0);
        signal oVar3S104: std_logic_vector(   0 downto 0);
        signal oVar3S105: std_logic_vector(   0 downto 0);
        signal oVar3S106: std_logic_vector(   0 downto 0);
        signal oVar3S107: std_logic_vector(   0 downto 0);
        signal oVar3S108: std_logic_vector(   0 downto 0);
        signal oVar3S109: std_logic_vector(   0 downto 0);
        signal oVar3S110: std_logic_vector(   0 downto 0);
        signal oVar3S111: std_logic_vector(   0 downto 0);
        signal oVar3S112: std_logic_vector(   0 downto 0);
        signal oVar3S113: std_logic_vector(   0 downto 0);
        signal oVar3S114: std_logic_vector(   0 downto 0);
        signal oVar3S115: std_logic_vector(   0 downto 0);
        signal oVar3S116: std_logic_vector(   0 downto 0);
        signal oVar3S118: std_logic_vector(   0 downto 0);
        signal oVar3S119: std_logic_vector(   0 downto 0);
        signal oVar3S120: std_logic_vector(   0 downto 0);
        signal oVar3S121: std_logic_vector(   0 downto 0);
        signal oVar3S122: std_logic_vector(   0 downto 0);
        signal oVar3S123: std_logic_vector(   0 downto 0);
        signal oVar3S124: std_logic_vector(   0 downto 0);
        signal oVar3S125: std_logic_vector(   0 downto 0);
        signal oVar3S126: std_logic_vector(   0 downto 0);
        signal oVar3S127: std_logic_vector(   0 downto 0);
        signal oVar3S129: std_logic_vector(   0 downto 0);
        signal oVar3S130: std_logic_vector(   0 downto 0);
        signal oVar3S131: std_logic_vector(   0 downto 0);
        signal oVar3S132: std_logic_vector(   0 downto 0);
        signal aVar3S0: std_logic_vector(   15 downto 0);
        signal aVar3S1: std_logic_vector(   15 downto 0);
        signal aVar3S2: std_logic_vector(   15 downto 0);
        signal aVar3S3: std_logic_vector(   15 downto 0);
        signal aVar3S4: std_logic_vector(   15 downto 0);
        signal aVar3S5: std_logic_vector(   15 downto 0);
        signal aVar3S6: std_logic_vector(   15 downto 0);
        signal aVar3S7: std_logic_vector(   15 downto 0);
        signal aVar3S8: std_logic_vector(   15 downto 0);
        signal aVar3S9: std_logic_vector(   15 downto 0);
        signal aVar3S10: std_logic_vector(   15 downto 0);
        signal aVar3S11: std_logic_vector(   15 downto 0);
        signal aVar3S12: std_logic_vector(   15 downto 0);
        signal aVar3S13: std_logic_vector(   15 downto 0);
        signal aVar3S14: std_logic_vector(   15 downto 0);
        signal aVar3S15: std_logic_vector(   15 downto 0);
        signal aVar4S0: std_logic_vector(   15 downto 0);
        signal aVar4S1: std_logic_vector(   15 downto 0);
        signal aVar4S2: std_logic_vector(   15 downto 0);
        signal aVar4S3: std_logic_vector(   15 downto 0);
        signal aVar4S4: std_logic_vector(   15 downto 0);
        signal aVar4S5: std_logic_vector(   15 downto 0);
        signal aVar4S6: std_logic_vector(   15 downto 0);
        signal aVar4S7: std_logic_vector(   15 downto 0);
        signal aVar5S0: std_logic_vector(   15 downto 0);
        signal aVar5S1: std_logic_vector(   15 downto 0);
        signal aVar5S2: std_logic_vector(   15 downto 0);
        signal aVar5S3: std_logic_vector(   15 downto 0);
        signal aVar6S0: std_logic_vector(   15 downto 0);
        signal aVar6S1: std_logic_vector(   15 downto 0);
        signal aVar7S0: std_logic_vector(   15 downto 0);
signal ADDM4K3S1: std_logic_vector(   7 downto 0);
signal ADDM4K3S0: std_logic_vector(   7 downto 0);
signal ADDM4K3S3: std_logic_vector(   7 downto 0);
signal ADDM4K3S2: std_logic_vector(   7 downto 0);
signal ADDM4K3S5: std_logic_vector(   7 downto 0);
signal ADDM4K3S4: std_logic_vector(   7 downto 0);
signal ADDM4K3S7: std_logic_vector(   7 downto 0);
signal ADDM4K3S6: std_logic_vector(   7 downto 0);
signal ADDM4K3S9: std_logic_vector(   7 downto 0);
signal ADDM4K3S8: std_logic_vector(   7 downto 0);
signal ADDM4K3S11: std_logic_vector(   7 downto 0);
signal ADDM4K3S10: std_logic_vector(   7 downto 0);
signal ADDM4K3S13: std_logic_vector(   7 downto 0);
signal ADDM4K3S12: std_logic_vector(   7 downto 0);
signal ADDM4K3S15: std_logic_vector(   7 downto 0);
signal ADDM4K3S14: std_logic_vector(   7 downto 0);
BEGIN
	A (19 downto 0) <= A_DIN_L (19 downto 0);
	B (8 downto 0) <= A_DIN_L (28 downto 20);
	B (17 downto 9) <= B_DIN_L (8 downto 0);
	D (15 downto 0) <= B_DIN_L (24 downto 9);
	E (15 downto 0) <= D_DIN_L (31 downto 16);
	C_DOUT_L (31 downto 0) <= output (31 downto 0);
	F_DOUT_L (31 downto 0) <=  output (31 downto 0);
lookuptable_LV1 : process(c1)
begin
 if c1'event and c1='1' then
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='1' )then
          cVar1S0S0P069P019P067P064(0) <='1';
          else
          cVar1S0S0P069P019P067P064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='1' )then
          cVar1S1S0P069P019P067P064(0) <='1';
          else
          cVar1S1S0P069P019P067P064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='1' )then
          cVar1S2S0P069P019P067P064(0) <='1';
          else
          cVar1S2S0P069P019P067P064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='0' )then
          cVar1S3S0P069P019P067N064(0) <='1';
          else
          cVar1S3S0P069P019P067N064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='0' )then
          cVar1S4S0P069P019P067N064(0) <='1';
          else
          cVar1S4S0P069P019P067N064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='0' )then
          cVar1S5S0P069P019P067N064(0) <='1';
          else
          cVar1S5S0P069P019P067N064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='1' AND E( 1)='0' )then
          cVar1S6S0P069P019P067N064(0) <='1';
          else
          cVar1S6S0P069P019P067N064(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='0' AND D( 9)='1' )then
          cVar1S7S0P069P019N067P063(0) <='1';
          else
          cVar1S7S0P069P019N067P063(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='1' AND D( 8)='0' AND D( 9)='1' )then
          cVar1S8S0P069P019N067P063(0) <='1';
          else
          cVar1S8S0P069P019N067P063(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='1' )then
          cVar1S9S0P069N019P036P017(0) <='1';
          else
          cVar1S9S0P069N019P036P017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='1' )then
          cVar1S10S0P069N019P036P017(0) <='1';
          else
          cVar1S10S0P069N019P036P017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='1' )then
          cVar1S11S0P069N019P036P017(0) <='1';
          else
          cVar1S11S0P069N019P036P017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='0' )then
          cVar1S12S0P069N019P036N017(0) <='1';
          else
          cVar1S12S0P069N019P036N017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='0' )then
          cVar1S13S0P069N019P036N017(0) <='1';
          else
          cVar1S13S0P069N019P036N017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='1' AND A( 1)='0' )then
          cVar1S14S0P069N019P036N017(0) <='1';
          else
          cVar1S14S0P069N019P036N017(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='0' AND A(10)='1' )then
          cVar1S15S0P069N019N036P018(0) <='1';
          else
          cVar1S15S0P069N019N036P018(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='0' AND A(10)='1' )then
          cVar1S16S0P069N019N036P018(0) <='1';
          else
          cVar1S16S0P069N019N036P018(0) <='0';
          end if;
        if(E( 8)='1' AND A( 0)='0' AND B( 9)='0' AND A(10)='0' )then
          cVar1S17S0P069N019N036N018(0) <='1';
          else
          cVar1S17S0P069N019N036N018(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S18S0N069P063P065P017(0) <='1';
          else
          cVar1S18S0N069P063P065P017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S19S0N069P063P065P017(0) <='1';
          else
          cVar1S19S0N069P063P065P017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S20S0N069P063P065P017(0) <='1';
          else
          cVar1S20S0N069P063P065P017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S21S0N069P063P065P017(0) <='1';
          else
          cVar1S21S0N069P063P065P017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S22S0N069P063P065N017(0) <='1';
          else
          cVar1S22S0N069P063P065N017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S23S0N069P063P065N017(0) <='1';
          else
          cVar1S23S0N069P063P065N017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S24S0N069P063P065N017(0) <='1';
          else
          cVar1S24S0N069P063P065N017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S25S0N069P063P065N017(0) <='1';
          else
          cVar1S25S0N069P063P065N017(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='0' AND E(10)='1' )then
          cVar1S26S0N069P063N065P061(0) <='1';
          else
          cVar1S26S0N069P063N065P061(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='1' AND E( 9)='0' AND E(10)='1' )then
          cVar1S27S0N069P063N065P061(0) <='1';
          else
          cVar1S27S0N069P063N065P061(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='1' AND D(10)='1' )then
          cVar1S28S0N069N063P061P059(0) <='1';
          else
          cVar1S28S0N069N063P061P059(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='1' AND D(10)='1' )then
          cVar1S29S0N069N063P061P059(0) <='1';
          else
          cVar1S29S0N069N063P061P059(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='1' AND D(10)='1' )then
          cVar1S30S0N069N063P061P059(0) <='1';
          else
          cVar1S30S0N069N063P061P059(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='1' AND D(10)='1' )then
          cVar1S31S0N069N063P061P059(0) <='1';
          else
          cVar1S31S0N069N063P061P059(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='1' )then
          cVar1S32S0N069N063N061P055(0) <='1';
          else
          cVar1S32S0N069N063N061P055(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='1' )then
          cVar1S33S0N069N063N061P055(0) <='1';
          else
          cVar1S33S0N069N063N061P055(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='1' )then
          cVar1S34S0N069N063N061P055(0) <='1';
          else
          cVar1S34S0N069N063N061P055(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='1' )then
          cVar1S35S0N069N063N061P055(0) <='1';
          else
          cVar1S35S0N069N063N061P055(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='0' )then
          cVar1S36S0N069N063N061N055(0) <='1';
          else
          cVar1S36S0N069N063N061N055(0) <='0';
          end if;
        if(E( 8)='0' AND D( 9)='0' AND E(10)='0' AND D(11)='0' )then
          cVar1S37S0N069N063N061N055(0) <='1';
          else
          cVar1S37S0N069N063N061N055(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='1' AND E( 0)='0' )then
          cVar1S0S1P052P050P010P068(0) <='1';
          else
          cVar1S0S1P052P050P010P068(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='1' AND E( 0)='0' )then
          cVar1S1S1P052P050P010P068(0) <='1';
          else
          cVar1S1S1P052P050P010P068(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='1' AND E( 0)='1' )then
          cVar1S2S1P052P050P010P068(0) <='1';
          else
          cVar1S2S1P052P050P010P068(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='1' AND E( 0)='1' )then
          cVar1S3S1P052P050P010P068(0) <='1';
          else
          cVar1S3S1P052P050P010P068(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar1S4S1P052P050N010P069(0) <='1';
          else
          cVar1S4S1P052P050N010P069(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar1S5S1P052P050N010P069(0) <='1';
          else
          cVar1S5S1P052P050N010P069(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='0' AND E( 8)='0' )then
          cVar1S6S1P052P050N010N069(0) <='1';
          else
          cVar1S6S1P052P050N010N069(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='1' AND A(14)='0' AND E( 8)='0' )then
          cVar1S7S1P052P050N010N069(0) <='1';
          else
          cVar1S7S1P052P050N010N069(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='0' AND B( 4)='1' )then
          cVar1S8S1P052N050P029nsss(0) <='1';
          else
          cVar1S8S1P052N050P029nsss(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='0' AND B( 4)='0' AND B(13)='1' )then
          cVar1S9S1P052N050N029P028(0) <='1';
          else
          cVar1S9S1P052N050N029P028(0) <='0';
          end if;
        if(E( 4)='1' AND D( 4)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S10S1P052N050N029N028(0) <='1';
          else
          cVar1S10S1P052N050N029N028(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='1' AND D( 9)='1' )then
          cVar1S11S1N052P056P031P063(0) <='1';
          else
          cVar1S11S1N052P056P031P063(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='1' AND D( 9)='1' )then
          cVar1S12S1N052P056P031P063(0) <='1';
          else
          cVar1S12S1N052P056P031P063(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='1' AND D( 9)='0' )then
          cVar1S13S1N052P056P031N063psss(0) <='1';
          else
          cVar1S13S1N052P056P031N063psss(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='0' AND B( 4)='1' )then
          cVar1S14S1N052P056N031P029(0) <='1';
          else
          cVar1S14S1N052P056N031P029(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='0' AND B( 4)='0' )then
          cVar1S15S1N052P056N031N029(0) <='1';
          else
          cVar1S15S1N052P056N031N029(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='0' AND B( 4)='0' )then
          cVar1S16S1N052P056N031N029(0) <='1';
          else
          cVar1S16S1N052P056N031N029(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='0' AND B( 4)='0' )then
          cVar1S17S1N052P056N031N029(0) <='1';
          else
          cVar1S17S1N052P056N031N029(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='1' AND B( 3)='0' AND B( 4)='0' )then
          cVar1S18S1N052P056N031N029(0) <='1';
          else
          cVar1S18S1N052P056N031N029(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='0' )then
          cVar1S19S1N052N056P060P065(0) <='1';
          else
          cVar1S19S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='0' )then
          cVar1S20S1N052N056P060P065(0) <='1';
          else
          cVar1S20S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='0' )then
          cVar1S21S1N052N056P060P065(0) <='1';
          else
          cVar1S21S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='0' )then
          cVar1S22S1N052N056P060P065(0) <='1';
          else
          cVar1S22S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='1' )then
          cVar1S23S1N052N056P060P065(0) <='1';
          else
          cVar1S23S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='1' )then
          cVar1S24S1N052N056P060P065(0) <='1';
          else
          cVar1S24S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='1' AND E( 9)='1' )then
          cVar1S25S1N052N056P060P065(0) <='1';
          else
          cVar1S25S1N052N056P060P065(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='1' )then
          cVar1S26S1N052N056N060P046(0) <='1';
          else
          cVar1S26S1N052N056N060P046(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='1' )then
          cVar1S27S1N052N056N060P046(0) <='1';
          else
          cVar1S27S1N052N056N060P046(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='1' )then
          cVar1S28S1N052N056N060P046(0) <='1';
          else
          cVar1S28S1N052N056N060P046(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='0' )then
          cVar1S29S1N052N056N060N046(0) <='1';
          else
          cVar1S29S1N052N056N060N046(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='0' )then
          cVar1S30S1N052N056N060N046(0) <='1';
          else
          cVar1S30S1N052N056N060N046(0) <='0';
          end if;
        if(E( 4)='0' AND E( 3)='0' AND E( 2)='0' AND D( 5)='0' )then
          cVar1S31S1N052N056N060N046(0) <='1';
          else
          cVar1S31S1N052N056N060N046(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='0' )then
          cVar1S0S2P068P067P066P035(0) <='1';
          else
          cVar1S0S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='0' )then
          cVar1S1S2P068P067P066P035(0) <='1';
          else
          cVar1S1S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='0' )then
          cVar1S2S2P068P067P066P035(0) <='1';
          else
          cVar1S2S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='0' )then
          cVar1S3S2P068P067P066P035(0) <='1';
          else
          cVar1S3S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='1' )then
          cVar1S4S2P068P067P066P035(0) <='1';
          else
          cVar1S4S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='1' )then
          cVar1S5S2P068P067P066P035(0) <='1';
          else
          cVar1S5S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='1' AND B( 1)='1' )then
          cVar1S6S2P068P067P066P035(0) <='1';
          else
          cVar1S6S2P068P067P066P035(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='0' AND D( 9)='1' )then
          cVar1S7S2P068P067N066P063(0) <='1';
          else
          cVar1S7S2P068P067N066P063(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='0' AND D( 9)='1' )then
          cVar1S8S2P068P067N066P063(0) <='1';
          else
          cVar1S8S2P068P067N066P063(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S9S2P068P067N066N063(0) <='1';
          else
          cVar1S9S2P068P067N066N063(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S10S2P068P067N066N063(0) <='1';
          else
          cVar1S10S2P068P067N066N063(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='1' )then
          cVar1S11S2P068P067P035P016(0) <='1';
          else
          cVar1S11S2P068P067P035P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='1' )then
          cVar1S12S2P068P067P035P016(0) <='1';
          else
          cVar1S12S2P068P067P035P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='1' )then
          cVar1S13S2P068P067P035P016(0) <='1';
          else
          cVar1S13S2P068P067P035P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='0' )then
          cVar1S14S2P068P067P035N016(0) <='1';
          else
          cVar1S14S2P068P067P035N016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='0' )then
          cVar1S15S2P068P067P035N016(0) <='1';
          else
          cVar1S15S2P068P067P035N016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='0' AND A(11)='0' )then
          cVar1S16S2P068P067P035N016(0) <='1';
          else
          cVar1S16S2P068P067P035N016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='1' AND B( 3)='1' )then
          cVar1S17S2P068P067P035P031nsss(0) <='1';
          else
          cVar1S17S2P068P067P035P031nsss(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND B( 1)='1' AND B( 3)='0' )then
          cVar1S18S2P068P067P035N031(0) <='1';
          else
          cVar1S18S2P068P067P035N031(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='0' AND E( 9)='1' )then
          cVar1S19S2N068P063P062P065(0) <='1';
          else
          cVar1S19S2N068P063P062P065(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='0' AND E( 9)='1' )then
          cVar1S20S2N068P063P062P065(0) <='1';
          else
          cVar1S20S2N068P063P062P065(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='0' AND E( 9)='1' )then
          cVar1S21S2N068P063P062P065(0) <='1';
          else
          cVar1S21S2N068P063P062P065(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='0' AND E( 9)='0' )then
          cVar1S22S2N068P063P062N065(0) <='1';
          else
          cVar1S22S2N068P063P062N065(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='0' AND E( 9)='0' )then
          cVar1S23S2N068P063P062N065(0) <='1';
          else
          cVar1S23S2N068P063P062N065(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='1' AND B( 1)='0' )then
          cVar1S24S2N068P063P062P035(0) <='1';
          else
          cVar1S24S2N068P063P062P035(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='1' AND B( 1)='1' )then
          cVar1S25S2N068P063P062P035(0) <='1';
          else
          cVar1S25S2N068P063P062P035(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='1' AND B( 1)='1' )then
          cVar1S26S2N068P063P062P035(0) <='1';
          else
          cVar1S26S2N068P063P062P035(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='1' AND B( 1)='1' )then
          cVar1S27S2N068P063P062P035(0) <='1';
          else
          cVar1S27S2N068P063P062P035(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='1' AND D( 1)='1' AND B( 1)='1' )then
          cVar1S28S2N068P063P062P035(0) <='1';
          else
          cVar1S28S2N068P063P062P035(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='1' AND B(13)='1' )then
          cVar1S29S2N068N063P051P028nsss(0) <='1';
          else
          cVar1S29S2N068N063P051P028nsss(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='1' AND B(13)='0' )then
          cVar1S30S2N068N063P051N028(0) <='1';
          else
          cVar1S30S2N068N063P051N028(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='1' AND B(13)='0' )then
          cVar1S31S2N068N063P051N028(0) <='1';
          else
          cVar1S31S2N068N063P051N028(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='1' AND B(13)='0' )then
          cVar1S32S2N068N063P051N028(0) <='1';
          else
          cVar1S32S2N068N063P051N028(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='1' )then
          cVar1S33S2N068N063N051P067(0) <='1';
          else
          cVar1S33S2N068N063N051P067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='1' )then
          cVar1S34S2N068N063N051P067(0) <='1';
          else
          cVar1S34S2N068N063N051P067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='1' )then
          cVar1S35S2N068N063N051P067(0) <='1';
          else
          cVar1S35S2N068N063N051P067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='1' )then
          cVar1S36S2N068N063N051P067(0) <='1';
          else
          cVar1S36S2N068N063N051P067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='0' )then
          cVar1S37S2N068N063N051N067(0) <='1';
          else
          cVar1S37S2N068N063N051N067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='0' )then
          cVar1S38S2N068N063N051N067(0) <='1';
          else
          cVar1S38S2N068N063N051N067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='0' )then
          cVar1S39S2N068N063N051N067(0) <='1';
          else
          cVar1S39S2N068N063N051N067(0) <='0';
          end if;
        if(E( 0)='0' AND D( 9)='0' AND D(12)='0' AND D( 8)='0' )then
          cVar1S40S2N068N063N051N067(0) <='1';
          else
          cVar1S40S2N068N063N051N067(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' )then
          cVar1S0S3P043P022nsss(0) <='1';
          else
          cVar1S0S3P043P022nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='1' AND A( 2)='0' )then
          cVar1S1S3P043N022P007P015(0) <='1';
          else
          cVar1S1S3P043N022P007P015(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='1' AND A( 2)='0' )then
          cVar1S2S3P043N022P007P015(0) <='1';
          else
          cVar1S2S3P043N022P007P015(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='1' AND A( 2)='1' )then
          cVar1S3S3P043N022P007P015psss(0) <='1';
          else
          cVar1S3S3P043N022P007P015psss(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='0' AND E(13)='0' )then
          cVar1S4S3P043N022N007P049(0) <='1';
          else
          cVar1S4S3P043N022N007P049(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='0' AND E(13)='0' )then
          cVar1S5S3P043N022N007P049(0) <='1';
          else
          cVar1S5S3P043N022N007P049(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND A( 6)='0' AND E(13)='0' )then
          cVar1S6S3P043N022N007P049(0) <='1';
          else
          cVar1S6S3P043N022N007P049(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='0' AND E( 2)='0' )then
          cVar1S7S3N043P067P068P060(0) <='1';
          else
          cVar1S7S3N043P067P068P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='0' AND E( 2)='0' )then
          cVar1S8S3N043P067P068P060(0) <='1';
          else
          cVar1S8S3N043P067P068P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='0' AND E( 2)='0' )then
          cVar1S9S3N043P067P068P060(0) <='1';
          else
          cVar1S9S3N043P067P068P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='0' AND E( 2)='1' )then
          cVar1S10S3N043P067P068P060(0) <='1';
          else
          cVar1S10S3N043P067P068P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='1' AND A(11)='1' )then
          cVar1S11S3N043P067P068P016(0) <='1';
          else
          cVar1S11S3N043P067P068P016(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='1' AND A(11)='1' )then
          cVar1S12S3N043P067P068P016(0) <='1';
          else
          cVar1S12S3N043P067P068P016(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='1' AND A(11)='0' )then
          cVar1S13S3N043P067P068N016(0) <='1';
          else
          cVar1S13S3N043P067P068N016(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='1' AND A(11)='0' )then
          cVar1S14S3N043P067P068N016(0) <='1';
          else
          cVar1S14S3N043P067P068N016(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='1' AND E( 0)='1' AND A(11)='0' )then
          cVar1S15S3N043P067P068N016(0) <='1';
          else
          cVar1S15S3N043P067P068N016(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='0' )then
          cVar1S16S3N043N067P034P062(0) <='1';
          else
          cVar1S16S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='0' )then
          cVar1S17S3N043N067P034P062(0) <='1';
          else
          cVar1S17S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='0' )then
          cVar1S18S3N043N067P034P062(0) <='1';
          else
          cVar1S18S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='0' )then
          cVar1S19S3N043N067P034P062(0) <='1';
          else
          cVar1S19S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='1' )then
          cVar1S20S3N043N067P034P062(0) <='1';
          else
          cVar1S20S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='1' AND D( 1)='1' )then
          cVar1S21S3N043N067P034P062(0) <='1';
          else
          cVar1S21S3N043N067P034P062(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='1' )then
          cVar1S22S3N043N067N034P051(0) <='1';
          else
          cVar1S22S3N043N067N034P051(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='1' )then
          cVar1S23S3N043N067N034P051(0) <='1';
          else
          cVar1S23S3N043N067N034P051(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='1' )then
          cVar1S24S3N043N067N034P051(0) <='1';
          else
          cVar1S24S3N043N067N034P051(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='0' )then
          cVar1S25S3N043N067N034N051(0) <='1';
          else
          cVar1S25S3N043N067N034N051(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='0' )then
          cVar1S26S3N043N067N034N051(0) <='1';
          else
          cVar1S26S3N043N067N034N051(0) <='0';
          end if;
        if(D(14)='0' AND D( 8)='0' AND B(10)='0' AND D(12)='0' )then
          cVar1S27S3N043N067N034N051(0) <='1';
          else
          cVar1S27S3N043N067N034N051(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='1' AND A(16)='1' )then
          cVar1S0S4P044P023P006nsss(0) <='1';
          else
          cVar1S0S4P044P023P006nsss(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='1' AND A(16)='0' AND A(17)='1' )then
          cVar1S1S4P044P023N006P004nsss(0) <='1';
          else
          cVar1S1S4P044P023N006P004nsss(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='1' AND A(16)='0' AND A(17)='0' )then
          cVar1S2S4P044P023N006N004(0) <='1';
          else
          cVar1S2S4P044P023N006N004(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='1' AND A(10)='0' )then
          cVar1S3S4P044N023P025P018(0) <='1';
          else
          cVar1S3S4P044N023P025P018(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='1' AND A(10)='0' )then
          cVar1S4S4P044N023P025P018(0) <='1';
          else
          cVar1S4S4P044N023P025P018(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='1' AND A(10)='1' )then
          cVar1S5S4P044N023P025P018psss(0) <='1';
          else
          cVar1S5S4P044N023P025P018psss(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='0' AND B(16)='1' )then
          cVar1S6S4P044N023N025P022(0) <='1';
          else
          cVar1S6S4P044N023N025P022(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='0' AND B(16)='0' )then
          cVar1S7S4P044N023N025N022(0) <='1';
          else
          cVar1S7S4P044N023N025N022(0) <='0';
          end if;
        if(E( 6)='1' AND B( 7)='0' AND B( 6)='0' AND B(16)='0' )then
          cVar1S8S4P044N023N025N022(0) <='1';
          else
          cVar1S8S4P044N023N025N022(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='0' AND D( 8)='0' )then
          cVar1S9S4N044P037P008P067(0) <='1';
          else
          cVar1S9S4N044P037P008P067(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='0' AND D( 8)='0' )then
          cVar1S10S4N044P037P008P067(0) <='1';
          else
          cVar1S10S4N044P037P008P067(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='0' AND D( 8)='0' )then
          cVar1S11S4N044P037P008P067(0) <='1';
          else
          cVar1S11S4N044P037P008P067(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='0' AND D( 8)='1' )then
          cVar1S12S4N044P037P008P067(0) <='1';
          else
          cVar1S12S4N044P037P008P067(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='0' AND D( 8)='1' )then
          cVar1S13S4N044P037P008P067(0) <='1';
          else
          cVar1S13S4N044P037P008P067(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='1' AND D( 4)='1' )then
          cVar1S14S4N044P037P008P050(0) <='1';
          else
          cVar1S14S4N044P037P008P050(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='1' AND D( 4)='0' )then
          cVar1S15S4N044P037P008N050(0) <='1';
          else
          cVar1S15S4N044P037P008N050(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='1' AND A(15)='1' AND D( 4)='0' )then
          cVar1S16S4N044P037P008N050(0) <='1';
          else
          cVar1S16S4N044P037P008N050(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='1' AND D( 0)='0' )then
          cVar1S17S4N044N037P031P066(0) <='1';
          else
          cVar1S17S4N044N037P031P066(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='1' AND D( 0)='0' )then
          cVar1S18S4N044N037P031P066(0) <='1';
          else
          cVar1S18S4N044N037P031P066(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='1' AND D( 0)='0' )then
          cVar1S19S4N044N037P031P066(0) <='1';
          else
          cVar1S19S4N044N037P031P066(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='1' AND D( 0)='0' )then
          cVar1S20S4N044N037P031P066(0) <='1';
          else
          cVar1S20S4N044N037P031P066(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='1' AND D( 0)='1' )then
          cVar1S21S4N044N037P031P066(0) <='1';
          else
          cVar1S21S4N044N037P031P066(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='1' )then
          cVar1S22S4N044N037N031P036(0) <='1';
          else
          cVar1S22S4N044N037N031P036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='1' )then
          cVar1S23S4N044N037N031P036(0) <='1';
          else
          cVar1S23S4N044N037N031P036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='1' )then
          cVar1S24S4N044N037N031P036(0) <='1';
          else
          cVar1S24S4N044N037N031P036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='1' )then
          cVar1S25S4N044N037N031P036(0) <='1';
          else
          cVar1S25S4N044N037N031P036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='0' )then
          cVar1S26S4N044N037N031N036(0) <='1';
          else
          cVar1S26S4N044N037N031N036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='0' )then
          cVar1S27S4N044N037N031N036(0) <='1';
          else
          cVar1S27S4N044N037N031N036(0) <='0';
          end if;
        if(E( 6)='0' AND B( 0)='0' AND B( 3)='0' AND B( 9)='0' )then
          cVar1S28S4N044N037N031N036(0) <='1';
          else
          cVar1S28S4N044N037N031N036(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='1' AND E( 4)='0' AND D( 4)='1' )then
          cVar1S0S5P027P048P052P050nsss(0) <='1';
          else
          cVar1S0S5P027P048P052P050nsss(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='1' AND E( 4)='0' AND D( 4)='0' )then
          cVar1S1S5P027P048P052N050(0) <='1';
          else
          cVar1S1S5P027P048P052N050(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='1' AND E( 4)='0' AND D( 4)='0' )then
          cVar1S2S5P027P048P052N050(0) <='1';
          else
          cVar1S2S5P027P048P052N050(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='1' AND E( 4)='0' AND D( 4)='0' )then
          cVar1S3S5P027P048P052N050(0) <='1';
          else
          cVar1S3S5P027P048P052N050(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S4S5P027P048P052P009nsss(0) <='1';
          else
          cVar1S4S5P027P048P052P009nsss(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='1' AND A(15)='1' )then
          cVar1S5S5P027N048P050P008nsss(0) <='1';
          else
          cVar1S5S5P027N048P050P008nsss(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S6S5P027N048P050N008(0) <='1';
          else
          cVar1S6S5P027N048P050N008(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S7S5P027N048P050N008(0) <='1';
          else
          cVar1S7S5P027N048P050N008(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S8S5P027N048P050N008(0) <='1';
          else
          cVar1S8S5P027N048P050N008(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='0' AND E(13)='1' )then
          cVar1S9S5P027N048N050P049(0) <='1';
          else
          cVar1S9S5P027N048N050P049(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='0' AND E(13)='0' )then
          cVar1S10S5P027N048N050N049(0) <='1';
          else
          cVar1S10S5P027N048N050N049(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='0' AND E(13)='0' )then
          cVar1S11S5P027N048N050N049(0) <='1';
          else
          cVar1S11S5P027N048N050N049(0) <='0';
          end if;
        if(B( 5)='1' AND E( 5)='0' AND D( 4)='0' AND E(13)='0' )then
          cVar1S12S5P027N048N050N049(0) <='1';
          else
          cVar1S12S5P027N048N050N049(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='1' )then
          cVar1S13S5N027P043P022nsss(0) <='1';
          else
          cVar1S13S5N027P043P022nsss(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='0' AND A( 6)='1' )then
          cVar1S14S5N027P043N022P007(0) <='1';
          else
          cVar1S14S5N027P043N022P007(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='0' AND A( 6)='0' )then
          cVar1S15S5N027P043N022N007(0) <='1';
          else
          cVar1S15S5N027P043N022N007(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='0' AND A( 6)='0' )then
          cVar1S16S5N027P043N022N007(0) <='1';
          else
          cVar1S16S5N027P043N022N007(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='0' AND A( 6)='0' )then
          cVar1S17S5N027P043N022N007(0) <='1';
          else
          cVar1S17S5N027P043N022N007(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='1' AND B(16)='0' AND A( 6)='0' )then
          cVar1S18S5N027P043N022N007(0) <='1';
          else
          cVar1S18S5N027P043N022N007(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='0' )then
          cVar1S19S5N027N043P036P015(0) <='1';
          else
          cVar1S19S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='0' )then
          cVar1S20S5N027N043P036P015(0) <='1';
          else
          cVar1S20S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='0' )then
          cVar1S21S5N027N043P036P015(0) <='1';
          else
          cVar1S21S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='0' )then
          cVar1S22S5N027N043P036P015(0) <='1';
          else
          cVar1S22S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='1' )then
          cVar1S23S5N027N043P036P015(0) <='1';
          else
          cVar1S23S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='1' )then
          cVar1S24S5N027N043P036P015(0) <='1';
          else
          cVar1S24S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='1' AND A( 2)='1' )then
          cVar1S25S5N027N043P036P015(0) <='1';
          else
          cVar1S25S5N027N043P036P015(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='1' )then
          cVar1S26S5N027N043N036P068(0) <='1';
          else
          cVar1S26S5N027N043N036P068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='1' )then
          cVar1S27S5N027N043N036P068(0) <='1';
          else
          cVar1S27S5N027N043N036P068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='1' )then
          cVar1S28S5N027N043N036P068(0) <='1';
          else
          cVar1S28S5N027N043N036P068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='0' )then
          cVar1S29S5N027N043N036N068(0) <='1';
          else
          cVar1S29S5N027N043N036N068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='0' )then
          cVar1S30S5N027N043N036N068(0) <='1';
          else
          cVar1S30S5N027N043N036N068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='0' )then
          cVar1S31S5N027N043N036N068(0) <='1';
          else
          cVar1S31S5N027N043N036N068(0) <='0';
          end if;
        if(B( 5)='0' AND D(14)='0' AND B( 9)='0' AND E( 0)='0' )then
          cVar1S32S5N027N043N036N068(0) <='1';
          else
          cVar1S32S5N027N043N036N068(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='1' )then
          cVar1S0S6P040P021nsss(0) <='1';
          else
          cVar1S0S6P040P021nsss(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='1' AND A(10)='1' )then
          cVar1S1S6P040N021P023P018nsss(0) <='1';
          else
          cVar1S1S6P040N021P023P018nsss(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='1' AND A(10)='0' )then
          cVar1S2S6P040N021P023N018(0) <='1';
          else
          cVar1S2S6P040N021P023N018(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S3S6P040N021N023P020(0) <='1';
          else
          cVar1S3S6P040N021N023P020(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S4S6P040N021N023P020(0) <='1';
          else
          cVar1S4S6P040N021N023P020(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S5S6P040N021N023N020(0) <='1';
          else
          cVar1S5S6P040N021N023N020(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S6S6P040N021N023N020(0) <='1';
          else
          cVar1S6S6P040N021N023N020(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='1' AND A(11)='0' )then
          cVar1S7S6N040P025P046P016(0) <='1';
          else
          cVar1S7S6N040P025P046P016(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='1' AND A(11)='1' )then
          cVar1S8S6N040P025P046P016(0) <='1';
          else
          cVar1S8S6N040P025P046P016(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='0' AND E( 6)='1' )then
          cVar1S9S6N040P025N046P044nsss(0) <='1';
          else
          cVar1S9S6N040P025N046P044nsss(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='0' AND E( 6)='0' )then
          cVar1S10S6N040P025N046N044(0) <='1';
          else
          cVar1S10S6N040P025N046N044(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='0' AND E( 6)='0' )then
          cVar1S11S6N040P025N046N044(0) <='1';
          else
          cVar1S11S6N040P025N046N044(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='1' AND D( 5)='0' AND E( 6)='0' )then
          cVar1S12S6N040P025N046N044(0) <='1';
          else
          cVar1S12S6N040P025N046N044(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='0' )then
          cVar1S13S6N040N025P056P055(0) <='1';
          else
          cVar1S13S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='0' )then
          cVar1S14S6N040N025P056P055(0) <='1';
          else
          cVar1S14S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='0' )then
          cVar1S15S6N040N025P056P055(0) <='1';
          else
          cVar1S15S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='1' )then
          cVar1S16S6N040N025P056P055(0) <='1';
          else
          cVar1S16S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='1' )then
          cVar1S17S6N040N025P056P055(0) <='1';
          else
          cVar1S17S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='1' )then
          cVar1S18S6N040N025P056P055(0) <='1';
          else
          cVar1S18S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='1' AND D(11)='1' )then
          cVar1S19S6N040N025P056P055(0) <='1';
          else
          cVar1S19S6N040N025P056P055(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='1' )then
          cVar1S20S6N040N025N056P060(0) <='1';
          else
          cVar1S20S6N040N025N056P060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='1' )then
          cVar1S21S6N040N025N056P060(0) <='1';
          else
          cVar1S21S6N040N025N056P060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='1' )then
          cVar1S22S6N040N025N056P060(0) <='1';
          else
          cVar1S22S6N040N025N056P060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='0' )then
          cVar1S23S6N040N025N056N060(0) <='1';
          else
          cVar1S23S6N040N025N056N060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='0' )then
          cVar1S24S6N040N025N056N060(0) <='1';
          else
          cVar1S24S6N040N025N056N060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='0' )then
          cVar1S25S6N040N025N056N060(0) <='1';
          else
          cVar1S25S6N040N025N056N060(0) <='0';
          end if;
        if(E( 7)='0' AND B( 6)='0' AND E( 3)='0' AND E( 2)='0' )then
          cVar1S26S6N040N025N056N060(0) <='1';
          else
          cVar1S26S6N040N025N056N060(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='1' )then
          cVar1S0S7P066P028P055nsss(0) <='1';
          else
          cVar1S0S7P066P028P055nsss(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='0' AND E(12)='1' )then
          cVar1S1S7P066P028N055P053nsss(0) <='1';
          else
          cVar1S1S7P066P028N055P053nsss(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='0' AND E(12)='0' )then
          cVar1S2S7P066P028N055N053(0) <='1';
          else
          cVar1S2S7P066P028N055N053(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='0' AND E(12)='0' )then
          cVar1S3S7P066P028N055N053(0) <='1';
          else
          cVar1S3S7P066P028N055N053(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='0' AND E(12)='0' )then
          cVar1S4S7P066P028N055N053(0) <='1';
          else
          cVar1S4S7P066P028N055N053(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='1' AND D(11)='0' AND E(12)='0' )then
          cVar1S5S7P066P028N055N053(0) <='1';
          else
          cVar1S5S7P066P028N055N053(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='1' AND B( 7)='1' )then
          cVar1S6S7P066N028P044P023nsss(0) <='1';
          else
          cVar1S6S7P066N028P044P023nsss(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S7S7P066N028P044N023(0) <='1';
          else
          cVar1S7S7P066N028P044N023(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S8S7P066N028P044N023(0) <='1';
          else
          cVar1S8S7P066N028P044N023(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S9S7P066N028P044N023(0) <='1';
          else
          cVar1S9S7P066N028P044N023(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S10S7P066N028P044N023(0) <='1';
          else
          cVar1S10S7P066N028P044N023(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S11S7P066N028N044P040(0) <='1';
          else
          cVar1S11S7P066N028N044P040(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S12S7P066N028N044P040(0) <='1';
          else
          cVar1S12S7P066N028N044P040(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S13S7P066N028N044P040(0) <='1';
          else
          cVar1S13S7P066N028N044P040(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S14S7P066N028N044N040(0) <='1';
          else
          cVar1S14S7P066N028N044N040(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S15S7P066N028N044N040(0) <='1';
          else
          cVar1S15S7P066N028N044N040(0) <='0';
          end if;
        if(D( 0)='0' AND B(13)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S16S7P066N028N044N040(0) <='1';
          else
          cVar1S16S7P066N028N044N040(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='0' AND D( 8)='0' )then
          cVar1S17S7P066P065P003P067(0) <='1';
          else
          cVar1S17S7P066P065P003P067(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='0' AND D( 8)='0' )then
          cVar1S18S7P066P065P003P067(0) <='1';
          else
          cVar1S18S7P066P065P003P067(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='0' AND D( 8)='1' )then
          cVar1S19S7P066P065P003P067(0) <='1';
          else
          cVar1S19S7P066P065P003P067(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='0' AND D( 8)='1' )then
          cVar1S20S7P066P065P003P067(0) <='1';
          else
          cVar1S20S7P066P065P003P067(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='1' AND E(15)='1' )then
          cVar1S21S7P066P065P003P041nsss(0) <='1';
          else
          cVar1S21S7P066P065P003P041nsss(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='0' AND A( 8)='1' AND E(15)='0' )then
          cVar1S22S7P066P065P003N041(0) <='1';
          else
          cVar1S22S7P066P065P003N041(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='0' AND A(10)='1' )then
          cVar1S23S7P066P065P068P018(0) <='1';
          else
          cVar1S23S7P066P065P068P018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S24S7P066P065P068N018(0) <='1';
          else
          cVar1S24S7P066P065P068N018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S25S7P066P065P068N018(0) <='1';
          else
          cVar1S25S7P066P065P068N018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='1' AND A(10)='0' )then
          cVar1S26S7P066P065P068P018(0) <='1';
          else
          cVar1S26S7P066P065P068P018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='1' AND A(10)='0' )then
          cVar1S27S7P066P065P068P018(0) <='1';
          else
          cVar1S27S7P066P065P068P018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='1' AND A(10)='1' )then
          cVar1S28S7P066P065P068P018(0) <='1';
          else
          cVar1S28S7P066P065P068P018(0) <='0';
          end if;
        if(D( 0)='1' AND E( 9)='1' AND E( 0)='1' AND A(10)='1' )then
          cVar1S29S7P066P065P068P018(0) <='1';
          else
          cVar1S29S7P066P065P068P018(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='1' AND E( 1)='1' )then
          cVar1S0S8P043P045P064nsss(0) <='1';
          else
          cVar1S0S8P043P045P064nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='1' AND E( 1)='0' AND B( 3)='0' )then
          cVar1S1S8P043P045N064P031(0) <='1';
          else
          cVar1S1S8P043P045N064P031(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='1' AND E( 1)='0' AND B( 3)='0' )then
          cVar1S2S8P043P045N064P031(0) <='1';
          else
          cVar1S2S8P043P045N064P031(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='1' AND E( 1)='0' AND B( 3)='0' )then
          cVar1S3S8P043P045N064P031(0) <='1';
          else
          cVar1S3S8P043P045N064P031(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='0' AND A( 7)='1' AND B(16)='1' )then
          cVar1S4S8P043N045P005P022nsss(0) <='1';
          else
          cVar1S4S8P043N045P005P022nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='0' AND A( 7)='1' AND B(16)='0' )then
          cVar1S5S8P043N045P005N022(0) <='1';
          else
          cVar1S5S8P043N045P005N022(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='0' AND A( 7)='0' AND B(16)='1' )then
          cVar1S6S8P043N045N005P022(0) <='1';
          else
          cVar1S6S8P043N045N005P022(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='0' AND A( 7)='0' AND B(16)='0' )then
          cVar1S7S8P043N045N005N022(0) <='1';
          else
          cVar1S7S8P043N045N005N022(0) <='0';
          end if;
        if(D(14)='1' AND E(14)='0' AND A( 7)='0' AND B(16)='0' )then
          cVar1S8S8P043N045N005N022(0) <='1';
          else
          cVar1S8S8P043N045N005N022(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='1' AND B( 8)='1' )then
          cVar1S9S8N043P003P040P021nsss(0) <='1';
          else
          cVar1S9S8N043P003P040P021nsss(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='1' AND B( 8)='0' )then
          cVar1S10S8N043P003P040N021(0) <='1';
          else
          cVar1S10S8N043P003P040N021(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='1' AND B( 8)='0' )then
          cVar1S11S8N043P003P040N021(0) <='1';
          else
          cVar1S11S8N043P003P040N021(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='1' AND B( 8)='0' )then
          cVar1S12S8N043P003P040N021(0) <='1';
          else
          cVar1S12S8N043P003P040N021(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='1' )then
          cVar1S13S8N043P003N040P026(0) <='1';
          else
          cVar1S13S8N043P003N040P026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='1' )then
          cVar1S14S8N043P003N040P026(0) <='1';
          else
          cVar1S14S8N043P003N040P026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='1' )then
          cVar1S15S8N043P003N040P026(0) <='1';
          else
          cVar1S15S8N043P003N040P026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='0' )then
          cVar1S16S8N043P003N040N026(0) <='1';
          else
          cVar1S16S8N043P003N040N026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='0' )then
          cVar1S17S8N043P003N040N026(0) <='1';
          else
          cVar1S17S8N043P003N040N026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='0' AND E( 7)='0' AND B(14)='0' )then
          cVar1S18S8N043P003N040N026(0) <='1';
          else
          cVar1S18S8N043P003N040N026(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='1' AND B(17)='1' )then
          cVar1S19S8N043P003P039P020nsss(0) <='1';
          else
          cVar1S19S8N043P003P039P020nsss(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='1' AND B(17)='0' )then
          cVar1S20S8N043P003P039N020(0) <='1';
          else
          cVar1S20S8N043P003P039N020(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='1' AND B(17)='0' )then
          cVar1S21S8N043P003P039N020(0) <='1';
          else
          cVar1S21S8N043P003P039N020(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='0' AND B( 9)='1' )then
          cVar1S22S8N043P003N039P036(0) <='1';
          else
          cVar1S22S8N043P003N039P036(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='0' AND B( 9)='0' )then
          cVar1S23S8N043P003N039N036(0) <='1';
          else
          cVar1S23S8N043P003N039N036(0) <='0';
          end if;
        if(D(14)='0' AND A( 8)='1' AND D(15)='0' AND B( 9)='0' )then
          cVar1S24S8N043P003N039N036(0) <='1';
          else
          cVar1S24S8N043P003N039N036(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='1' )then
          cVar1S0S9P032P015P062P059(0) <='1';
          else
          cVar1S0S9P032P015P062P059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='1' )then
          cVar1S1S9P032P015P062P059(0) <='1';
          else
          cVar1S1S9P032P015P062P059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='1' )then
          cVar1S2S9P032P015P062P059(0) <='1';
          else
          cVar1S2S9P032P015P062P059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='1' )then
          cVar1S3S9P032P015P062P059(0) <='1';
          else
          cVar1S3S9P032P015P062P059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='0' )then
          cVar1S4S9P032P015P062N059(0) <='1';
          else
          cVar1S4S9P032P015P062N059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='0' )then
          cVar1S5S9P032P015P062N059(0) <='1';
          else
          cVar1S5S9P032P015P062N059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='0' )then
          cVar1S6S9P032P015P062N059(0) <='1';
          else
          cVar1S6S9P032P015P062N059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND D(10)='0' )then
          cVar1S7S9P032P015P062N059(0) <='1';
          else
          cVar1S7S9P032P015P062N059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='1' AND D(11)='0' )then
          cVar1S8S9P032P015P062P055(0) <='1';
          else
          cVar1S8S9P032P015P062P055(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='1' AND D(11)='0' )then
          cVar1S9S9P032P015P062P055(0) <='1';
          else
          cVar1S9S9P032P015P062P055(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='1' AND D(10)='1' )then
          cVar1S10S9P032P015P063P059nsss(0) <='1';
          else
          cVar1S10S9P032P015P063P059nsss(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='1' AND D(10)='0' )then
          cVar1S11S9P032P015P063N059(0) <='1';
          else
          cVar1S11S9P032P015P063N059(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='1' )then
          cVar1S12S9P032P015N063P068(0) <='1';
          else
          cVar1S12S9P032P015N063P068(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='1' )then
          cVar1S13S9P032P015N063P068(0) <='1';
          else
          cVar1S13S9P032P015N063P068(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='0' )then
          cVar1S14S9P032P015N063N068(0) <='1';
          else
          cVar1S14S9P032P015N063N068(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='0' )then
          cVar1S15S9P032P015N063N068(0) <='1';
          else
          cVar1S15S9P032P015N063N068(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='0' )then
          cVar1S16S9P032P015N063N068(0) <='1';
          else
          cVar1S16S9P032P015N063N068(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND E( 0)='0' )then
          cVar1S17S9P032P015N063N068(0) <='1';
          else
          cVar1S17S9P032P015N063N068(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='1' AND D( 1)='1' )then
          cVar1S18S9N032P043P045P062nsss(0) <='1';
          else
          cVar1S18S9N032P043P045P062nsss(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='1' AND D( 1)='0' )then
          cVar1S19S9N032P043P045N062(0) <='1';
          else
          cVar1S19S9N032P043P045N062(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='1' AND D( 1)='0' )then
          cVar1S20S9N032P043P045N062(0) <='1';
          else
          cVar1S20S9N032P043P045N062(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='0' AND A( 7)='1' )then
          cVar1S21S9N032P043N045P005nsss(0) <='1';
          else
          cVar1S21S9N032P043N045P005nsss(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='0' AND A( 7)='0' )then
          cVar1S22S9N032P043N045N005(0) <='1';
          else
          cVar1S22S9N032P043N045N005(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='0' AND A( 7)='0' )then
          cVar1S23S9N032P043N045N005(0) <='1';
          else
          cVar1S23S9N032P043N045N005(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='1' AND E(14)='0' AND A( 7)='0' )then
          cVar1S24S9N032P043N045N005(0) <='1';
          else
          cVar1S24S9N032P043N045N005(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='1' AND B( 7)='1' )then
          cVar1S25S9N032N043P044P023nsss(0) <='1';
          else
          cVar1S25S9N032N043P044P023nsss(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S26S9N032N043P044N023(0) <='1';
          else
          cVar1S26S9N032N043P044N023(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S27S9N032N043P044N023(0) <='1';
          else
          cVar1S27S9N032N043P044N023(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S28S9N032N043P044N023(0) <='1';
          else
          cVar1S28S9N032N043P044N023(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S29S9N032N043N044P040(0) <='1';
          else
          cVar1S29S9N032N043N044P040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S30S9N032N043N044P040(0) <='1';
          else
          cVar1S30S9N032N043N044P040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S31S9N032N043N044P040(0) <='1';
          else
          cVar1S31S9N032N043N044P040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S32S9N032N043N044N040(0) <='1';
          else
          cVar1S32S9N032N043N044N040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S33S9N032N043N044N040(0) <='1';
          else
          cVar1S33S9N032N043N044N040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S34S9N032N043N044N040(0) <='1';
          else
          cVar1S34S9N032N043N044N040(0) <='0';
          end if;
        if(B(11)='0' AND D(14)='0' AND E( 6)='0' AND E( 7)='0' )then
          cVar1S35S9N032N043N044N040(0) <='1';
          else
          cVar1S35S9N032N043N044N040(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='1' )then
          cVar1S0S10P032P015P062P061(0) <='1';
          else
          cVar1S0S10P032P015P062P061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='1' )then
          cVar1S1S10P032P015P062P061(0) <='1';
          else
          cVar1S1S10P032P015P062P061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='1' )then
          cVar1S2S10P032P015P062P061(0) <='1';
          else
          cVar1S2S10P032P015P062P061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='1' )then
          cVar1S3S10P032P015P062P061(0) <='1';
          else
          cVar1S3S10P032P015P062P061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='0' )then
          cVar1S4S10P032P015P062N061(0) <='1';
          else
          cVar1S4S10P032P015P062N061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='0' AND E(10)='0' )then
          cVar1S5S10P032P015P062N061(0) <='1';
          else
          cVar1S5S10P032P015P062N061(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='1' AND D(11)='0' )then
          cVar1S6S10P032P015P062P055(0) <='1';
          else
          cVar1S6S10P032P015P062P055(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='0' AND D( 1)='1' AND D(11)='0' )then
          cVar1S7S10P032P015P062P055(0) <='1';
          else
          cVar1S7S10P032P015P062P055(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='1' AND E(11)='0' )then
          cVar1S8S10P032P015P063P057(0) <='1';
          else
          cVar1S8S10P032P015P063P057(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='1' AND E(11)='0' )then
          cVar1S9S10P032P015P063P057(0) <='1';
          else
          cVar1S9S10P032P015P063P057(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='1' AND E(11)='0' )then
          cVar1S10S10P032P015P063P057(0) <='1';
          else
          cVar1S10S10P032P015P063P057(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND A(10)='1' )then
          cVar1S11S10P032P015N063P018(0) <='1';
          else
          cVar1S11S10P032P015N063P018(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND A(10)='1' )then
          cVar1S12S10P032P015N063P018(0) <='1';
          else
          cVar1S12S10P032P015N063P018(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND A(10)='0' )then
          cVar1S13S10P032P015N063N018(0) <='1';
          else
          cVar1S13S10P032P015N063N018(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND A(10)='0' )then
          cVar1S14S10P032P015N063N018(0) <='1';
          else
          cVar1S14S10P032P015N063N018(0) <='0';
          end if;
        if(B(11)='1' AND A( 2)='1' AND D( 9)='0' AND A(10)='0' )then
          cVar1S15S10P032P015N063N018(0) <='1';
          else
          cVar1S15S10P032P015N063N018(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='1' )then
          cVar1S16S10N032P040P021nsss(0) <='1';
          else
          cVar1S16S10N032P040P021nsss(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S17S10N032P040N021P010(0) <='1';
          else
          cVar1S17S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S18S10N032P040N021P010(0) <='1';
          else
          cVar1S18S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S19S10N032P040N021P010(0) <='1';
          else
          cVar1S19S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S20S10N032P040N021P010(0) <='1';
          else
          cVar1S20S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='1' )then
          cVar1S21S10N032P040N021P010(0) <='1';
          else
          cVar1S21S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='1' AND B( 8)='0' AND A(14)='1' )then
          cVar1S22S10N032P040N021P010(0) <='1';
          else
          cVar1S22S10N032P040N021P010(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='1' )then
          cVar1S23S10N032N040P043P062(0) <='1';
          else
          cVar1S23S10N032N040P043P062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='1' )then
          cVar1S24S10N032N040P043P062(0) <='1';
          else
          cVar1S24S10N032N040P043P062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='0' )then
          cVar1S25S10N032N040P043N062(0) <='1';
          else
          cVar1S25S10N032N040P043N062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='0' )then
          cVar1S26S10N032N040P043N062(0) <='1';
          else
          cVar1S26S10N032N040P043N062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='0' )then
          cVar1S27S10N032N040P043N062(0) <='1';
          else
          cVar1S27S10N032N040P043N062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='1' AND D( 1)='0' )then
          cVar1S28S10N032N040P043N062(0) <='1';
          else
          cVar1S28S10N032N040P043N062(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='1' )then
          cVar1S29S10N032N040N043P033(0) <='1';
          else
          cVar1S29S10N032N040N043P033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='1' )then
          cVar1S30S10N032N040N043P033(0) <='1';
          else
          cVar1S30S10N032N040N043P033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='1' )then
          cVar1S31S10N032N040N043P033(0) <='1';
          else
          cVar1S31S10N032N040N043P033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='0' )then
          cVar1S32S10N032N040N043N033(0) <='1';
          else
          cVar1S32S10N032N040N043N033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='0' )then
          cVar1S33S10N032N040N043N033(0) <='1';
          else
          cVar1S33S10N032N040N043N033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='0' )then
          cVar1S34S10N032N040N043N033(0) <='1';
          else
          cVar1S34S10N032N040N043N033(0) <='0';
          end if;
        if(B(11)='0' AND E( 7)='0' AND D(14)='0' AND B( 2)='0' )then
          cVar1S35S10N032N040N043N033(0) <='1';
          else
          cVar1S35S10N032N040N043N033(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='1' AND D( 5)='1' )then
          cVar1S0S11P027P008P046nsss(0) <='1';
          else
          cVar1S0S11P027P008P046nsss(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='1' AND D( 5)='0' AND D( 4)='1' )then
          cVar1S1S11P027P008N046P050nsss(0) <='1';
          else
          cVar1S1S11P027P008N046P050nsss(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='1' AND D( 5)='0' AND D( 4)='0' )then
          cVar1S2S11P027P008N046N050(0) <='1';
          else
          cVar1S2S11P027P008N046N050(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='1' AND E( 4)='0' )then
          cVar1S3S11P027N008P050P052(0) <='1';
          else
          cVar1S3S11P027N008P050P052(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='1' AND E( 4)='1' )then
          cVar1S4S11P027N008P050P052(0) <='1';
          else
          cVar1S4S11P027N008P050P052(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='1' AND E( 4)='1' )then
          cVar1S5S11P027N008P050P052(0) <='1';
          else
          cVar1S5S11P027N008P050P052(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='0' AND A(10)='1' )then
          cVar1S6S11P027N008N050P018(0) <='1';
          else
          cVar1S6S11P027N008N050P018(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='0' AND A(10)='1' )then
          cVar1S7S11P027N008N050P018(0) <='1';
          else
          cVar1S7S11P027N008N050P018(0) <='0';
          end if;
        if(B( 5)='1' AND A(15)='0' AND D( 4)='0' AND A(10)='0' )then
          cVar1S8S11P027N008N050N018(0) <='1';
          else
          cVar1S8S11P027N008N050N018(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='1' AND A( 7)='1' )then
          cVar1S9S11N027P039P020P005nsss(0) <='1';
          else
          cVar1S9S11N027P039P020P005nsss(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='1' AND A( 7)='0' )then
          cVar1S10S11N027P039P020N005(0) <='1';
          else
          cVar1S10S11N027P039P020N005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='0' AND A( 3)='0' )then
          cVar1S11S11N027P039N020P013(0) <='1';
          else
          cVar1S11S11N027P039N020P013(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='0' AND A( 3)='0' )then
          cVar1S12S11N027P039N020P013(0) <='1';
          else
          cVar1S12S11N027P039N020P013(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='0' AND A( 3)='0' )then
          cVar1S13S11N027P039N020P013(0) <='1';
          else
          cVar1S13S11N027P039N020P013(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(17)='0' AND A( 3)='1' )then
          cVar1S14S11N027P039N020P013(0) <='1';
          else
          cVar1S14S11N027P039N020P013(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='0' AND B(10)='1' )then
          cVar1S15S11N027N039P020P034(0) <='1';
          else
          cVar1S15S11N027N039P020P034(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='0' AND B(10)='1' )then
          cVar1S16S11N027N039P020P034(0) <='1';
          else
          cVar1S16S11N027N039P020P034(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='0' AND B(10)='0' )then
          cVar1S17S11N027N039P020N034(0) <='1';
          else
          cVar1S17S11N027N039P020N034(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='0' AND B(10)='0' )then
          cVar1S18S11N027N039P020N034(0) <='1';
          else
          cVar1S18S11N027N039P020N034(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='0' AND B(10)='0' )then
          cVar1S19S11N027N039P020N034(0) <='1';
          else
          cVar1S19S11N027N039P020N034(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='1' AND E( 7)='1' )then
          cVar1S20S11N027N039P020P040(0) <='1';
          else
          cVar1S20S11N027N039P020P040(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='1' AND E( 7)='1' )then
          cVar1S21S11N027N039P020P040(0) <='1';
          else
          cVar1S21S11N027N039P020P040(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='1' AND E( 7)='0' )then
          cVar1S22S11N027N039P020N040(0) <='1';
          else
          cVar1S22S11N027N039P020N040(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND B(17)='1' AND E( 7)='0' )then
          cVar1S23S11N027N039P020N040(0) <='1';
          else
          cVar1S23S11N027N039P020N040(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='0' )then
          cVar1S0S12P035P068P032P015(0) <='1';
          else
          cVar1S0S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='0' )then
          cVar1S1S12P035P068P032P015(0) <='1';
          else
          cVar1S1S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='0' )then
          cVar1S2S12P035P068P032P015(0) <='1';
          else
          cVar1S2S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='1' )then
          cVar1S3S12P035P068P032P015(0) <='1';
          else
          cVar1S3S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='1' )then
          cVar1S4S12P035P068P032P015(0) <='1';
          else
          cVar1S4S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='1' AND A( 2)='1' )then
          cVar1S5S12P035P068P032P015(0) <='1';
          else
          cVar1S5S12P035P068P032P015(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='1' )then
          cVar1S6S12P035P068N032P036(0) <='1';
          else
          cVar1S6S12P035P068N032P036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='1' )then
          cVar1S7S12P035P068N032P036(0) <='1';
          else
          cVar1S7S12P035P068N032P036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='1' )then
          cVar1S8S12P035P068N032P036(0) <='1';
          else
          cVar1S8S12P035P068N032P036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='1' )then
          cVar1S9S12P035P068N032P036(0) <='1';
          else
          cVar1S9S12P035P068N032P036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='0' )then
          cVar1S10S12P035P068N032N036(0) <='1';
          else
          cVar1S10S12P035P068N032N036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='0' )then
          cVar1S11S12P035P068N032N036(0) <='1';
          else
          cVar1S11S12P035P068N032N036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='0' )then
          cVar1S12S12P035P068N032N036(0) <='1';
          else
          cVar1S12S12P035P068N032N036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='0' AND B(11)='0' AND B( 9)='0' )then
          cVar1S13S12P035P068N032N036(0) <='1';
          else
          cVar1S13S12P035P068N032N036(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='0' )then
          cVar1S14S12P035P068P028P067(0) <='1';
          else
          cVar1S14S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='0' )then
          cVar1S15S12P035P068P028P067(0) <='1';
          else
          cVar1S15S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='0' )then
          cVar1S16S12P035P068P028P067(0) <='1';
          else
          cVar1S16S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='0' )then
          cVar1S17S12P035P068P028P067(0) <='1';
          else
          cVar1S17S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='1' )then
          cVar1S18S12P035P068P028P067(0) <='1';
          else
          cVar1S18S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='0' AND D( 8)='1' )then
          cVar1S19S12P035P068P028P067(0) <='1';
          else
          cVar1S19S12P035P068P028P067(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='1' AND A(10)='0' )then
          cVar1S20S12P035P068P028P018(0) <='1';
          else
          cVar1S20S12P035P068P028P018(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='1' AND A(10)='0' )then
          cVar1S21S12P035P068P028P018(0) <='1';
          else
          cVar1S21S12P035P068P028P018(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='1' AND A(10)='1' )then
          cVar1S22S12P035P068P028P018(0) <='1';
          else
          cVar1S22S12P035P068P028P018(0) <='0';
          end if;
        if(B( 1)='0' AND E( 0)='1' AND B(13)='1' AND A(10)='1' )then
          cVar1S23S12P035P068P028P018(0) <='1';
          else
          cVar1S23S12P035P068P028P018(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='0' )then
          cVar1S24S12P035P067P066P061(0) <='1';
          else
          cVar1S24S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='0' )then
          cVar1S25S12P035P067P066P061(0) <='1';
          else
          cVar1S25S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='0' )then
          cVar1S26S12P035P067P066P061(0) <='1';
          else
          cVar1S26S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='1' )then
          cVar1S27S12P035P067P066P061(0) <='1';
          else
          cVar1S27S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='1' )then
          cVar1S28S12P035P067P066P061(0) <='1';
          else
          cVar1S28S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='0' AND E(10)='1' )then
          cVar1S29S12P035P067P066P061(0) <='1';
          else
          cVar1S29S12P035P067P066P061(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='1' AND B( 0)='1' )then
          cVar1S30S12P035P067P066P037(0) <='1';
          else
          cVar1S30S12P035P067P066P037(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='1' AND B( 0)='1' )then
          cVar1S31S12P035P067P066P037(0) <='1';
          else
          cVar1S31S12P035P067P066P037(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='0' AND D( 0)='1' AND B( 0)='0' )then
          cVar1S32S12P035P067P066N037(0) <='1';
          else
          cVar1S32S12P035P067P066N037(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='1' AND A(12)='0' )then
          cVar1S33S12P035P067P068P014(0) <='1';
          else
          cVar1S33S12P035P067P068P014(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='1' AND A(12)='1' )then
          cVar1S34S12P035P067P068P014(0) <='1';
          else
          cVar1S34S12P035P067P068P014(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='1' AND A(12)='1' )then
          cVar1S35S12P035P067P068P014(0) <='1';
          else
          cVar1S35S12P035P067P068P014(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S36S12P035P067N068P018(0) <='1';
          else
          cVar1S36S12P035P067N068P018(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S37S12P035P067N068P018(0) <='1';
          else
          cVar1S37S12P035P067N068P018(0) <='0';
          end if;
        if(B( 1)='1' AND D( 8)='1' AND E( 0)='0' AND A(10)='1' )then
          cVar1S38S12P035P067N068P018(0) <='1';
          else
          cVar1S38S12P035P067N068P018(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='1' AND A(14)='1' )then
          cVar1S0S13P064P037P029P010(0) <='1';
          else
          cVar1S0S13P064P037P029P010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='1' AND A(14)='1' )then
          cVar1S1S13P064P037P029P010(0) <='1';
          else
          cVar1S1S13P064P037P029P010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='1' AND A(14)='0' )then
          cVar1S2S13P064P037P029N010(0) <='1';
          else
          cVar1S2S13P064P037P029N010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='1' AND A(14)='0' )then
          cVar1S3S13P064P037P029N010(0) <='1';
          else
          cVar1S3S13P064P037P029N010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='1' AND A(14)='0' )then
          cVar1S4S13P064P037P029N010(0) <='1';
          else
          cVar1S4S13P064P037P029N010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='1' )then
          cVar1S5S13P064P037N029P046(0) <='1';
          else
          cVar1S5S13P064P037N029P046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='1' )then
          cVar1S6S13P064P037N029P046(0) <='1';
          else
          cVar1S6S13P064P037N029P046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='1' )then
          cVar1S7S13P064P037N029P046(0) <='1';
          else
          cVar1S7S13P064P037N029P046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='0' )then
          cVar1S8S13P064P037N029N046(0) <='1';
          else
          cVar1S8S13P064P037N029N046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='0' )then
          cVar1S9S13P064P037N029N046(0) <='1';
          else
          cVar1S9S13P064P037N029N046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='0' AND B( 4)='0' AND D( 5)='0' )then
          cVar1S10S13P064P037N029N046(0) <='1';
          else
          cVar1S10S13P064P037N029N046(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='1' AND D( 0)='1' )then
          cVar1S11S13P064P037P067P066(0) <='1';
          else
          cVar1S11S13P064P037P067P066(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='1' AND D( 0)='1' )then
          cVar1S12S13P064P037P067P066(0) <='1';
          else
          cVar1S12S13P064P037P067P066(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S13S13P064P037P067N066(0) <='1';
          else
          cVar1S13S13P064P037P067N066(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S14S13P064P037P067N066(0) <='1';
          else
          cVar1S14S13P064P037P067N066(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S15S13P064P037P067N066(0) <='1';
          else
          cVar1S15S13P064P037P067N066(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='0' AND E( 2)='1' )then
          cVar1S16S13P064P037N067P060(0) <='1';
          else
          cVar1S16S13P064P037N067P060(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='0' AND E( 2)='1' )then
          cVar1S17S13P064P037N067P060(0) <='1';
          else
          cVar1S17S13P064P037N067P060(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='0' AND E( 2)='0' )then
          cVar1S18S13P064P037N067N060(0) <='1';
          else
          cVar1S18S13P064P037N067N060(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='0' AND E( 2)='0' )then
          cVar1S19S13P064P037N067N060(0) <='1';
          else
          cVar1S19S13P064P037N067N060(0) <='0';
          end if;
        if(E( 1)='0' AND B( 0)='1' AND D( 8)='0' AND E( 2)='0' )then
          cVar1S20S13P064P037N067N060(0) <='1';
          else
          cVar1S20S13P064P037N067N060(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='0' AND E(10)='0' )then
          cVar1S21S13P064P010P063P061(0) <='1';
          else
          cVar1S21S13P064P010P063P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='0' AND E(10)='0' )then
          cVar1S22S13P064P010P063P061(0) <='1';
          else
          cVar1S22S13P064P010P063P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='0' AND E(10)='0' )then
          cVar1S23S13P064P010P063P061(0) <='1';
          else
          cVar1S23S13P064P010P063P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='0' AND E(10)='1' )then
          cVar1S24S13P064P010P063P061(0) <='1';
          else
          cVar1S24S13P064P010P063P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='0' AND E(10)='1' )then
          cVar1S25S13P064P010P063P061(0) <='1';
          else
          cVar1S25S13P064P010P063P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='1' )then
          cVar1S26S13P064P010P063P018(0) <='1';
          else
          cVar1S26S13P064P010P063P018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='1' )then
          cVar1S27S13P064P010P063P018(0) <='1';
          else
          cVar1S27S13P064P010P063P018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='1' )then
          cVar1S28S13P064P010P063P018(0) <='1';
          else
          cVar1S28S13P064P010P063P018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='0' )then
          cVar1S29S13P064P010P063N018(0) <='1';
          else
          cVar1S29S13P064P010P063N018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='0' )then
          cVar1S30S13P064P010P063N018(0) <='1';
          else
          cVar1S30S13P064P010P063N018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='0' )then
          cVar1S31S13P064P010P063N018(0) <='1';
          else
          cVar1S31S13P064P010P063N018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='0' AND D( 9)='1' AND A(10)='0' )then
          cVar1S32S13P064P010P063N018(0) <='1';
          else
          cVar1S32S13P064P010P063N018(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='1' AND B(11)='1' AND E(10)='1' )then
          cVar1S33S13P064P010P032P061nsss(0) <='1';
          else
          cVar1S33S13P064P010P032P061nsss(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='1' AND B(11)='0' AND E(10)='0' )then
          cVar1S34S13P064P010N032P061(0) <='1';
          else
          cVar1S34S13P064P010N032P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='1' AND B(11)='0' AND E(10)='0' )then
          cVar1S35S13P064P010N032P061(0) <='1';
          else
          cVar1S35S13P064P010N032P061(0) <='0';
          end if;
        if(E( 1)='1' AND A(14)='1' AND B(11)='0' AND E(10)='0' )then
          cVar1S36S13P064P010N032P061(0) <='1';
          else
          cVar1S36S13P064P010N032P061(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='1' )then
          cVar1S0S14P030P057P063nsss(0) <='1';
          else
          cVar1S0S14P030P057P063nsss(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='0' )then
          cVar1S1S14P030P057N063P013(0) <='1';
          else
          cVar1S1S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='0' )then
          cVar1S2S14P030P057N063P013(0) <='1';
          else
          cVar1S2S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='0' )then
          cVar1S3S14P030P057N063P013(0) <='1';
          else
          cVar1S3S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='0' )then
          cVar1S4S14P030P057N063P013(0) <='1';
          else
          cVar1S4S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='1' )then
          cVar1S5S14P030P057N063P013(0) <='1';
          else
          cVar1S5S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='1' )then
          cVar1S6S14P030P057N063P013(0) <='1';
          else
          cVar1S6S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='1' AND D( 9)='0' AND A( 3)='1' )then
          cVar1S7S14P030P057N063P013(0) <='1';
          else
          cVar1S7S14P030P057N063P013(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='1' AND B( 0)='0' )then
          cVar1S8S14P030N057P056P037(0) <='1';
          else
          cVar1S8S14P030N057P056P037(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='1' AND B( 0)='0' )then
          cVar1S9S14P030N057P056P037(0) <='1';
          else
          cVar1S9S14P030N057P056P037(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='1' AND B( 0)='1' )then
          cVar1S10S14P030N057P056P037(0) <='1';
          else
          cVar1S10S14P030N057P056P037(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='0' AND E(10)='1' )then
          cVar1S11S14P030N057N056P061(0) <='1';
          else
          cVar1S11S14P030N057N056P061(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='0' AND E(10)='1' )then
          cVar1S12S14P030N057N056P061(0) <='1';
          else
          cVar1S12S14P030N057N056P061(0) <='0';
          end if;
        if(B(12)='1' AND E(11)='0' AND E( 3)='0' AND E(10)='0' )then
          cVar1S13S14P030N057N056N061(0) <='1';
          else
          cVar1S13S14P030N057N056N061(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='1' AND A(13)='0' )then
          cVar1S14S14N030P029P010P012(0) <='1';
          else
          cVar1S14S14N030P029P010P012(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='1' AND A(13)='0' )then
          cVar1S15S14N030P029P010P012(0) <='1';
          else
          cVar1S15S14N030P029P010P012(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='1' AND A(13)='1' )then
          cVar1S16S14N030P029P010P012(0) <='1';
          else
          cVar1S16S14N030P029P010P012(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='1' AND A(13)='1' )then
          cVar1S17S14N030P029P010P012(0) <='1';
          else
          cVar1S17S14N030P029P010P012(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='0' AND E(12)='1' )then
          cVar1S18S14N030P029N010P053(0) <='1';
          else
          cVar1S18S14N030P029N010P053(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='0' AND E(12)='1' )then
          cVar1S19S14N030P029N010P053(0) <='1';
          else
          cVar1S19S14N030P029N010P053(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='0' AND E(12)='1' )then
          cVar1S20S14N030P029N010P053(0) <='1';
          else
          cVar1S20S14N030P029N010P053(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='0' AND E(12)='0' )then
          cVar1S21S14N030P029N010N053(0) <='1';
          else
          cVar1S21S14N030P029N010N053(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='1' AND A(14)='0' AND E(12)='0' )then
          cVar1S22S14N030P029N010N053(0) <='1';
          else
          cVar1S22S14N030P029N010N053(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='1' AND E( 0)='0' )then
          cVar1S23S14N030N029P046P068(0) <='1';
          else
          cVar1S23S14N030N029P046P068(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='1' AND E( 0)='0' )then
          cVar1S24S14N030N029P046P068(0) <='1';
          else
          cVar1S24S14N030N029P046P068(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='1' AND E( 0)='1' )then
          cVar1S25S14N030N029P046P068(0) <='1';
          else
          cVar1S25S14N030N029P046P068(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='1' AND E( 0)='1' )then
          cVar1S26S14N030N029P046P068(0) <='1';
          else
          cVar1S26S14N030N029P046P068(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='1' AND E( 0)='1' )then
          cVar1S27S14N030N029P046P068(0) <='1';
          else
          cVar1S27S14N030N029P046P068(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='1' )then
          cVar1S28S14N030N029N046P037(0) <='1';
          else
          cVar1S28S14N030N029N046P037(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='1' )then
          cVar1S29S14N030N029N046P037(0) <='1';
          else
          cVar1S29S14N030N029N046P037(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='1' )then
          cVar1S30S14N030N029N046P037(0) <='1';
          else
          cVar1S30S14N030N029N046P037(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='0' )then
          cVar1S31S14N030N029N046N037(0) <='1';
          else
          cVar1S31S14N030N029N046N037(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='0' )then
          cVar1S32S14N030N029N046N037(0) <='1';
          else
          cVar1S32S14N030N029N046N037(0) <='0';
          end if;
        if(B(12)='0' AND B( 4)='0' AND D( 5)='0' AND B( 0)='0' )then
          cVar1S33S14N030N029N046N037(0) <='1';
          else
          cVar1S33S14N030N029N046N037(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='1' AND B(17)='1' )then
          cVar1S0S15P037P039P020nsss(0) <='1';
          else
          cVar1S0S15P037P039P020nsss(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S15P037P039N020P022nsss(0) <='1';
          else
          cVar1S1S15P037P039N020P022nsss(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S2S15P037P039N020N022(0) <='1';
          else
          cVar1S2S15P037P039N020N022(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S3S15P037P039N020N022(0) <='1';
          else
          cVar1S3S15P037P039N020N022(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S4S15P037P039N020N022(0) <='1';
          else
          cVar1S4S15P037P039N020N022(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='1' AND D( 4)='1' )then
          cVar1S5S15P037N039P027P050(0) <='1';
          else
          cVar1S5S15P037N039P027P050(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='1' AND D( 4)='1' )then
          cVar1S6S15P037N039P027P050(0) <='1';
          else
          cVar1S6S15P037N039P027P050(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='1' AND D( 4)='0' )then
          cVar1S7S15P037N039P027N050(0) <='1';
          else
          cVar1S7S15P037N039P027N050(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='1' AND D( 4)='0' )then
          cVar1S8S15P037N039P027N050(0) <='1';
          else
          cVar1S8S15P037N039P027N050(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='1' )then
          cVar1S9S15P037N039N027P026(0) <='1';
          else
          cVar1S9S15P037N039N027P026(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='1' )then
          cVar1S10S15P037N039N027P026(0) <='1';
          else
          cVar1S10S15P037N039N027P026(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='1' )then
          cVar1S11S15P037N039N027P026(0) <='1';
          else
          cVar1S11S15P037N039N027P026(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='0' )then
          cVar1S12S15P037N039N027N026(0) <='1';
          else
          cVar1S12S15P037N039N027N026(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='0' )then
          cVar1S13S15P037N039N027N026(0) <='1';
          else
          cVar1S13S15P037N039N027N026(0) <='0';
          end if;
        if(B( 0)='0' AND D(15)='0' AND B( 5)='0' AND B(14)='0' )then
          cVar1S14S15P037N039N027N026(0) <='1';
          else
          cVar1S14S15P037N039N027N026(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='1' AND A(11)='1' )then
          cVar1S15S15P037P030P057P016nsss(0) <='1';
          else
          cVar1S15S15P037P030P057P016nsss(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='1' AND A(11)='0' )then
          cVar1S16S15P037P030P057N016(0) <='1';
          else
          cVar1S16S15P037P030P057N016(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='1' AND A(11)='0' )then
          cVar1S17S15P037P030P057N016(0) <='1';
          else
          cVar1S17S15P037P030P057N016(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='1' AND A(11)='0' )then
          cVar1S18S15P037P030P057N016(0) <='1';
          else
          cVar1S18S15P037P030P057N016(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='0' AND E( 9)='1' )then
          cVar1S19S15P037P030N057P065(0) <='1';
          else
          cVar1S19S15P037P030N057P065(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='1' AND E(11)='0' AND E( 9)='1' )then
          cVar1S20S15P037P030N057P065(0) <='1';
          else
          cVar1S20S15P037P030N057P065(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='1' )then
          cVar1S21S15P037N030P055P009(0) <='1';
          else
          cVar1S21S15P037N030P055P009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='1' )then
          cVar1S22S15P037N030P055P009(0) <='1';
          else
          cVar1S22S15P037N030P055P009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='1' )then
          cVar1S23S15P037N030P055P009(0) <='1';
          else
          cVar1S23S15P037N030P055P009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='0' )then
          cVar1S24S15P037N030P055N009(0) <='1';
          else
          cVar1S24S15P037N030P055N009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='0' )then
          cVar1S25S15P037N030P055N009(0) <='1';
          else
          cVar1S25S15P037N030P055N009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='0' AND A( 5)='0' )then
          cVar1S26S15P037N030P055N009(0) <='1';
          else
          cVar1S26S15P037N030P055N009(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='1' AND B( 3)='1' )then
          cVar1S27S15P037N030P055P031(0) <='1';
          else
          cVar1S27S15P037N030P055P031(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='1' AND B( 3)='1' )then
          cVar1S28S15P037N030P055P031(0) <='1';
          else
          cVar1S28S15P037N030P055P031(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='1' AND B( 3)='0' )then
          cVar1S29S15P037N030P055N031(0) <='1';
          else
          cVar1S29S15P037N030P055N031(0) <='0';
          end if;
        if(B( 0)='1' AND B(12)='0' AND D(11)='1' AND B( 3)='0' )then
          cVar1S30S15P037N030P055N031(0) <='1';
          else
          cVar1S30S15P037N030P055N031(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' AND A( 6)='1' )then
          cVar1S0S16P043P022P007nsss(0) <='1';
          else
          cVar1S0S16P043P022P007nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' AND A( 6)='0' AND A( 0)='1' )then
          cVar1S1S16P043P022N007P019(0) <='1';
          else
          cVar1S1S16P043P022N007P019(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' AND A( 6)='0' AND A( 0)='1' )then
          cVar1S2S16P043P022N007P019(0) <='1';
          else
          cVar1S2S16P043P022N007P019(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' AND A( 6)='0' AND A( 0)='0' )then
          cVar1S3S16P043P022N007N019(0) <='1';
          else
          cVar1S3S16P043P022N007N019(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='1' AND A( 6)='0' AND A( 0)='0' )then
          cVar1S4S16P043P022N007N019(0) <='1';
          else
          cVar1S4S16P043P022N007N019(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND D( 1)='1' AND A(11)='1' )then
          cVar1S5S16P043N022P062P016nsss(0) <='1';
          else
          cVar1S5S16P043N022P062P016nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND D( 1)='1' AND A(11)='0' )then
          cVar1S6S16P043N022P062N016(0) <='1';
          else
          cVar1S6S16P043N022P062N016(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND D( 1)='0' AND A(16)='1' )then
          cVar1S7S16P043N022N062P006(0) <='1';
          else
          cVar1S7S16P043N022N062P006(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND D( 1)='0' AND A(16)='1' )then
          cVar1S8S16P043N022N062P006(0) <='1';
          else
          cVar1S8S16P043N022N062P006(0) <='0';
          end if;
        if(D(14)='1' AND B(16)='0' AND D( 1)='0' AND A(16)='0' )then
          cVar1S9S16P043N022N062N006(0) <='1';
          else
          cVar1S9S16P043N022N062N006(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='1' )then
          cVar1S10S16N043P030P057P063(0) <='1';
          else
          cVar1S10S16N043P030P057P063(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S11S16N043P030P057N063(0) <='1';
          else
          cVar1S11S16N043P030P057N063(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S12S16N043P030P057N063(0) <='1';
          else
          cVar1S12S16N043P030P057N063(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S13S16N043P030P057N063(0) <='1';
          else
          cVar1S13S16N043P030P057N063(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S14S16N043P030P057N063(0) <='1';
          else
          cVar1S14S16N043P030P057N063(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S15S16N043P030N057P029(0) <='1';
          else
          cVar1S15S16N043P030N057P029(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S16S16N043P030N057P029(0) <='1';
          else
          cVar1S16S16N043P030N057P029(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S17S16N043P030N057P029(0) <='1';
          else
          cVar1S17S16N043P030N057P029(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S18S16N043P030N057P029(0) <='1';
          else
          cVar1S18S16N043P030N057P029(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='1' )then
          cVar1S19S16N043P030N057P029(0) <='1';
          else
          cVar1S19S16N043P030N057P029(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='1' AND B(17)='1' )then
          cVar1S20S16N043N030P039P020(0) <='1';
          else
          cVar1S20S16N043N030P039P020(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='1' AND B(17)='1' )then
          cVar1S21S16N043N030P039P020(0) <='1';
          else
          cVar1S21S16N043N030P039P020(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='1' AND B(17)='0' )then
          cVar1S22S16N043N030P039N020(0) <='1';
          else
          cVar1S22S16N043N030P039N020(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='1' AND B(17)='0' )then
          cVar1S23S16N043N030P039N020(0) <='1';
          else
          cVar1S23S16N043N030P039N020(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='1' )then
          cVar1S24S16N043N030N039P034(0) <='1';
          else
          cVar1S24S16N043N030N039P034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='1' )then
          cVar1S25S16N043N030N039P034(0) <='1';
          else
          cVar1S25S16N043N030N039P034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='1' )then
          cVar1S26S16N043N030N039P034(0) <='1';
          else
          cVar1S26S16N043N030N039P034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='1' )then
          cVar1S27S16N043N030N039P034(0) <='1';
          else
          cVar1S27S16N043N030N039P034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='0' )then
          cVar1S28S16N043N030N039N034(0) <='1';
          else
          cVar1S28S16N043N030N039N034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='0' )then
          cVar1S29S16N043N030N039N034(0) <='1';
          else
          cVar1S29S16N043N030N039N034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='0' )then
          cVar1S30S16N043N030N039N034(0) <='1';
          else
          cVar1S30S16N043N030N039N034(0) <='0';
          end if;
        if(D(14)='0' AND B(12)='0' AND D(15)='0' AND B(10)='0' )then
          cVar1S31S16N043N030N039N034(0) <='1';
          else
          cVar1S31S16N043N030N039N034(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='0' AND B( 3)='0' )then
          cVar1S0S17P001P032P068P031(0) <='1';
          else
          cVar1S0S17P001P032P068P031(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='0' AND B( 3)='0' )then
          cVar1S1S17P001P032P068P031(0) <='1';
          else
          cVar1S1S17P001P032P068P031(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='0' AND B( 3)='0' )then
          cVar1S2S17P001P032P068P031(0) <='1';
          else
          cVar1S2S17P001P032P068P031(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='0' AND B( 3)='1' )then
          cVar1S3S17P001P032P068P031(0) <='1';
          else
          cVar1S3S17P001P032P068P031(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='0' AND B( 3)='1' )then
          cVar1S4S17P001P032P068P031(0) <='1';
          else
          cVar1S4S17P001P032P068P031(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='1' AND D( 0)='1' )then
          cVar1S5S17P001P032P068P066(0) <='1';
          else
          cVar1S5S17P001P032P068P066(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='1' AND D( 0)='1' )then
          cVar1S6S17P001P032P068P066(0) <='1';
          else
          cVar1S6S17P001P032P068P066(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='1' AND D( 0)='1' )then
          cVar1S7S17P001P032P068P066(0) <='1';
          else
          cVar1S7S17P001P032P068P066(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='1' AND E( 0)='1' AND D( 0)='0' )then
          cVar1S8S17P001P032P068N066(0) <='1';
          else
          cVar1S8S17P001P032P068N066(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='1' )then
          cVar1S9S17P001N032P000P019(0) <='1';
          else
          cVar1S9S17P001N032P000P019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='1' )then
          cVar1S10S17P001N032P000P019(0) <='1';
          else
          cVar1S10S17P001N032P000P019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='1' )then
          cVar1S11S17P001N032P000P019(0) <='1';
          else
          cVar1S11S17P001N032P000P019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='1' )then
          cVar1S12S17P001N032P000P019(0) <='1';
          else
          cVar1S12S17P001N032P000P019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='0' )then
          cVar1S13S17P001N032P000N019(0) <='1';
          else
          cVar1S13S17P001N032P000N019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='0' )then
          cVar1S14S17P001N032P000N019(0) <='1';
          else
          cVar1S14S17P001N032P000N019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='0' )then
          cVar1S15S17P001N032P000N019(0) <='1';
          else
          cVar1S15S17P001N032P000N019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='0' AND A( 0)='0' )then
          cVar1S16S17P001N032P000N019(0) <='1';
          else
          cVar1S16S17P001N032P000N019(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='1' )then
          cVar1S17S17P001N032P000P069(0) <='1';
          else
          cVar1S17S17P001N032P000P069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='1' )then
          cVar1S18S17P001N032P000P069(0) <='1';
          else
          cVar1S18S17P001N032P000P069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='1' )then
          cVar1S19S17P001N032P000P069(0) <='1';
          else
          cVar1S19S17P001N032P000P069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='0' )then
          cVar1S20S17P001N032P000N069(0) <='1';
          else
          cVar1S20S17P001N032P000N069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='0' )then
          cVar1S21S17P001N032P000N069(0) <='1';
          else
          cVar1S21S17P001N032P000N069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='0' )then
          cVar1S22S17P001N032P000N069(0) <='1';
          else
          cVar1S22S17P001N032P000N069(0) <='0';
          end if;
        if(A( 9)='0' AND B(11)='0' AND A(19)='1' AND E( 8)='0' )then
          cVar1S23S17P001N032P000N069(0) <='1';
          else
          cVar1S23S17P001N032P000N069(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='0' AND E(15)='1' )then
          cVar1S24S17P001P015P041nsss(0) <='1';
          else
          cVar1S24S17P001P015P041nsss(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='0' AND E(15)='0' AND D(10)='0' )then
          cVar1S25S17P001P015N041P059(0) <='1';
          else
          cVar1S25S17P001P015N041P059(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='0' AND E(15)='0' AND D(10)='0' )then
          cVar1S26S17P001P015N041P059(0) <='1';
          else
          cVar1S26S17P001P015N041P059(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='0' AND E(15)='0' AND D(10)='0' )then
          cVar1S27S17P001P015N041P059(0) <='1';
          else
          cVar1S27S17P001P015N041P059(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='0' AND E(15)='0' AND D(10)='0' )then
          cVar1S28S17P001P015N041P059(0) <='1';
          else
          cVar1S28S17P001P015N041P059(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='1' AND A(13)='1' AND D( 0)='0' )then
          cVar1S29S17P001P015P012P066(0) <='1';
          else
          cVar1S29S17P001P015P012P066(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='1' AND A(13)='1' AND D( 0)='0' )then
          cVar1S30S17P001P015P012P066(0) <='1';
          else
          cVar1S30S17P001P015P012P066(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='1' AND A(13)='1' AND D( 0)='1' )then
          cVar1S31S17P001P015P012P066(0) <='1';
          else
          cVar1S31S17P001P015P012P066(0) <='0';
          end if;
        if(A( 9)='1' AND A( 2)='1' AND A(13)='0' AND D( 9)='0' )then
          cVar1S32S17P001P015N012P063(0) <='1';
          else
          cVar1S32S17P001P015N012P063(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='1' )then
          cVar1S0S18P067P037P069P031(0) <='1';
          else
          cVar1S0S18P067P037P069P031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='1' )then
          cVar1S1S18P067P037P069P031(0) <='1';
          else
          cVar1S1S18P067P037P069P031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='1' )then
          cVar1S2S18P067P037P069P031(0) <='1';
          else
          cVar1S2S18P067P037P069P031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='1' )then
          cVar1S3S18P067P037P069P031(0) <='1';
          else
          cVar1S3S18P067P037P069P031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='0' )then
          cVar1S4S18P067P037P069N031(0) <='1';
          else
          cVar1S4S18P067P037P069N031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='0' )then
          cVar1S5S18P067P037P069N031(0) <='1';
          else
          cVar1S5S18P067P037P069N031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='0' )then
          cVar1S6S18P067P037P069N031(0) <='1';
          else
          cVar1S6S18P067P037P069N031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='0' AND B( 3)='0' )then
          cVar1S7S18P067P037P069N031(0) <='1';
          else
          cVar1S7S18P067P037P069N031(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='1' AND A( 1)='1' )then
          cVar1S8S18P067P037P069P017(0) <='1';
          else
          cVar1S8S18P067P037P069P017(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='1' AND A( 1)='1' )then
          cVar1S9S18P067P037P069P017(0) <='1';
          else
          cVar1S9S18P067P037P069P017(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='1' AND A( 1)='0' )then
          cVar1S10S18P067P037P069N017(0) <='1';
          else
          cVar1S10S18P067P037P069N017(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='0' AND E( 8)='1' AND A( 1)='0' )then
          cVar1S11S18P067P037P069N017(0) <='1';
          else
          cVar1S11S18P067P037P069N017(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='0' )then
          cVar1S12S18P067P037P016P018(0) <='1';
          else
          cVar1S12S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='0' )then
          cVar1S13S18P067P037P016P018(0) <='1';
          else
          cVar1S13S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='0' )then
          cVar1S14S18P067P037P016P018(0) <='1';
          else
          cVar1S14S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='0' )then
          cVar1S15S18P067P037P016P018(0) <='1';
          else
          cVar1S15S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='1' )then
          cVar1S16S18P067P037P016P018(0) <='1';
          else
          cVar1S16S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='1' AND A(10)='1' )then
          cVar1S17S18P067P037P016P018(0) <='1';
          else
          cVar1S17S18P067P037P016P018(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='0' AND A( 0)='1' )then
          cVar1S18S18P067P037N016P019(0) <='1';
          else
          cVar1S18S18P067P037N016P019(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='0' AND A( 0)='1' )then
          cVar1S19S18P067P037N016P019(0) <='1';
          else
          cVar1S19S18P067P037N016P019(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='0' AND A( 0)='0' )then
          cVar1S20S18P067P037N016N019(0) <='1';
          else
          cVar1S20S18P067P037N016N019(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='0' AND A( 0)='0' )then
          cVar1S21S18P067P037N016N019(0) <='1';
          else
          cVar1S21S18P067P037N016N019(0) <='0';
          end if;
        if(D( 8)='0' AND B( 0)='1' AND A(11)='0' AND A( 0)='0' )then
          cVar1S22S18P067P037N016N019(0) <='1';
          else
          cVar1S22S18P067P037N016N019(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='0' )then
          cVar1S23S18P067P007P069P036(0) <='1';
          else
          cVar1S23S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='0' )then
          cVar1S24S18P067P007P069P036(0) <='1';
          else
          cVar1S24S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='0' )then
          cVar1S25S18P067P007P069P036(0) <='1';
          else
          cVar1S25S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='1' )then
          cVar1S26S18P067P007P069P036(0) <='1';
          else
          cVar1S26S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='1' )then
          cVar1S27S18P067P007P069P036(0) <='1';
          else
          cVar1S27S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='1' AND B( 9)='1' )then
          cVar1S28S18P067P007P069P036(0) <='1';
          else
          cVar1S28S18P067P007P069P036(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='0' AND A(10)='1' )then
          cVar1S29S18P067P007N069P018(0) <='1';
          else
          cVar1S29S18P067P007N069P018(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='0' AND A(10)='1' )then
          cVar1S30S18P067P007N069P018(0) <='1';
          else
          cVar1S30S18P067P007N069P018(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='0' AND A(10)='0' )then
          cVar1S31S18P067P007N069N018(0) <='1';
          else
          cVar1S31S18P067P007N069N018(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='0' AND E( 8)='0' AND A(10)='0' )then
          cVar1S32S18P067P007N069N018(0) <='1';
          else
          cVar1S32S18P067P007N069N018(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='1' AND E(13)='1' )then
          cVar1S33S18P067P007P049nsss(0) <='1';
          else
          cVar1S33S18P067P007P049nsss(0) <='0';
          end if;
        if(D( 8)='1' AND A( 6)='1' AND E(13)='0' AND E( 6)='0' )then
          cVar1S34S18P067P007N049P044(0) <='1';
          else
          cVar1S34S18P067P007N049P044(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='0' AND E( 2)='1' )then
          cVar1S0S19P031P012P008P060(0) <='1';
          else
          cVar1S0S19P031P012P008P060(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='0' AND E( 2)='1' )then
          cVar1S1S19P031P012P008P060(0) <='1';
          else
          cVar1S1S19P031P012P008P060(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='0' AND E( 2)='0' )then
          cVar1S2S19P031P012P008N060(0) <='1';
          else
          cVar1S2S19P031P012P008N060(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='0' AND E( 2)='0' )then
          cVar1S3S19P031P012P008N060(0) <='1';
          else
          cVar1S3S19P031P012P008N060(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='0' AND E( 2)='0' )then
          cVar1S4S19P031P012P008N060(0) <='1';
          else
          cVar1S4S19P031P012P008N060(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='1' AND B( 2)='0' )then
          cVar1S5S19P031P012P008P033(0) <='1';
          else
          cVar1S5S19P031P012P008P033(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='1' AND A(15)='1' AND B( 2)='0' )then
          cVar1S6S19P031P012P008P033(0) <='1';
          else
          cVar1S6S19P031P012P008P033(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='1' AND D(10)='0' )then
          cVar1S7S19P031N012P013P059(0) <='1';
          else
          cVar1S7S19P031N012P013P059(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='1' AND D(10)='0' )then
          cVar1S8S19P031N012P013P059(0) <='1';
          else
          cVar1S8S19P031N012P013P059(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='1' AND D(10)='0' )then
          cVar1S9S19P031N012P013P059(0) <='1';
          else
          cVar1S9S19P031N012P013P059(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='1' AND D(10)='1' )then
          cVar1S10S19P031N012P013P059(0) <='1';
          else
          cVar1S10S19P031N012P013P059(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='1' AND D(10)='1' )then
          cVar1S11S19P031N012P013P059(0) <='1';
          else
          cVar1S11S19P031N012P013P059(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='0' AND D( 3)='1' )then
          cVar1S12S19P031N012N013P054(0) <='1';
          else
          cVar1S12S19P031N012N013P054(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='0' AND D( 3)='1' )then
          cVar1S13S19P031N012N013P054(0) <='1';
          else
          cVar1S13S19P031N012N013P054(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='0' AND D( 3)='0' )then
          cVar1S14S19P031N012N013N054(0) <='1';
          else
          cVar1S14S19P031N012N013N054(0) <='0';
          end if;
        if(B( 3)='1' AND A(13)='0' AND A( 3)='0' AND D( 3)='0' )then
          cVar1S15S19P031N012N013N054(0) <='1';
          else
          cVar1S15S19P031N012N013N054(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S16S19N031P036P007P037(0) <='1';
          else
          cVar1S16S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S17S19N031P036P007P037(0) <='1';
          else
          cVar1S17S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S18S19N031P036P007P037(0) <='1';
          else
          cVar1S18S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S19S19N031P036P007P037(0) <='1';
          else
          cVar1S19S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='1' )then
          cVar1S20S19N031P036P007P037(0) <='1';
          else
          cVar1S20S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='0' AND B( 0)='1' )then
          cVar1S21S19N031P036P007P037(0) <='1';
          else
          cVar1S21S19N031P036P007P037(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='1' AND A(15)='0' )then
          cVar1S22S19N031P036P007P008(0) <='1';
          else
          cVar1S22S19N031P036P007P008(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='1' AND A(15)='1' )then
          cVar1S23S19N031P036P007P008(0) <='1';
          else
          cVar1S23S19N031P036P007P008(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='1' AND A( 6)='1' AND A(15)='1' )then
          cVar1S24S19N031P036P007P008(0) <='1';
          else
          cVar1S24S19N031P036P007P008(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='1' )then
          cVar1S25S19N031N036P045P007(0) <='1';
          else
          cVar1S25S19N031N036P045P007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='1' )then
          cVar1S26S19N031N036P045P007(0) <='1';
          else
          cVar1S26S19N031N036P045P007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='1' )then
          cVar1S27S19N031N036P045P007(0) <='1';
          else
          cVar1S27S19N031N036P045P007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='0' )then
          cVar1S28S19N031N036P045N007(0) <='1';
          else
          cVar1S28S19N031N036P045N007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='0' )then
          cVar1S29S19N031N036P045N007(0) <='1';
          else
          cVar1S29S19N031N036P045N007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='1' AND A( 6)='0' )then
          cVar1S30S19N031N036P045N007(0) <='1';
          else
          cVar1S30S19N031N036P045N007(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='1' )then
          cVar1S31S19N031N036N045P053(0) <='1';
          else
          cVar1S31S19N031N036N045P053(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='1' )then
          cVar1S32S19N031N036N045P053(0) <='1';
          else
          cVar1S32S19N031N036N045P053(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='1' )then
          cVar1S33S19N031N036N045P053(0) <='1';
          else
          cVar1S33S19N031N036N045P053(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='0' )then
          cVar1S34S19N031N036N045N053(0) <='1';
          else
          cVar1S34S19N031N036N045N053(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='0' )then
          cVar1S35S19N031N036N045N053(0) <='1';
          else
          cVar1S35S19N031N036N045N053(0) <='0';
          end if;
        if(B( 3)='0' AND B( 9)='0' AND E(14)='0' AND E(12)='0' )then
          cVar1S36S19N031N036N045N053(0) <='1';
          else
          cVar1S36S19N031N036N045N053(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='1' AND A( 3)='0' )then
          cVar1S0S20P032P031P016P013(0) <='1';
          else
          cVar1S0S20P032P031P016P013(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='1' AND A( 3)='0' )then
          cVar1S1S20P032P031P016P013(0) <='1';
          else
          cVar1S1S20P032P031P016P013(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='1' AND A( 3)='0' )then
          cVar1S2S20P032P031P016P013(0) <='1';
          else
          cVar1S2S20P032P031P016P013(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='1' AND A( 3)='1' )then
          cVar1S3S20P032P031P016P013(0) <='1';
          else
          cVar1S3S20P032P031P016P013(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='1' AND A( 3)='1' )then
          cVar1S4S20P032P031P016P013(0) <='1';
          else
          cVar1S4S20P032P031P016P013(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S5S20P032P031N016P018(0) <='1';
          else
          cVar1S5S20P032P031N016P018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S6S20P032P031N016P018(0) <='1';
          else
          cVar1S6S20P032P031N016P018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S7S20P032P031N016P018(0) <='1';
          else
          cVar1S7S20P032P031N016P018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='0' )then
          cVar1S8S20P032P031N016N018(0) <='1';
          else
          cVar1S8S20P032P031N016N018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='0' )then
          cVar1S9S20P032P031N016N018(0) <='1';
          else
          cVar1S9S20P032P031N016N018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='0' AND A(11)='0' AND A(10)='0' )then
          cVar1S10S20P032P031N016N018(0) <='1';
          else
          cVar1S10S20P032P031N016N018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='1' AND A( 8)='0' AND A(10)='1' )then
          cVar1S11S20P032P031P003P018(0) <='1';
          else
          cVar1S11S20P032P031P003P018(0) <='0';
          end if;
        if(B(11)='1' AND B( 3)='1' AND A( 8)='0' AND A(10)='0' )then
          cVar1S12S20P032P031P003N018(0) <='1';
          else
          cVar1S12S20P032P031P003N018(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='1' )then
          cVar1S13S20N032P036P024P047(0) <='1';
          else
          cVar1S13S20N032P036P024P047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='1' )then
          cVar1S14S20N032P036P024P047(0) <='1';
          else
          cVar1S14S20N032P036P024P047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='1' )then
          cVar1S15S20N032P036P024P047(0) <='1';
          else
          cVar1S15S20N032P036P024P047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='0' )then
          cVar1S16S20N032P036P024N047(0) <='1';
          else
          cVar1S16S20N032P036P024N047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='0' )then
          cVar1S17S20N032P036P024N047(0) <='1';
          else
          cVar1S17S20N032P036P024N047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='1' AND D(13)='0' )then
          cVar1S18S20N032P036P024N047(0) <='1';
          else
          cVar1S18S20N032P036P024N047(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='1' )then
          cVar1S19S20N032P036N024P019(0) <='1';
          else
          cVar1S19S20N032P036N024P019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='1' )then
          cVar1S20S20N032P036N024P019(0) <='1';
          else
          cVar1S20S20N032P036N024P019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='1' )then
          cVar1S21S20N032P036N024P019(0) <='1';
          else
          cVar1S21S20N032P036N024P019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='1' )then
          cVar1S22S20N032P036N024P019(0) <='1';
          else
          cVar1S22S20N032P036N024P019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='0' )then
          cVar1S23S20N032P036N024N019(0) <='1';
          else
          cVar1S23S20N032P036N024N019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='0' )then
          cVar1S24S20N032P036N024N019(0) <='1';
          else
          cVar1S24S20N032P036N024N019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='0' )then
          cVar1S25S20N032P036N024N019(0) <='1';
          else
          cVar1S25S20N032P036N024N019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='0' AND B(15)='0' AND A( 0)='0' )then
          cVar1S26S20N032P036N024N019(0) <='1';
          else
          cVar1S26S20N032P036N024N019(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='0' AND B( 4)='0' )then
          cVar1S27S20N032P036P010P029(0) <='1';
          else
          cVar1S27S20N032P036P010P029(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='0' AND B( 4)='0' )then
          cVar1S28S20N032P036P010P029(0) <='1';
          else
          cVar1S28S20N032P036P010P029(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='0' AND B( 4)='0' )then
          cVar1S29S20N032P036P010P029(0) <='1';
          else
          cVar1S29S20N032P036P010P029(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='0' AND B( 4)='1' )then
          cVar1S30S20N032P036P010P029(0) <='1';
          else
          cVar1S30S20N032P036P010P029(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='0' AND B( 4)='1' )then
          cVar1S31S20N032P036P010P029(0) <='1';
          else
          cVar1S31S20N032P036P010P029(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='1' AND D(11)='1' )then
          cVar1S32S20N032P036P010P055(0) <='1';
          else
          cVar1S32S20N032P036P010P055(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='1' AND D(11)='1' )then
          cVar1S33S20N032P036P010P055(0) <='1';
          else
          cVar1S33S20N032P036P010P055(0) <='0';
          end if;
        if(B(11)='0' AND B( 9)='1' AND A(14)='1' AND D(11)='0' )then
          cVar1S34S20N032P036P010N055(0) <='1';
          else
          cVar1S34S20N032P036P010N055(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S0S21P024P047P066P063(0) <='1';
          else
          cVar1S0S21P024P047P066P063(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S1S21P024P047P066P063(0) <='1';
          else
          cVar1S1S21P024P047P066P063(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S2S21P024P047P066P063(0) <='1';
          else
          cVar1S2S21P024P047P066P063(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND A( 6)='1' )then
          cVar1S3S21P024P047P066P007nsss(0) <='1';
          else
          cVar1S3S21P024P047P066P007nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND A( 6)='0' )then
          cVar1S4S21P024P047P066N007(0) <='1';
          else
          cVar1S4S21P024P047P066N007(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND D(14)='1' )then
          cVar1S5S21P024N047P010P043(0) <='1';
          else
          cVar1S5S21P024N047P010P043(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND D(14)='1' )then
          cVar1S6S21P024N047P010P043(0) <='1';
          else
          cVar1S6S21P024N047P010P043(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND D(14)='0' )then
          cVar1S7S21P024N047P010N043(0) <='1';
          else
          cVar1S7S21P024N047P010N043(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND D(14)='0' )then
          cVar1S8S21P024N047P010N043(0) <='1';
          else
          cVar1S8S21P024N047P010N043(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND D(14)='0' )then
          cVar1S9S21P024N047P010N043(0) <='1';
          else
          cVar1S9S21P024N047P010N043(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B(11)='1' )then
          cVar1S10S21P024N047P010P032nsss(0) <='1';
          else
          cVar1S10S21P024N047P010P032nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B(11)='0' )then
          cVar1S11S21P024N047P010N032(0) <='1';
          else
          cVar1S11S21P024N047P010N032(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='1' )then
          cVar1S12S21N024P030P057P063(0) <='1';
          else
          cVar1S12S21N024P030P057P063(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S13S21N024P030P057N063(0) <='1';
          else
          cVar1S13S21N024P030P057N063(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S14S21N024P030P057N063(0) <='1';
          else
          cVar1S14S21N024P030P057N063(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S15S21N024P030P057N063(0) <='1';
          else
          cVar1S15S21N024P030P057N063(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='1' AND D( 9)='0' )then
          cVar1S16S21N024P030P057N063(0) <='1';
          else
          cVar1S16S21N024P030P057N063(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S17S21N024P030N057P029(0) <='1';
          else
          cVar1S17S21N024P030N057P029(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S18S21N024P030N057P029(0) <='1';
          else
          cVar1S18S21N024P030N057P029(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S19S21N024P030N057P029(0) <='1';
          else
          cVar1S19S21N024P030N057P029(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='1' AND E(11)='0' AND B( 4)='0' )then
          cVar1S20S21N024P030N057P029(0) <='1';
          else
          cVar1S20S21N024P030N057P029(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='0' )then
          cVar1S21S21N024N030P031P019(0) <='1';
          else
          cVar1S21S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='0' )then
          cVar1S22S21N024N030P031P019(0) <='1';
          else
          cVar1S22S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='0' )then
          cVar1S23S21N024N030P031P019(0) <='1';
          else
          cVar1S23S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='1' )then
          cVar1S24S21N024N030P031P019(0) <='1';
          else
          cVar1S24S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='1' )then
          cVar1S25S21N024N030P031P019(0) <='1';
          else
          cVar1S25S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='1' AND A( 0)='1' )then
          cVar1S26S21N024N030P031P019(0) <='1';
          else
          cVar1S26S21N024N030P031P019(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='0' )then
          cVar1S27S21N024N030N031P055(0) <='1';
          else
          cVar1S27S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='0' )then
          cVar1S28S21N024N030N031P055(0) <='1';
          else
          cVar1S28S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='0' )then
          cVar1S29S21N024N030N031P055(0) <='1';
          else
          cVar1S29S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='0' )then
          cVar1S30S21N024N030N031P055(0) <='1';
          else
          cVar1S30S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='1' )then
          cVar1S31S21N024N030N031P055(0) <='1';
          else
          cVar1S31S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='1' )then
          cVar1S32S21N024N030N031P055(0) <='1';
          else
          cVar1S32S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='0' AND B(12)='0' AND B( 3)='0' AND D(11)='1' )then
          cVar1S33S21N024N030N031P055(0) <='1';
          else
          cVar1S33S21N024N030N031P055(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' )then
          cVar1S0S22P024P047P066nsss(0) <='1';
          else
          cVar1S0S22P024P047P066nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND E( 0)='1' )then
          cVar1S1S22P024P047P066P068(0) <='1';
          else
          cVar1S1S22P024P047P066P068(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND E( 0)='1' )then
          cVar1S2S22P024P047P066P068(0) <='1';
          else
          cVar1S2S22P024P047P066P068(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND A( 9)='0' )then
          cVar1S3S22P024N047P010P001(0) <='1';
          else
          cVar1S3S22P024N047P010P001(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND A( 9)='0' )then
          cVar1S4S22P024N047P010P001(0) <='1';
          else
          cVar1S4S22P024N047P010P001(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND A( 9)='0' )then
          cVar1S5S22P024N047P010P001(0) <='1';
          else
          cVar1S5S22P024N047P010P001(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B(11)='1' )then
          cVar1S6S22P024N047P010P032nsss(0) <='1';
          else
          cVar1S6S22P024N047P010P032nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B(11)='0' )then
          cVar1S7S22P024N047P010N032(0) <='1';
          else
          cVar1S7S22P024N047P010N032(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='0' AND B(16)='1' )then
          cVar1S8S22N024P067P017P022(0) <='1';
          else
          cVar1S8S22N024P067P017P022(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='0' AND B(16)='1' )then
          cVar1S9S22N024P067P017P022(0) <='1';
          else
          cVar1S9S22N024P067P017P022(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='0' AND B(16)='1' )then
          cVar1S10S22N024P067P017P022(0) <='1';
          else
          cVar1S10S22N024P067P017P022(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='0' AND B(16)='0' )then
          cVar1S11S22N024P067P017N022(0) <='1';
          else
          cVar1S11S22N024P067P017N022(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='0' AND B(16)='0' )then
          cVar1S12S22N024P067P017N022(0) <='1';
          else
          cVar1S12S22N024P067P017N022(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='1' )then
          cVar1S13S22N024P067P017P014(0) <='1';
          else
          cVar1S13S22N024P067P017P014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='1' )then
          cVar1S14S22N024P067P017P014(0) <='1';
          else
          cVar1S14S22N024P067P017P014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='0' )then
          cVar1S15S22N024P067P017N014(0) <='1';
          else
          cVar1S15S22N024P067P017N014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='0' )then
          cVar1S16S22N024P067P017N014(0) <='1';
          else
          cVar1S16S22N024P067P017N014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='0' )then
          cVar1S17S22N024P067P017N014(0) <='1';
          else
          cVar1S17S22N024P067P017N014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='0' AND A( 1)='1' AND A(12)='0' )then
          cVar1S18S22N024P067P017N014(0) <='1';
          else
          cVar1S18S22N024P067P017N014(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='0' )then
          cVar1S19S22N024P067P060P064(0) <='1';
          else
          cVar1S19S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='0' )then
          cVar1S20S22N024P067P060P064(0) <='1';
          else
          cVar1S20S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='0' )then
          cVar1S21S22N024P067P060P064(0) <='1';
          else
          cVar1S21S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='0' )then
          cVar1S22S22N024P067P060P064(0) <='1';
          else
          cVar1S22S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='1' )then
          cVar1S23S22N024P067P060P064(0) <='1';
          else
          cVar1S23S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='1' AND E( 1)='1' )then
          cVar1S24S22N024P067P060P064(0) <='1';
          else
          cVar1S24S22N024P067P060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='1' )then
          cVar1S25S22N024P067N060P064(0) <='1';
          else
          cVar1S25S22N024P067N060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='1' )then
          cVar1S26S22N024P067N060P064(0) <='1';
          else
          cVar1S26S22N024P067N060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='1' )then
          cVar1S27S22N024P067N060P064(0) <='1';
          else
          cVar1S27S22N024P067N060P064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='0' )then
          cVar1S28S22N024P067N060N064(0) <='1';
          else
          cVar1S28S22N024P067N060N064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='0' )then
          cVar1S29S22N024P067N060N064(0) <='1';
          else
          cVar1S29S22N024P067N060N064(0) <='0';
          end if;
        if(B(15)='0' AND D( 8)='1' AND E( 2)='0' AND E( 1)='0' )then
          cVar1S30S22N024P067N060N064(0) <='1';
          else
          cVar1S30S22N024P067N060N064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND D( 9)='0' )then
          cVar1S0S23P024P047P066P063nsss(0) <='1';
          else
          cVar1S0S23P024P047P066P063nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND A( 6)='1' )then
          cVar1S1S23P024P047P066P007nsss(0) <='1';
          else
          cVar1S1S23P024P047P066P007nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND A( 6)='0' )then
          cVar1S2S23P024P047P066N007(0) <='1';
          else
          cVar1S2S23P024P047P066N007(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND A( 6)='0' )then
          cVar1S3S23P024P047P066N007(0) <='1';
          else
          cVar1S3S23P024P047P066N007(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E(13)='0' )then
          cVar1S4S23P024N047P010P049(0) <='1';
          else
          cVar1S4S23P024N047P010P049(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E(13)='0' )then
          cVar1S5S23P024N047P010P049(0) <='1';
          else
          cVar1S5S23P024N047P010P049(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E(13)='0' )then
          cVar1S6S23P024N047P010P049(0) <='1';
          else
          cVar1S6S23P024N047P010P049(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND A(10)='0' )then
          cVar1S7S23P024N047P010P018(0) <='1';
          else
          cVar1S7S23P024N047P010P018(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='0' AND A( 6)='0' )then
          cVar1S8S23N024P069P047P007(0) <='1';
          else
          cVar1S8S23N024P069P047P007(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='0' AND A( 6)='0' )then
          cVar1S9S23N024P069P047P007(0) <='1';
          else
          cVar1S9S23N024P069P047P007(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='0' AND A( 6)='0' )then
          cVar1S10S23N024P069P047P007(0) <='1';
          else
          cVar1S10S23N024P069P047P007(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='0' AND A( 6)='1' )then
          cVar1S11S23N024P069P047P007(0) <='1';
          else
          cVar1S11S23N024P069P047P007(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='1' AND D( 9)='0' )then
          cVar1S12S23N024P069P047P063(0) <='1';
          else
          cVar1S12S23N024P069P047P063(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='1' AND D( 9)='0' )then
          cVar1S13S23N024P069P047P063(0) <='1';
          else
          cVar1S13S23N024P069P047P063(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='1' AND D(13)='1' AND D( 9)='0' )then
          cVar1S14S23N024P069P047P063(0) <='1';
          else
          cVar1S14S23N024P069P047P063(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='1' AND D(14)='1' )then
          cVar1S15S23N024N069P022P043nsss(0) <='1';
          else
          cVar1S15S23N024N069P022P043nsss(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='1' AND D(14)='0' )then
          cVar1S16S23N024N069P022N043(0) <='1';
          else
          cVar1S16S23N024N069P022N043(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='1' AND D(14)='0' )then
          cVar1S17S23N024N069P022N043(0) <='1';
          else
          cVar1S17S23N024N069P022N043(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='0' AND B( 9)='1' )then
          cVar1S18S23N024N069N022P036(0) <='1';
          else
          cVar1S18S23N024N069N022P036(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='0' AND B( 9)='1' )then
          cVar1S19S23N024N069N022P036(0) <='1';
          else
          cVar1S19S23N024N069N022P036(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='0' AND B( 9)='0' )then
          cVar1S20S23N024N069N022N036(0) <='1';
          else
          cVar1S20S23N024N069N022N036(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='0' AND B( 9)='0' )then
          cVar1S21S23N024N069N022N036(0) <='1';
          else
          cVar1S21S23N024N069N022N036(0) <='0';
          end if;
        if(B(15)='0' AND E( 8)='0' AND B(16)='0' AND B( 9)='0' )then
          cVar1S22S23N024N069N022N036(0) <='1';
          else
          cVar1S22S23N024N069N022N036(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND E( 2)='0' )then
          cVar1S0S24P024P047P066P060(0) <='1';
          else
          cVar1S0S24P024P047P066P060(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND E( 2)='0' )then
          cVar1S1S24P024P047P066P060(0) <='1';
          else
          cVar1S1S24P024P047P066P060(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='0' AND E( 2)='1' )then
          cVar1S2S24P024P047P066P060psss(0) <='1';
          else
          cVar1S2S24P024P047P066P060psss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND E( 8)='1' )then
          cVar1S3S24P024P047P066P069nsss(0) <='1';
          else
          cVar1S3S24P024P047P066P069nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND E( 8)='0' )then
          cVar1S4S24P024P047P066N069(0) <='1';
          else
          cVar1S4S24P024P047P066N069(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='1' AND D( 0)='1' AND E( 8)='0' )then
          cVar1S5S24P024P047P066N069(0) <='1';
          else
          cVar1S5S24P024P047P066N069(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='1' )then
          cVar1S6S24P024N047P010P064(0) <='1';
          else
          cVar1S6S24P024N047P010P064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='1' )then
          cVar1S7S24P024N047P010P064(0) <='1';
          else
          cVar1S7S24P024N047P010P064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='1' )then
          cVar1S8S24P024N047P010P064(0) <='1';
          else
          cVar1S8S24P024N047P010P064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='0' )then
          cVar1S9S24P024N047P010N064(0) <='1';
          else
          cVar1S9S24P024N047P010N064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='0' )then
          cVar1S10S24P024N047P010N064(0) <='1';
          else
          cVar1S10S24P024N047P010N064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='0' AND E( 1)='0' )then
          cVar1S11S24P024N047P010N064(0) <='1';
          else
          cVar1S11S24P024N047P010N064(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B( 6)='1' )then
          cVar1S12S24P024N047P010P025nsss(0) <='1';
          else
          cVar1S12S24P024N047P010P025nsss(0) <='0';
          end if;
        if(B(15)='1' AND D(13)='0' AND A(14)='1' AND B( 6)='0' )then
          cVar1S13S24P024N047P010N025(0) <='1';
          else
          cVar1S13S24P024N047P010N025(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='1' AND B( 1)='0' )then
          cVar1S14S24N024P040P021P035nsss(0) <='1';
          else
          cVar1S14S24N024P040P021P035nsss(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='1' )then
          cVar1S15S24N024P040N021P037(0) <='1';
          else
          cVar1S15S24N024P040N021P037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='1' )then
          cVar1S16S24N024P040N021P037(0) <='1';
          else
          cVar1S16S24N024P040N021P037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='1' )then
          cVar1S17S24N024P040N021P037(0) <='1';
          else
          cVar1S17S24N024P040N021P037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='0' )then
          cVar1S18S24N024P040N021N037(0) <='1';
          else
          cVar1S18S24N024P040N021N037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='0' )then
          cVar1S19S24N024P040N021N037(0) <='1';
          else
          cVar1S19S24N024P040N021N037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='1' AND B( 8)='0' AND B( 0)='0' )then
          cVar1S20S24N024P040N021N037(0) <='1';
          else
          cVar1S20S24N024P040N021N037(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='0' AND D(15)='1' )then
          cVar1S21S24N024N040P002P039(0) <='1';
          else
          cVar1S21S24N024N040P002P039(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='0' AND D(15)='1' )then
          cVar1S22S24N024N040P002P039(0) <='1';
          else
          cVar1S22S24N024N040P002P039(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='0' AND D(15)='1' )then
          cVar1S23S24N024N040P002P039(0) <='1';
          else
          cVar1S23S24N024N040P002P039(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='0' AND D(15)='0' )then
          cVar1S24S24N024N040P002N039(0) <='1';
          else
          cVar1S24S24N024N040P002N039(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='0' AND D(15)='0' )then
          cVar1S25S24N024N040P002N039(0) <='1';
          else
          cVar1S25S24N024N040P002N039(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='1' AND E(12)='1' )then
          cVar1S26S24N024N040P002P053(0) <='1';
          else
          cVar1S26S24N024N040P002P053(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='1' AND E(12)='0' )then
          cVar1S27S24N024N040P002N053(0) <='1';
          else
          cVar1S27S24N024N040P002N053(0) <='0';
          end if;
        if(B(15)='0' AND E( 7)='0' AND A(18)='1' AND E(12)='0' )then
          cVar1S28S24N024N040P002N053(0) <='1';
          else
          cVar1S28S24N024N040P002N053(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='1' AND D( 1)='0' )then
          cVar1S0S25P001P031P012P062(0) <='1';
          else
          cVar1S0S25P001P031P012P062(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='1' AND D( 1)='0' )then
          cVar1S1S25P001P031P012P062(0) <='1';
          else
          cVar1S1S25P001P031P012P062(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='1' AND D( 1)='0' )then
          cVar1S2S25P001P031P012P062(0) <='1';
          else
          cVar1S2S25P001P031P012P062(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='1' AND D( 1)='0' )then
          cVar1S3S25P001P031P012P062(0) <='1';
          else
          cVar1S3S25P001P031P012P062(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='1' AND D( 1)='1' )then
          cVar1S4S25P001P031P012P062(0) <='1';
          else
          cVar1S4S25P001P031P012P062(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='0' AND A( 3)='1' )then
          cVar1S5S25P001P031N012P013(0) <='1';
          else
          cVar1S5S25P001P031N012P013(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='0' AND A( 3)='1' )then
          cVar1S6S25P001P031N012P013(0) <='1';
          else
          cVar1S6S25P001P031N012P013(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='0' AND A( 3)='0' )then
          cVar1S7S25P001P031N012N013(0) <='1';
          else
          cVar1S7S25P001P031N012N013(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='1' AND A(13)='0' AND A( 3)='0' )then
          cVar1S8S25P001P031N012N013(0) <='1';
          else
          cVar1S8S25P001P031N012N013(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='1' )then
          cVar1S9S25P001N031P030P063(0) <='1';
          else
          cVar1S9S25P001N031P030P063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='1' )then
          cVar1S10S25P001N031P030P063(0) <='1';
          else
          cVar1S10S25P001N031P030P063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='0' )then
          cVar1S11S25P001N031P030N063(0) <='1';
          else
          cVar1S11S25P001N031P030N063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='0' )then
          cVar1S12S25P001N031P030N063(0) <='1';
          else
          cVar1S12S25P001N031P030N063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='0' )then
          cVar1S13S25P001N031P030N063(0) <='1';
          else
          cVar1S13S25P001N031P030N063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='1' AND D( 9)='0' )then
          cVar1S14S25P001N031P030N063(0) <='1';
          else
          cVar1S14S25P001N031P030N063(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='0' )then
          cVar1S15S25P001N031N030P055(0) <='1';
          else
          cVar1S15S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='0' )then
          cVar1S16S25P001N031N030P055(0) <='1';
          else
          cVar1S16S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='0' )then
          cVar1S17S25P001N031N030P055(0) <='1';
          else
          cVar1S17S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='0' )then
          cVar1S18S25P001N031N030P055(0) <='1';
          else
          cVar1S18S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='1' )then
          cVar1S19S25P001N031N030P055(0) <='1';
          else
          cVar1S19S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='1' )then
          cVar1S20S25P001N031N030P055(0) <='1';
          else
          cVar1S20S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='1' )then
          cVar1S21S25P001N031N030P055(0) <='1';
          else
          cVar1S21S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='0' AND B( 3)='0' AND B(12)='0' AND D(11)='1' )then
          cVar1S22S25P001N031N030P055(0) <='1';
          else
          cVar1S22S25P001N031N030P055(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='1' AND A(13)='1' )then
          cVar1S23S25P001P023P067P012(0) <='1';
          else
          cVar1S23S25P001P023P067P012(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='1' AND A(13)='0' )then
          cVar1S24S25P001P023P067N012(0) <='1';
          else
          cVar1S24S25P001P023P067N012(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='1' AND A(13)='0' )then
          cVar1S25S25P001P023P067N012(0) <='1';
          else
          cVar1S25S25P001P023P067N012(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='0' AND E(15)='1' )then
          cVar1S26S25P001P023N067P041nsss(0) <='1';
          else
          cVar1S26S25P001P023N067P041nsss(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='0' AND E(15)='0' )then
          cVar1S27S25P001P023N067N041(0) <='1';
          else
          cVar1S27S25P001P023N067N041(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='0' AND E(15)='0' )then
          cVar1S28S25P001P023N067N041(0) <='1';
          else
          cVar1S28S25P001P023N067N041(0) <='0';
          end if;
        if(A( 9)='1' AND B( 7)='0' AND D( 8)='0' AND E(15)='0' )then
          cVar1S29S25P001P023N067N041(0) <='1';
          else
          cVar1S29S25P001P023N067N041(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='1' AND D( 2)='0' )then
          cVar1S0S26P015P017P034P058(0) <='1';
          else
          cVar1S0S26P015P017P034P058(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='1' AND D( 2)='1' )then
          cVar1S1S26P015P017P034P058(0) <='1';
          else
          cVar1S1S26P015P017P034P058(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='1' AND D( 2)='1' )then
          cVar1S2S26P015P017P034P058(0) <='1';
          else
          cVar1S2S26P015P017P034P058(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='0' AND B( 2)='1' )then
          cVar1S3S26P015P017N034P033(0) <='1';
          else
          cVar1S3S26P015P017N034P033(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='0' AND B( 2)='0' )then
          cVar1S4S26P015P017N034N033(0) <='1';
          else
          cVar1S4S26P015P017N034N033(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='0' AND B( 2)='0' )then
          cVar1S5S26P015P017N034N033(0) <='1';
          else
          cVar1S5S26P015P017N034N033(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='0' AND B( 2)='0' )then
          cVar1S6S26P015P017N034N033(0) <='1';
          else
          cVar1S6S26P015P017N034N033(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND B(10)='0' AND B( 2)='0' )then
          cVar1S7S26P015P017N034N033(0) <='1';
          else
          cVar1S7S26P015P017N034N033(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='0' AND A( 9)='0' )then
          cVar1S8S26P015P017P006P001(0) <='1';
          else
          cVar1S8S26P015P017P006P001(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='0' AND A( 9)='0' )then
          cVar1S9S26P015P017P006P001(0) <='1';
          else
          cVar1S9S26P015P017P006P001(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='0' AND A( 9)='0' )then
          cVar1S10S26P015P017P006P001(0) <='1';
          else
          cVar1S10S26P015P017P006P001(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='0' AND A( 9)='1' )then
          cVar1S11S26P015P017P006P001(0) <='1';
          else
          cVar1S11S26P015P017P006P001(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='1' AND D( 1)='1' )then
          cVar1S12S26P015P017P006P062(0) <='1';
          else
          cVar1S12S26P015P017P006P062(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='1' AND D( 1)='1' )then
          cVar1S13S26P015P017P006P062(0) <='1';
          else
          cVar1S13S26P015P017P006P062(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='1' AND D( 1)='0' )then
          cVar1S14S26P015P017P006N062(0) <='1';
          else
          cVar1S14S26P015P017P006N062(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='1' AND D( 1)='0' )then
          cVar1S15S26P015P017P006N062(0) <='1';
          else
          cVar1S15S26P015P017P006N062(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(16)='1' AND D( 1)='0' )then
          cVar1S16S26P015P017P006N062(0) <='1';
          else
          cVar1S16S26P015P017P006N062(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='1' AND A( 1)='1' )then
          cVar1S17S26N015P031P012P017(0) <='1';
          else
          cVar1S17S26N015P031P012P017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='1' AND A( 1)='1' )then
          cVar1S18S26N015P031P012P017(0) <='1';
          else
          cVar1S18S26N015P031P012P017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='1' AND A( 1)='0' )then
          cVar1S19S26N015P031P012N017(0) <='1';
          else
          cVar1S19S26N015P031P012N017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='1' AND A( 1)='0' )then
          cVar1S20S26N015P031P012N017(0) <='1';
          else
          cVar1S20S26N015P031P012N017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='1' AND A( 1)='0' )then
          cVar1S21S26N015P031P012N017(0) <='1';
          else
          cVar1S21S26N015P031P012N017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='1' )then
          cVar1S22S26N015P031N012P014(0) <='1';
          else
          cVar1S22S26N015P031N012P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='1' )then
          cVar1S23S26N015P031N012P014(0) <='1';
          else
          cVar1S23S26N015P031N012P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='1' )then
          cVar1S24S26N015P031N012P014(0) <='1';
          else
          cVar1S24S26N015P031N012P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='0' )then
          cVar1S25S26N015P031N012N014(0) <='1';
          else
          cVar1S25S26N015P031N012N014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='0' )then
          cVar1S26S26N015P031N012N014(0) <='1';
          else
          cVar1S26S26N015P031N012N014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='0' )then
          cVar1S27S26N015P031N012N014(0) <='1';
          else
          cVar1S27S26N015P031N012N014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='1' AND A(13)='0' AND A(12)='0' )then
          cVar1S28S26N015P031N012N014(0) <='1';
          else
          cVar1S28S26N015P031N012N014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='1' )then
          cVar1S29S26N015N031P030P059(0) <='1';
          else
          cVar1S29S26N015N031P030P059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='1' )then
          cVar1S30S26N015N031P030P059(0) <='1';
          else
          cVar1S30S26N015N031P030P059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='1' )then
          cVar1S31S26N015N031P030P059(0) <='1';
          else
          cVar1S31S26N015N031P030P059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='0' )then
          cVar1S32S26N015N031P030N059(0) <='1';
          else
          cVar1S32S26N015N031P030N059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='0' )then
          cVar1S33S26N015N031P030N059(0) <='1';
          else
          cVar1S33S26N015N031P030N059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='1' AND D(10)='0' )then
          cVar1S34S26N015N031P030N059(0) <='1';
          else
          cVar1S34S26N015N031P030N059(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S35S26N015N031N030P007(0) <='1';
          else
          cVar1S35S26N015N031N030P007(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S36S26N015N031N030P007(0) <='1';
          else
          cVar1S36S26N015N031N030P007(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S37S26N015N031N030P007(0) <='1';
          else
          cVar1S37S26N015N031N030P007(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S38S26N015N031N030N007(0) <='1';
          else
          cVar1S38S26N015N031N030N007(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S39S26N015N031N030N007(0) <='1';
          else
          cVar1S39S26N015N031N030N007(0) <='0';
          end if;
        if(A( 2)='0' AND B( 3)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S40S26N015N031N030N007(0) <='1';
          else
          cVar1S40S26N015N031N030N007(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='1' AND A( 6)='1' )then
          cVar1S0S27P002P022P043P007nsss(0) <='1';
          else
          cVar1S0S27P002P022P043P007nsss(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='1' AND A( 6)='0' )then
          cVar1S1S27P002P022P043N007(0) <='1';
          else
          cVar1S1S27P002P022P043N007(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='1' AND A( 6)='0' )then
          cVar1S2S27P002P022P043N007(0) <='1';
          else
          cVar1S2S27P002P022P043N007(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='1' AND A( 6)='0' )then
          cVar1S3S27P002P022P043N007(0) <='1';
          else
          cVar1S3S27P002P022P043N007(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='0' AND D( 6)='1' )then
          cVar1S4S27P002P022N043P042(0) <='1';
          else
          cVar1S4S27P002P022N043P042(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='0' AND D( 6)='1' )then
          cVar1S5S27P002P022N043P042(0) <='1';
          else
          cVar1S5S27P002P022N043P042(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='0' AND D( 6)='0' )then
          cVar1S6S27P002P022N043N042(0) <='1';
          else
          cVar1S6S27P002P022N043N042(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='1' AND D(14)='0' AND D( 6)='0' )then
          cVar1S7S27P002P022N043N042(0) <='1';
          else
          cVar1S7S27P002P022N043N042(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S8S27P002N022P027P026(0) <='1';
          else
          cVar1S8S27P002N022P027P026(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S9S27P002N022P027P026(0) <='1';
          else
          cVar1S9S27P002N022P027P026(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S10S27P002N022P027P026(0) <='1';
          else
          cVar1S10S27P002N022P027P026(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='1' AND B(14)='1' )then
          cVar1S11S27P002N022P027P026(0) <='1';
          else
          cVar1S11S27P002N022P027P026(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='1' )then
          cVar1S12S27P002N022N027P032(0) <='1';
          else
          cVar1S12S27P002N022N027P032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='1' )then
          cVar1S13S27P002N022N027P032(0) <='1';
          else
          cVar1S13S27P002N022N027P032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='1' )then
          cVar1S14S27P002N022N027P032(0) <='1';
          else
          cVar1S14S27P002N022N027P032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='0' )then
          cVar1S15S27P002N022N027N032(0) <='1';
          else
          cVar1S15S27P002N022N027N032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='0' )then
          cVar1S16S27P002N022N027N032(0) <='1';
          else
          cVar1S16S27P002N022N027N032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='0' )then
          cVar1S17S27P002N022N027N032(0) <='1';
          else
          cVar1S17S27P002N022N027N032(0) <='0';
          end if;
        if(A(18)='0' AND B(16)='0' AND B( 5)='0' AND B(11)='0' )then
          cVar1S18S27P002N022N027N032(0) <='1';
          else
          cVar1S18S27P002N022N027N032(0) <='0';
          end if;
        if(A(18)='1' AND E( 7)='1' AND B( 8)='1' )then
          cVar1S19S27P002P040P021nsss(0) <='1';
          else
          cVar1S19S27P002P040P021nsss(0) <='0';
          end if;
        if(A(18)='1' AND E( 7)='1' AND B( 8)='0' AND D( 7)='1' )then
          cVar1S20S27P002P040N021P038nsss(0) <='1';
          else
          cVar1S20S27P002P040N021P038nsss(0) <='0';
          end if;
        if(A(18)='1' AND E( 7)='0' AND D( 4)='0' AND E( 5)='1' )then
          cVar1S21S27P002N040P050P048(0) <='1';
          else
          cVar1S21S27P002N040P050P048(0) <='0';
          end if;
        if(A(18)='1' AND E( 7)='0' AND D( 4)='0' AND E( 5)='0' )then
          cVar1S22S27P002N040P050N048(0) <='1';
          else
          cVar1S22S27P002N040P050N048(0) <='0';
          end if;
        if(A(18)='1' AND E( 7)='0' AND D( 4)='0' AND E( 5)='0' )then
          cVar1S23S27P002N040P050N048(0) <='1';
          else
          cVar1S23S27P002N040P050N048(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='1' AND E(13)='0' )then
          cVar1S0S28P032P002P016P049(0) <='1';
          else
          cVar1S0S28P032P002P016P049(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='1' AND E(13)='0' )then
          cVar1S1S28P032P002P016P049(0) <='1';
          else
          cVar1S1S28P032P002P016P049(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='1' )then
          cVar1S2S28P032P002N016P063(0) <='1';
          else
          cVar1S2S28P032P002N016P063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='1' )then
          cVar1S3S28P032P002N016P063(0) <='1';
          else
          cVar1S3S28P032P002N016P063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='1' )then
          cVar1S4S28P032P002N016P063(0) <='1';
          else
          cVar1S4S28P032P002N016P063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='0' )then
          cVar1S5S28P032P002N016N063(0) <='1';
          else
          cVar1S5S28P032P002N016N063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='0' )then
          cVar1S6S28P032P002N016N063(0) <='1';
          else
          cVar1S6S28P032P002N016N063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='0' )then
          cVar1S7S28P032P002N016N063(0) <='1';
          else
          cVar1S7S28P032P002N016N063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='0' AND A(11)='0' AND D( 9)='0' )then
          cVar1S8S28P032P002N016N063(0) <='1';
          else
          cVar1S8S28P032P002N016N063(0) <='0';
          end if;
        if(B(11)='1' AND A(18)='1' AND A(10)='0' AND B( 1)='1' )then
          cVar1S9S28P032P002P018P035nsss(0) <='1';
          else
          cVar1S9S28P032P002P018P035nsss(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='1' AND B(14)='0' AND A(19)='0' )then
          cVar1S10S28N032P027P026P000(0) <='1';
          else
          cVar1S10S28N032P027P026P000(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='1' AND B(14)='0' AND A(19)='0' )then
          cVar1S11S28N032P027P026P000(0) <='1';
          else
          cVar1S11S28N032P027P026P000(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='1' AND B(14)='0' AND A(19)='1' )then
          cVar1S12S28N032P027P026P000(0) <='1';
          else
          cVar1S12S28N032P027P026P000(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='1' AND B(14)='1' AND B( 9)='0' )then
          cVar1S13S28N032P027P026P036(0) <='1';
          else
          cVar1S13S28N032P027P026P036(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='1' AND B(14)='1' AND B( 9)='0' )then
          cVar1S14S28N032P027P026P036(0) <='1';
          else
          cVar1S14S28N032P027P026P036(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='1' AND E( 8)='0' )then
          cVar1S15S28N032N027P022P069(0) <='1';
          else
          cVar1S15S28N032N027P022P069(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='1' AND E( 8)='0' )then
          cVar1S16S28N032N027P022P069(0) <='1';
          else
          cVar1S16S28N032N027P022P069(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='1' AND E( 8)='0' )then
          cVar1S17S28N032N027P022P069(0) <='1';
          else
          cVar1S17S28N032N027P022P069(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='1' AND E( 8)='1' )then
          cVar1S18S28N032N027P022P069(0) <='1';
          else
          cVar1S18S28N032N027P022P069(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='1' )then
          cVar1S19S28N032N027N022P030(0) <='1';
          else
          cVar1S19S28N032N027N022P030(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='1' )then
          cVar1S20S28N032N027N022P030(0) <='1';
          else
          cVar1S20S28N032N027N022P030(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='1' )then
          cVar1S21S28N032N027N022P030(0) <='1';
          else
          cVar1S21S28N032N027N022P030(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='0' )then
          cVar1S22S28N032N027N022N030(0) <='1';
          else
          cVar1S22S28N032N027N022N030(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='0' )then
          cVar1S23S28N032N027N022N030(0) <='1';
          else
          cVar1S23S28N032N027N022N030(0) <='0';
          end if;
        if(B(11)='0' AND B( 5)='0' AND B(16)='0' AND B(12)='0' )then
          cVar1S24S28N032N027N022N030(0) <='1';
          else
          cVar1S24S28N032N027N022N030(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='1' AND B( 1)='0' AND A(18)='1' )then
          cVar1S0S29P040P021P035P002nsss(0) <='1';
          else
          cVar1S0S29P040P021P035P002nsss(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='1' AND B( 1)='0' AND A(18)='0' )then
          cVar1S1S29P040P021P035N002(0) <='1';
          else
          cVar1S1S29P040P021P035N002(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='1' AND B( 1)='0' AND A(18)='0' )then
          cVar1S2S29P040P021P035N002(0) <='1';
          else
          cVar1S2S29P040P021P035N002(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='1' AND B( 1)='0' AND A(18)='0' )then
          cVar1S3S29P040P021P035N002(0) <='1';
          else
          cVar1S3S29P040P021P035N002(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='1' AND A( 7)='0' )then
          cVar1S4S29P040N021P037P005(0) <='1';
          else
          cVar1S4S29P040N021P037P005(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='1' AND A( 7)='0' )then
          cVar1S5S29P040N021P037P005(0) <='1';
          else
          cVar1S5S29P040N021P037P005(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='1' AND A( 7)='0' )then
          cVar1S6S29P040N021P037P005(0) <='1';
          else
          cVar1S6S29P040N021P037P005(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='0' AND A( 1)='1' )then
          cVar1S7S29P040N021N037P017(0) <='1';
          else
          cVar1S7S29P040N021N037P017(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='0' AND A( 1)='1' )then
          cVar1S8S29P040N021N037P017(0) <='1';
          else
          cVar1S8S29P040N021N037P017(0) <='0';
          end if;
        if(E( 7)='1' AND B( 8)='0' AND B( 0)='0' AND A( 1)='0' )then
          cVar1S9S29P040N021N037N017(0) <='1';
          else
          cVar1S9S29P040N021N037N017(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='0' )then
          cVar1S10S29N040P038P021P002(0) <='1';
          else
          cVar1S10S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='0' )then
          cVar1S11S29N040P038P021P002(0) <='1';
          else
          cVar1S11S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='0' )then
          cVar1S12S29N040P038P021P002(0) <='1';
          else
          cVar1S12S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='0' )then
          cVar1S13S29N040P038P021P002(0) <='1';
          else
          cVar1S13S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='1' )then
          cVar1S14S29N040P038P021P002(0) <='1';
          else
          cVar1S14S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='1' )then
          cVar1S15S29N040P038P021P002(0) <='1';
          else
          cVar1S15S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='0' AND A(18)='1' )then
          cVar1S16S29N040P038P021P002(0) <='1';
          else
          cVar1S16S29N040P038P021P002(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='1' AND A(14)='0' )then
          cVar1S17S29N040P038P021P010(0) <='1';
          else
          cVar1S17S29N040P038P021P010(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='0' AND B( 8)='1' AND A(14)='1' )then
          cVar1S18S29N040P038P021P010(0) <='1';
          else
          cVar1S18S29N040P038P021P010(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='1' AND B(14)='1' )then
          cVar1S19S29N040P038P026nsss(0) <='1';
          else
          cVar1S19S29N040P038P026nsss(0) <='0';
          end if;
        if(E( 7)='0' AND D( 7)='1' AND B(14)='0' AND D(10)='0' )then
          cVar1S20S29N040P038N026N059(0) <='1';
          else
          cVar1S20S29N040P038N026N059(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='1' AND E( 9)='0' )then
          cVar1S0S30P068P047P049P065(0) <='1';
          else
          cVar1S0S30P068P047P049P065(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='1' AND E( 9)='0' )then
          cVar1S1S30P068P047P049P065(0) <='1';
          else
          cVar1S1S30P068P047P049P065(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='1' AND E( 9)='0' )then
          cVar1S2S30P068P047P049P065(0) <='1';
          else
          cVar1S2S30P068P047P049P065(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='1' AND E( 9)='1' )then
          cVar1S3S30P068P047P049P065(0) <='1';
          else
          cVar1S3S30P068P047P049P065(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='1' AND E( 9)='1' )then
          cVar1S4S30P068P047P049P065(0) <='1';
          else
          cVar1S4S30P068P047P049P065(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='0' AND B(15)='1' )then
          cVar1S5S30P068P047N049P024(0) <='1';
          else
          cVar1S5S30P068P047N049P024(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='0' AND B(15)='0' )then
          cVar1S6S30P068P047N049N024(0) <='1';
          else
          cVar1S6S30P068P047N049N024(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='1' AND E(13)='0' AND B(15)='0' )then
          cVar1S7S30P068P047N049N024(0) <='1';
          else
          cVar1S7S30P068P047N049N024(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='1' AND D( 0)='0' )then
          cVar1S8S30P068N047P052P066(0) <='1';
          else
          cVar1S8S30P068N047P052P066(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='1' AND D( 0)='0' )then
          cVar1S9S30P068N047P052P066(0) <='1';
          else
          cVar1S9S30P068N047P052P066(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='1' AND D( 0)='0' )then
          cVar1S10S30P068N047P052P066(0) <='1';
          else
          cVar1S10S30P068N047P052P066(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='1' AND D( 0)='0' )then
          cVar1S11S30P068N047P052P066(0) <='1';
          else
          cVar1S11S30P068N047P052P066(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='1' AND D( 0)='1' )then
          cVar1S12S30P068N047P052P066(0) <='1';
          else
          cVar1S12S30P068N047P052P066(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='1' )then
          cVar1S13S30P068N047N052P036(0) <='1';
          else
          cVar1S13S30P068N047N052P036(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='1' )then
          cVar1S14S30P068N047N052P036(0) <='1';
          else
          cVar1S14S30P068N047N052P036(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='1' )then
          cVar1S15S30P068N047N052P036(0) <='1';
          else
          cVar1S15S30P068N047N052P036(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='0' )then
          cVar1S16S30P068N047N052N036(0) <='1';
          else
          cVar1S16S30P068N047N052N036(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='0' )then
          cVar1S17S30P068N047N052N036(0) <='1';
          else
          cVar1S17S30P068N047N052N036(0) <='0';
          end if;
        if(E( 0)='0' AND D(13)='0' AND E( 4)='0' AND B( 9)='0' )then
          cVar1S18S30P068N047N052N036(0) <='1';
          else
          cVar1S18S30P068N047N052N036(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S19S30P068P055P019P047(0) <='1';
          else
          cVar1S19S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S20S30P068P055P019P047(0) <='1';
          else
          cVar1S20S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S21S30P068P055P019P047(0) <='1';
          else
          cVar1S21S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S22S30P068P055P019P047(0) <='1';
          else
          cVar1S22S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='1' )then
          cVar1S23S30P068P055P019P047(0) <='1';
          else
          cVar1S23S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='1' )then
          cVar1S24S30P068P055P019P047(0) <='1';
          else
          cVar1S24S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='1' AND D(13)='1' )then
          cVar1S25S30P068P055P019P047(0) <='1';
          else
          cVar1S25S30P068P055P019P047(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='0' AND D(12)='1' )then
          cVar1S26S30P068P055N019P051(0) <='1';
          else
          cVar1S26S30P068P055N019P051(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='0' AND D(12)='1' )then
          cVar1S27S30P068P055N019P051(0) <='1';
          else
          cVar1S27S30P068P055N019P051(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='0' AND D(12)='0' )then
          cVar1S28S30P068P055N019N051(0) <='1';
          else
          cVar1S28S30P068P055N019N051(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='0' AND D(12)='0' )then
          cVar1S29S30P068P055N019N051(0) <='1';
          else
          cVar1S29S30P068P055N019N051(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='0' AND A( 0)='0' AND D(12)='0' )then
          cVar1S30S30P068P055N019N051(0) <='1';
          else
          cVar1S30S30P068P055N019N051(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='1' AND A(10)='0' )then
          cVar1S31S30P068P055P016P018(0) <='1';
          else
          cVar1S31S30P068P055P016P018(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='1' AND A(10)='1' )then
          cVar1S32S30P068P055P016P018(0) <='1';
          else
          cVar1S32S30P068P055P016P018(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='1' AND A(10)='1' )then
          cVar1S33S30P068P055P016P018(0) <='1';
          else
          cVar1S33S30P068P055P016P018(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='0' AND E(13)='0' )then
          cVar1S34S30P068P055N016P049(0) <='1';
          else
          cVar1S34S30P068P055N016P049(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='0' AND E(13)='0' )then
          cVar1S35S30P068P055N016P049(0) <='1';
          else
          cVar1S35S30P068P055N016P049(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='0' AND E(13)='0' )then
          cVar1S36S30P068P055N016P049(0) <='1';
          else
          cVar1S36S30P068P055N016P049(0) <='0';
          end if;
        if(E( 0)='1' AND D(11)='1' AND A(11)='0' AND E(13)='0' )then
          cVar1S37S30P068P055N016P049(0) <='1';
          else
          cVar1S37S30P068P055N016P049(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='0' )then
          cVar1S0S31P036P063P005P048(0) <='1';
          else
          cVar1S0S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='0' )then
          cVar1S1S31P036P063P005P048(0) <='1';
          else
          cVar1S1S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='0' )then
          cVar1S2S31P036P063P005P048(0) <='1';
          else
          cVar1S2S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='0' )then
          cVar1S3S31P036P063P005P048(0) <='1';
          else
          cVar1S3S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='1' )then
          cVar1S4S31P036P063P005P048(0) <='1';
          else
          cVar1S4S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='0' AND E( 5)='1' )then
          cVar1S5S31P036P063P005P048(0) <='1';
          else
          cVar1S5S31P036P063P005P048(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='1' AND B( 1)='1' )then
          cVar1S6S31P036P063P005P035nsss(0) <='1';
          else
          cVar1S6S31P036P063P005P035nsss(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='1' AND A( 7)='1' AND B( 1)='0' )then
          cVar1S7S31P036P063P005N035(0) <='1';
          else
          cVar1S7S31P036P063P005N035(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='1' )then
          cVar1S8S31P036N063P016P064(0) <='1';
          else
          cVar1S8S31P036N063P016P064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='1' )then
          cVar1S9S31P036N063P016P064(0) <='1';
          else
          cVar1S9S31P036N063P016P064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='1' )then
          cVar1S10S31P036N063P016P064(0) <='1';
          else
          cVar1S10S31P036N063P016P064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='1' )then
          cVar1S11S31P036N063P016P064(0) <='1';
          else
          cVar1S11S31P036N063P016P064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='0' )then
          cVar1S12S31P036N063P016N064(0) <='1';
          else
          cVar1S12S31P036N063P016N064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='0' )then
          cVar1S13S31P036N063P016N064(0) <='1';
          else
          cVar1S13S31P036N063P016N064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='0' )then
          cVar1S14S31P036N063P016N064(0) <='1';
          else
          cVar1S14S31P036N063P016N064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='1' AND E( 1)='0' )then
          cVar1S15S31P036N063P016N064(0) <='1';
          else
          cVar1S15S31P036N063P016N064(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S16S31P036N063N016P018(0) <='1';
          else
          cVar1S16S31P036N063N016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S17S31P036N063N016P018(0) <='1';
          else
          cVar1S17S31P036N063N016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S18S31P036N063N016P018(0) <='1';
          else
          cVar1S18S31P036N063N016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='1' )then
          cVar1S19S31P036N063N016P018(0) <='1';
          else
          cVar1S19S31P036N063N016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='0' )then
          cVar1S20S31P036N063N016N018(0) <='1';
          else
          cVar1S20S31P036N063N016N018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 9)='0' AND A(11)='0' AND A(10)='0' )then
          cVar1S21S31P036N063N016N018(0) <='1';
          else
          cVar1S21S31P036N063N016N018(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='0' AND E( 5)='0' )then
          cVar1S22S31N036P052P068P048(0) <='1';
          else
          cVar1S22S31N036P052P068P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='0' AND E( 5)='0' )then
          cVar1S23S31N036P052P068P048(0) <='1';
          else
          cVar1S23S31N036P052P068P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='0' AND E( 5)='0' )then
          cVar1S24S31N036P052P068P048(0) <='1';
          else
          cVar1S24S31N036P052P068P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='0' AND E( 5)='0' )then
          cVar1S25S31N036P052P068P048(0) <='1';
          else
          cVar1S25S31N036P052P068P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='0' AND E( 5)='1' )then
          cVar1S26S31N036P052P068P048(0) <='1';
          else
          cVar1S26S31N036P052P068P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='1' AND D(11)='0' )then
          cVar1S27S31N036P052P068P055(0) <='1';
          else
          cVar1S27S31N036P052P068P055(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='1' AND E( 0)='1' AND D(11)='0' )then
          cVar1S28S31N036P052P068P055(0) <='1';
          else
          cVar1S28S31N036P052P068P055(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S29S31N036N052P018P016(0) <='1';
          else
          cVar1S29S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S30S31N036N052P018P016(0) <='1';
          else
          cVar1S30S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S31S31N036N052P018P016(0) <='1';
          else
          cVar1S31S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S32S31N036N052P018P016(0) <='1';
          else
          cVar1S32S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='1' )then
          cVar1S33S31N036N052P018P016(0) <='1';
          else
          cVar1S33S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='1' )then
          cVar1S34S31N036N052P018P016(0) <='1';
          else
          cVar1S34S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='1' AND A(11)='1' )then
          cVar1S35S31N036N052P018P016(0) <='1';
          else
          cVar1S35S31N036N052P018P016(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='1' )then
          cVar1S36S31N036N052N018P014(0) <='1';
          else
          cVar1S36S31N036N052N018P014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='1' )then
          cVar1S37S31N036N052N018P014(0) <='1';
          else
          cVar1S37S31N036N052N018P014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='1' )then
          cVar1S38S31N036N052N018P014(0) <='1';
          else
          cVar1S38S31N036N052N018P014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='1' )then
          cVar1S39S31N036N052N018P014(0) <='1';
          else
          cVar1S39S31N036N052N018P014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='0' )then
          cVar1S40S31N036N052N018N014(0) <='1';
          else
          cVar1S40S31N036N052N018N014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='0' )then
          cVar1S41S31N036N052N018N014(0) <='1';
          else
          cVar1S41S31N036N052N018N014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='0' )then
          cVar1S42S31N036N052N018N014(0) <='1';
          else
          cVar1S42S31N036N052N018N014(0) <='0';
          end if;
        if(B( 9)='0' AND E( 4)='0' AND A(10)='0' AND A(12)='0' )then
          cVar1S43S31N036N052N018N014(0) <='1';
          else
          cVar1S43S31N036N052N018N014(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='1' AND A(16)='0' AND B( 5)='0' )then
          cVar1S0S32P036P066P006P027(0) <='1';
          else
          cVar1S0S32P036P066P006P027(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='1' AND A(16)='0' AND B( 5)='0' )then
          cVar1S1S32P036P066P006P027(0) <='1';
          else
          cVar1S1S32P036P066P006P027(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='1' AND A(16)='0' AND B( 5)='1' )then
          cVar1S2S32P036P066P006P027(0) <='1';
          else
          cVar1S2S32P036P066P006P027(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='1' AND A(16)='1' AND D(10)='0' )then
          cVar1S3S32P036P066P006P059(0) <='1';
          else
          cVar1S3S32P036P066P006P059(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='1' AND A(10)='0' )then
          cVar1S4S32P036N066P016P018(0) <='1';
          else
          cVar1S4S32P036N066P016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='1' AND A(10)='0' )then
          cVar1S5S32P036N066P016P018(0) <='1';
          else
          cVar1S5S32P036N066P016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='1' AND A(10)='0' )then
          cVar1S6S32P036N066P016P018(0) <='1';
          else
          cVar1S6S32P036N066P016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='1' AND A(10)='1' )then
          cVar1S7S32P036N066P016P018(0) <='1';
          else
          cVar1S7S32P036N066P016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='1' AND A(10)='1' )then
          cVar1S8S32P036N066P016P018(0) <='1';
          else
          cVar1S8S32P036N066P016P018(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='0' AND E( 0)='0' )then
          cVar1S9S32P036N066N016P068(0) <='1';
          else
          cVar1S9S32P036N066N016P068(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='0' AND E( 0)='0' )then
          cVar1S10S32P036N066N016P068(0) <='1';
          else
          cVar1S10S32P036N066N016P068(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='0' AND E( 0)='0' )then
          cVar1S11S32P036N066N016P068(0) <='1';
          else
          cVar1S11S32P036N066N016P068(0) <='0';
          end if;
        if(B( 9)='1' AND D( 0)='0' AND A(11)='0' AND E( 0)='1' )then
          cVar1S12S32P036N066N016P068(0) <='1';
          else
          cVar1S12S32P036N066N016P068(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='0' )then
          cVar1S13S32N036P060P048P063(0) <='1';
          else
          cVar1S13S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='0' )then
          cVar1S14S32N036P060P048P063(0) <='1';
          else
          cVar1S14S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='0' )then
          cVar1S15S32N036P060P048P063(0) <='1';
          else
          cVar1S15S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='1' )then
          cVar1S16S32N036P060P048P063(0) <='1';
          else
          cVar1S16S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='1' )then
          cVar1S17S32N036P060P048P063(0) <='1';
          else
          cVar1S17S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='1' )then
          cVar1S18S32N036P060P048P063(0) <='1';
          else
          cVar1S18S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='0' AND D( 9)='1' )then
          cVar1S19S32N036P060P048P063(0) <='1';
          else
          cVar1S19S32N036P060P048P063(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='1' AND A(16)='1' )then
          cVar1S20S32N036P060P048P006nsss(0) <='1';
          else
          cVar1S20S32N036P060P048P006nsss(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='1' AND E( 5)='1' AND A(16)='0' )then
          cVar1S21S32N036P060P048N006(0) <='1';
          else
          cVar1S21S32N036P060P048N006(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S22S32N036N060P058P054(0) <='1';
          else
          cVar1S22S32N036N060P058P054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S23S32N036N060P058P054(0) <='1';
          else
          cVar1S23S32N036N060P058P054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S24S32N036N060P058P054(0) <='1';
          else
          cVar1S24S32N036N060P058P054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S25S32N036N060P058P054(0) <='1';
          else
          cVar1S25S32N036N060P058P054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='0' )then
          cVar1S26S32N036N060P058N054(0) <='1';
          else
          cVar1S26S32N036N060P058N054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='0' )then
          cVar1S27S32N036N060P058N054(0) <='1';
          else
          cVar1S27S32N036N060P058N054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='0' AND D( 3)='0' )then
          cVar1S28S32N036N060P058N054(0) <='1';
          else
          cVar1S28S32N036N060P058N054(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='1' AND E( 3)='1' )then
          cVar1S29S32N036N060P058P056(0) <='1';
          else
          cVar1S29S32N036N060P058P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='1' AND E( 3)='1' )then
          cVar1S30S32N036N060P058P056(0) <='1';
          else
          cVar1S30S32N036N060P058P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='1' AND E( 3)='1' )then
          cVar1S31S32N036N060P058P056(0) <='1';
          else
          cVar1S31S32N036N060P058P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 2)='0' AND D( 2)='1' AND E( 3)='0' )then
          cVar1S32S32N036N060P058N056(0) <='1';
          else
          cVar1S32S32N036N060P058N056(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='1' AND A(10)='1' )then
          cVar1S0S33P034P049P026P018nsss(0) <='1';
          else
          cVar1S0S33P034P049P026P018nsss(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='1' AND A(10)='0' )then
          cVar1S1S33P034P049P026N018(0) <='1';
          else
          cVar1S1S33P034P049P026N018(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='1' AND A(10)='0' )then
          cVar1S2S33P034P049P026N018(0) <='1';
          else
          cVar1S2S33P034P049P026N018(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='0' AND B(15)='1' )then
          cVar1S3S33P034P049N026P024(0) <='1';
          else
          cVar1S3S33P034P049N026P024(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='0' AND B(15)='1' )then
          cVar1S4S33P034P049N026P024(0) <='1';
          else
          cVar1S4S33P034P049N026P024(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S5S33P034P049N026N024(0) <='1';
          else
          cVar1S5S33P034P049N026N024(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S6S33P034P049N026N024(0) <='1';
          else
          cVar1S6S33P034P049N026N024(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S7S33P034P049N026N024(0) <='1';
          else
          cVar1S7S33P034P049N026N024(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='1' )then
          cVar1S8S33P034N049P028P011(0) <='1';
          else
          cVar1S8S33P034N049P028P011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='1' )then
          cVar1S9S33P034N049P028P011(0) <='1';
          else
          cVar1S9S33P034N049P028P011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='0' )then
          cVar1S10S33P034N049P028N011(0) <='1';
          else
          cVar1S10S33P034N049P028N011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='0' )then
          cVar1S11S33P034N049P028N011(0) <='1';
          else
          cVar1S11S33P034N049P028N011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='0' )then
          cVar1S12S33P034N049P028N011(0) <='1';
          else
          cVar1S12S33P034N049P028N011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='1' AND A( 4)='0' )then
          cVar1S13S33P034N049P028N011(0) <='1';
          else
          cVar1S13S33P034N049P028N011(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='1' )then
          cVar1S14S33P034N049N028P066(0) <='1';
          else
          cVar1S14S33P034N049N028P066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='1' )then
          cVar1S15S33P034N049N028P066(0) <='1';
          else
          cVar1S15S33P034N049N028P066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='1' )then
          cVar1S16S33P034N049N028P066(0) <='1';
          else
          cVar1S16S33P034N049N028P066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='0' )then
          cVar1S17S33P034N049N028N066(0) <='1';
          else
          cVar1S17S33P034N049N028N066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='0' )then
          cVar1S18S33P034N049N028N066(0) <='1';
          else
          cVar1S18S33P034N049N028N066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='0' )then
          cVar1S19S33P034N049N028N066(0) <='1';
          else
          cVar1S19S33P034N049N028N066(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND B(13)='0' AND D( 0)='0' )then
          cVar1S20S33P034N049N028N066(0) <='1';
          else
          cVar1S20S33P034N049N028N066(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='1' )then
          cVar1S21S33P034P014P044P069(0) <='1';
          else
          cVar1S21S33P034P014P044P069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='1' )then
          cVar1S22S33P034P014P044P069(0) <='1';
          else
          cVar1S22S33P034P014P044P069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='1' )then
          cVar1S23S33P034P014P044P069(0) <='1';
          else
          cVar1S23S33P034P014P044P069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='0' )then
          cVar1S24S33P034P014P044N069(0) <='1';
          else
          cVar1S24S33P034P014P044N069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='0' )then
          cVar1S25S33P034P014P044N069(0) <='1';
          else
          cVar1S25S33P034P014P044N069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='1' AND E( 6)='0' AND E( 8)='0' )then
          cVar1S26S33P034P014P044N069(0) <='1';
          else
          cVar1S26S33P034P014P044N069(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='0' AND E(14)='1' AND D( 1)='1' )then
          cVar1S27S33P034N014P045P062nsss(0) <='1';
          else
          cVar1S27S33P034N014P045P062nsss(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='0' AND E(14)='1' AND D( 1)='0' )then
          cVar1S28S33P034N014P045N062(0) <='1';
          else
          cVar1S28S33P034N014P045N062(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='0' AND E(14)='0' AND D( 5)='0' )then
          cVar1S29S33P034N014N045P046(0) <='1';
          else
          cVar1S29S33P034N014N045P046(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='0' AND E(14)='0' AND D( 5)='0' )then
          cVar1S30S33P034N014N045P046(0) <='1';
          else
          cVar1S30S33P034N014N045P046(0) <='0';
          end if;
        if(B(10)='1' AND A(12)='0' AND E(14)='0' AND D( 5)='1' )then
          cVar1S31S33P034N014N045P046(0) <='1';
          else
          cVar1S31S33P034N014N045P046(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='1' AND D( 3)='0' )then
          cVar1S0S34P034P068P032P054(0) <='1';
          else
          cVar1S0S34P034P068P032P054(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='1' AND D( 3)='0' )then
          cVar1S1S34P034P068P032P054(0) <='1';
          else
          cVar1S1S34P034P068P032P054(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='1' AND D( 3)='0' )then
          cVar1S2S34P034P068P032P054(0) <='1';
          else
          cVar1S2S34P034P068P032P054(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='1' AND D( 3)='1' )then
          cVar1S3S34P034P068P032P054(0) <='1';
          else
          cVar1S3S34P034P068P032P054(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='1' AND D( 3)='1' )then
          cVar1S4S34P034P068P032P054(0) <='1';
          else
          cVar1S4S34P034P068P032P054(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='0' )then
          cVar1S5S34P034P068N032P059(0) <='1';
          else
          cVar1S5S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='0' )then
          cVar1S6S34P034P068N032P059(0) <='1';
          else
          cVar1S6S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='1' )then
          cVar1S7S34P034P068N032P059(0) <='1';
          else
          cVar1S7S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='1' )then
          cVar1S8S34P034P068N032P059(0) <='1';
          else
          cVar1S8S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='1' )then
          cVar1S9S34P034P068N032P059(0) <='1';
          else
          cVar1S9S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='0' AND B(11)='0' AND D(10)='1' )then
          cVar1S10S34P034P068N032P059(0) <='1';
          else
          cVar1S10S34P034P068N032P059(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar1S11S34P034P068P019P064(0) <='1';
          else
          cVar1S11S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar1S12S34P034P068P019P064(0) <='1';
          else
          cVar1S12S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar1S13S34P034P068P019P064(0) <='1';
          else
          cVar1S13S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='1' )then
          cVar1S14S34P034P068P019P064(0) <='1';
          else
          cVar1S14S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='1' )then
          cVar1S15S34P034P068P019P064(0) <='1';
          else
          cVar1S15S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='0' AND E( 1)='1' )then
          cVar1S16S34P034P068P019P064(0) <='1';
          else
          cVar1S16S34P034P068P019P064(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='0' )then
          cVar1S17S34P034P068P019P036(0) <='1';
          else
          cVar1S17S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='0' )then
          cVar1S18S34P034P068P019P036(0) <='1';
          else
          cVar1S18S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='0' )then
          cVar1S19S34P034P068P019P036(0) <='1';
          else
          cVar1S19S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='1' )then
          cVar1S20S34P034P068P019P036(0) <='1';
          else
          cVar1S20S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='1' )then
          cVar1S21S34P034P068P019P036(0) <='1';
          else
          cVar1S21S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='1' )then
          cVar1S22S34P034P068P019P036(0) <='1';
          else
          cVar1S22S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='0' AND E( 0)='1' AND A( 0)='1' AND B( 9)='1' )then
          cVar1S23S34P034P068P019P036(0) <='1';
          else
          cVar1S23S34P034P068P019P036(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S24S34P034P062P065P018(0) <='1';
          else
          cVar1S24S34P034P062P065P018(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S25S34P034P062P065P018(0) <='1';
          else
          cVar1S25S34P034P062P065P018(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S26S34P034P062P065P018(0) <='1';
          else
          cVar1S26S34P034P062P065P018(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='0' AND A(10)='1' )then
          cVar1S27S34P034P062P065P018(0) <='1';
          else
          cVar1S27S34P034P062P065P018(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='0' AND A(10)='1' )then
          cVar1S28S34P034P062P065P018(0) <='1';
          else
          cVar1S28S34P034P062P065P018(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S29S34P034P062P065P017(0) <='1';
          else
          cVar1S29S34P034P062P065P017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S30S34P034P062P065P017(0) <='1';
          else
          cVar1S30S34P034P062P065P017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='1' )then
          cVar1S31S34P034P062P065P017(0) <='1';
          else
          cVar1S31S34P034P062P065P017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S32S34P034P062P065N017(0) <='1';
          else
          cVar1S32S34P034P062P065N017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S33S34P034P062P065N017(0) <='1';
          else
          cVar1S33S34P034P062P065N017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S34S34P034P062P065N017(0) <='1';
          else
          cVar1S34S34P034P062P065N017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar1S35S34P034P062P065N017(0) <='1';
          else
          cVar1S35S34P034P062P065N017(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='1' )then
          cVar1S36S34P034N062P008P063(0) <='1';
          else
          cVar1S36S34P034N062P008P063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='1' )then
          cVar1S37S34P034N062P008P063(0) <='1';
          else
          cVar1S37S34P034N062P008P063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='1' )then
          cVar1S38S34P034N062P008P063(0) <='1';
          else
          cVar1S38S34P034N062P008P063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='0' )then
          cVar1S39S34P034N062P008N063(0) <='1';
          else
          cVar1S39S34P034N062P008N063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='0' )then
          cVar1S40S34P034N062P008N063(0) <='1';
          else
          cVar1S40S34P034N062P008N063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='0' AND D( 9)='0' )then
          cVar1S41S34P034N062P008N063(0) <='1';
          else
          cVar1S41S34P034N062P008N063(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='1' AND B(14)='1' )then
          cVar1S42S34P034N062P008P026(0) <='1';
          else
          cVar1S42S34P034N062P008P026(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='1' AND B(14)='0' )then
          cVar1S43S34P034N062P008N026(0) <='1';
          else
          cVar1S43S34P034N062P008N026(0) <='0';
          end if;
        if(B(10)='1' AND D( 1)='0' AND A(15)='1' AND B(14)='0' )then
          cVar1S44S34P034N062P008N026(0) <='1';
          else
          cVar1S44S34P034N062P008N026(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='1' AND A( 3)='1' )then
          cVar1S0S35P061P064P030P013nsss(0) <='1';
          else
          cVar1S0S35P061P064P030P013nsss(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='1' AND A( 3)='0' )then
          cVar1S1S35P061P064P030N013(0) <='1';
          else
          cVar1S1S35P061P064P030N013(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='1' AND A( 3)='0' )then
          cVar1S2S35P061P064P030N013(0) <='1';
          else
          cVar1S2S35P061P064P030N013(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S3S35P061P064N030P057(0) <='1';
          else
          cVar1S3S35P061P064N030P057(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S4S35P061P064N030P057(0) <='1';
          else
          cVar1S4S35P061P064N030P057(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S5S35P061P064N030P057(0) <='1';
          else
          cVar1S5S35P061P064N030P057(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S6S35P061P064N030P057(0) <='1';
          else
          cVar1S6S35P061P064N030P057(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='0' AND B(12)='0' AND E(11)='1' )then
          cVar1S7S35P061P064N030P057(0) <='1';
          else
          cVar1S7S35P061P064N030P057(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='1' AND D( 2)='0' AND A(15)='1' )then
          cVar1S8S35P061P064P058P008nsss(0) <='1';
          else
          cVar1S8S35P061P064P058P008nsss(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='1' AND D( 2)='0' AND A(15)='0' )then
          cVar1S9S35P061P064P058N008(0) <='1';
          else
          cVar1S9S35P061P064P058N008(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='1' AND D( 2)='0' AND A(15)='0' )then
          cVar1S10S35P061P064P058N008(0) <='1';
          else
          cVar1S10S35P061P064P058N008(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='1' AND D( 2)='0' AND A(15)='0' )then
          cVar1S11S35P061P064P058N008(0) <='1';
          else
          cVar1S11S35P061P064P058N008(0) <='0';
          end if;
        if(E(10)='1' AND E( 1)='1' AND D( 2)='1' AND D( 9)='1' )then
          cVar1S12S35P061P064P058P063(0) <='1';
          else
          cVar1S12S35P061P064P058P063(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='1' AND B(14)='0' AND A( 6)='0' )then
          cVar1S13S35N061P057P026P007(0) <='1';
          else
          cVar1S13S35N061P057P026P007(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='1' AND B(14)='0' AND A( 6)='0' )then
          cVar1S14S35N061P057P026P007(0) <='1';
          else
          cVar1S14S35N061P057P026P007(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='1' AND B(14)='0' AND A( 6)='0' )then
          cVar1S15S35N061P057P026P007(0) <='1';
          else
          cVar1S15S35N061P057P026P007(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='1' AND B(14)='0' AND A( 6)='1' )then
          cVar1S16S35N061P057P026P007(0) <='1';
          else
          cVar1S16S35N061P057P026P007(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='1' AND B(14)='1' AND B(12)='0' )then
          cVar1S17S35N061P057P026N030(0) <='1';
          else
          cVar1S17S35N061P057P026N030(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='0' )then
          cVar1S18S35N061N057P064P065(0) <='1';
          else
          cVar1S18S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='0' )then
          cVar1S19S35N061N057P064P065(0) <='1';
          else
          cVar1S19S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='0' )then
          cVar1S20S35N061N057P064P065(0) <='1';
          else
          cVar1S20S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='0' )then
          cVar1S21S35N061N057P064P065(0) <='1';
          else
          cVar1S21S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='1' )then
          cVar1S22S35N061N057P064P065(0) <='1';
          else
          cVar1S22S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='1' AND E( 9)='1' )then
          cVar1S23S35N061N057P064P065(0) <='1';
          else
          cVar1S23S35N061N057P064P065(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='0' AND D( 9)='1' )then
          cVar1S24S35N061N057N064P063(0) <='1';
          else
          cVar1S24S35N061N057N064P063(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='0' AND D( 9)='1' )then
          cVar1S25S35N061N057N064P063(0) <='1';
          else
          cVar1S25S35N061N057N064P063(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='0' AND D( 9)='0' )then
          cVar1S26S35N061N057N064N063(0) <='1';
          else
          cVar1S26S35N061N057N064N063(0) <='0';
          end if;
        if(E(10)='0' AND E(11)='0' AND E( 1)='0' AND D( 9)='0' )then
          cVar1S27S35N061N057N064N063(0) <='1';
          else
          cVar1S27S35N061N057N064N063(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='1' AND D( 0)='0' )then
          cVar1S0S36P063P062P065P066(0) <='1';
          else
          cVar1S0S36P063P062P065P066(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='1' AND D( 0)='0' )then
          cVar1S1S36P063P062P065P066(0) <='1';
          else
          cVar1S1S36P063P062P065P066(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='1' AND D( 0)='0' )then
          cVar1S2S36P063P062P065P066(0) <='1';
          else
          cVar1S2S36P063P062P065P066(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='1' AND D( 0)='0' )then
          cVar1S3S36P063P062P065P066(0) <='1';
          else
          cVar1S3S36P063P062P065P066(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='1' AND D( 0)='1' )then
          cVar1S4S36P063P062P065P066(0) <='1';
          else
          cVar1S4S36P063P062P065P066(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='0' AND A( 6)='0' )then
          cVar1S5S36P063P062N065P007(0) <='1';
          else
          cVar1S5S36P063P062N065P007(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='0' AND A( 6)='0' )then
          cVar1S6S36P063P062N065P007(0) <='1';
          else
          cVar1S6S36P063P062N065P007(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='0' AND A( 6)='0' )then
          cVar1S7S36P063P062N065P007(0) <='1';
          else
          cVar1S7S36P063P062N065P007(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND E( 9)='0' AND A( 6)='1' )then
          cVar1S8S36P063P062N065P007(0) <='1';
          else
          cVar1S8S36P063P062N065P007(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S9S36P063P062P048P054(0) <='1';
          else
          cVar1S9S36P063P062P048P054(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S10S36P063P062P048P054(0) <='1';
          else
          cVar1S10S36P063P062P048P054(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S11S36P063P062P048P054(0) <='1';
          else
          cVar1S11S36P063P062P048P054(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S12S36P063P062P048P054(0) <='1';
          else
          cVar1S12S36P063P062P048P054(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='0' AND D( 3)='1' )then
          cVar1S13S36P063P062P048P054(0) <='1';
          else
          cVar1S13S36P063P062P048P054(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 5)='1' AND D( 5)='1' )then
          cVar1S14S36P063P062P048P046(0) <='1';
          else
          cVar1S14S36P063P062P048P046(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='1' )then
          cVar1S15S36N063P067P064P019(0) <='1';
          else
          cVar1S15S36N063P067P064P019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='1' )then
          cVar1S16S36N063P067P064P019(0) <='1';
          else
          cVar1S16S36N063P067P064P019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='1' )then
          cVar1S17S36N063P067P064P019(0) <='1';
          else
          cVar1S17S36N063P067P064P019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='1' )then
          cVar1S18S36N063P067P064P019(0) <='1';
          else
          cVar1S18S36N063P067P064P019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='0' )then
          cVar1S19S36N063P067P064N019(0) <='1';
          else
          cVar1S19S36N063P067P064N019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='0' )then
          cVar1S20S36N063P067P064N019(0) <='1';
          else
          cVar1S20S36N063P067P064N019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='0' AND A( 0)='0' )then
          cVar1S21S36N063P067P064N019(0) <='1';
          else
          cVar1S21S36N063P067P064N019(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='1' AND B( 0)='1' )then
          cVar1S22S36N063P067P064P037(0) <='1';
          else
          cVar1S22S36N063P067P064P037(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='1' AND B( 0)='1' )then
          cVar1S23S36N063P067P064P037(0) <='1';
          else
          cVar1S23S36N063P067P064P037(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='1' AND B( 0)='0' )then
          cVar1S24S36N063P067P064N037(0) <='1';
          else
          cVar1S24S36N063P067P064N037(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='1' AND E( 1)='1' AND B( 0)='0' )then
          cVar1S25S36N063P067P064N037(0) <='1';
          else
          cVar1S25S36N063P067P064N037(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='1' AND D(12)='1' )then
          cVar1S26S36N063N067P053P051(0) <='1';
          else
          cVar1S26S36N063N067P053P051(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='1' AND D(12)='1' )then
          cVar1S27S36N063N067P053P051(0) <='1';
          else
          cVar1S27S36N063N067P053P051(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='1' AND D(12)='1' )then
          cVar1S28S36N063N067P053P051(0) <='1';
          else
          cVar1S28S36N063N067P053P051(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='1' AND D(12)='0' )then
          cVar1S29S36N063N067P053N051(0) <='1';
          else
          cVar1S29S36N063N067P053N051(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='0' AND B(16)='1' )then
          cVar1S30S36N063N067N053P022(0) <='1';
          else
          cVar1S30S36N063N067N053P022(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='0' AND B(16)='1' )then
          cVar1S31S36N063N067N053P022(0) <='1';
          else
          cVar1S31S36N063N067N053P022(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='0' AND B(16)='0' )then
          cVar1S32S36N063N067N053N022(0) <='1';
          else
          cVar1S32S36N063N067N053N022(0) <='0';
          end if;
        if(D( 9)='0' AND D( 8)='0' AND E(12)='0' AND B(16)='0' )then
          cVar1S33S36N063N067N053N022(0) <='1';
          else
          cVar1S33S36N063N067N053N022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='1' )then
          cVar1S0S37P065P067P000P068(0) <='1';
          else
          cVar1S0S37P065P067P000P068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='1' )then
          cVar1S1S37P065P067P000P068(0) <='1';
          else
          cVar1S1S37P065P067P000P068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='1' )then
          cVar1S2S37P065P067P000P068(0) <='1';
          else
          cVar1S2S37P065P067P000P068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='0' )then
          cVar1S3S37P065P067P000N068(0) <='1';
          else
          cVar1S3S37P065P067P000N068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='0' )then
          cVar1S4S37P065P067P000N068(0) <='1';
          else
          cVar1S4S37P065P067P000N068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='0' AND E( 0)='0' )then
          cVar1S5S37P065P067P000N068(0) <='1';
          else
          cVar1S5S37P065P067P000N068(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='0' AND A(19)='1' AND E(12)='0' )then
          cVar1S6S37P065P067P000P053(0) <='1';
          else
          cVar1S6S37P065P067P000P053(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='0' AND E( 3)='1' )then
          cVar1S7S37P065P067P062P056(0) <='1';
          else
          cVar1S7S37P065P067P062P056(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='0' AND E( 3)='0' )then
          cVar1S8S37P065P067P062N056(0) <='1';
          else
          cVar1S8S37P065P067P062N056(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='0' AND E( 3)='0' )then
          cVar1S9S37P065P067P062N056(0) <='1';
          else
          cVar1S9S37P065P067P062N056(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='0' AND E( 3)='0' )then
          cVar1S10S37P065P067P062N056(0) <='1';
          else
          cVar1S10S37P065P067P062N056(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='0' AND E( 3)='0' )then
          cVar1S11S37P065P067P062N056(0) <='1';
          else
          cVar1S11S37P065P067P062N056(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='1' AND A(10)='0' )then
          cVar1S12S37P065P067P062P018(0) <='1';
          else
          cVar1S12S37P065P067P062P018(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='1' AND A(10)='0' )then
          cVar1S13S37P065P067P062P018(0) <='1';
          else
          cVar1S13S37P065P067P062P018(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='1' AND A(10)='0' )then
          cVar1S14S37P065P067P062P018(0) <='1';
          else
          cVar1S14S37P065P067P062P018(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='1' AND A(10)='1' )then
          cVar1S15S37P065P067P062P018(0) <='1';
          else
          cVar1S15S37P065P067P062P018(0) <='0';
          end if;
        if(E( 9)='0' AND D( 8)='1' AND D( 1)='1' AND A(10)='1' )then
          cVar1S16S37P065P067P062P018(0) <='1';
          else
          cVar1S16S37P065P067P062P018(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='1' AND E( 8)='1' )then
          cVar1S17S37P065P060P058P069(0) <='1';
          else
          cVar1S17S37P065P060P058P069(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='1' AND E( 8)='0' )then
          cVar1S18S37P065P060P058N069(0) <='1';
          else
          cVar1S18S37P065P060P058N069(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='1' AND E( 8)='0' )then
          cVar1S19S37P065P060P058N069(0) <='1';
          else
          cVar1S19S37P065P060P058N069(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='1' AND E( 8)='0' )then
          cVar1S20S37P065P060P058N069(0) <='1';
          else
          cVar1S20S37P065P060P058N069(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='1' AND E( 8)='0' )then
          cVar1S21S37P065P060P058N069(0) <='1';
          else
          cVar1S21S37P065P060P058N069(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='1' AND D( 2)='0' AND A(10)='0' )then
          cVar1S22S37P065P060N058P018(0) <='1';
          else
          cVar1S22S37P065P060N058P018(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='1' )then
          cVar1S23S37P065N060P062P063(0) <='1';
          else
          cVar1S23S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='1' )then
          cVar1S24S37P065N060P062P063(0) <='1';
          else
          cVar1S24S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='1' )then
          cVar1S25S37P065N060P062P063(0) <='1';
          else
          cVar1S25S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='0' )then
          cVar1S26S37P065N060P062N063(0) <='1';
          else
          cVar1S26S37P065N060P062N063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='0' )then
          cVar1S27S37P065N060P062N063(0) <='1';
          else
          cVar1S27S37P065N060P062N063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='0' AND D( 9)='0' )then
          cVar1S28S37P065N060P062N063(0) <='1';
          else
          cVar1S28S37P065N060P062N063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='1' AND D( 9)='0' )then
          cVar1S29S37P065N060P062P063(0) <='1';
          else
          cVar1S29S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='1' AND D( 9)='0' )then
          cVar1S30S37P065N060P062P063(0) <='1';
          else
          cVar1S30S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='1' AND D( 9)='0' )then
          cVar1S31S37P065N060P062P063(0) <='1';
          else
          cVar1S31S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='1' AND D( 9)='0' )then
          cVar1S32S37P065N060P062P063(0) <='1';
          else
          cVar1S32S37P065N060P062P063(0) <='0';
          end if;
        if(E( 9)='1' AND E( 2)='0' AND D( 1)='1' AND D( 9)='1' )then
          cVar1S33S37P065N060P062P063(0) <='1';
          else
          cVar1S33S37P065N060P062P063(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='1' AND A(16)='0' )then
          cVar1S0S38P019P069P015P006(0) <='1';
          else
          cVar1S0S38P019P069P015P006(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='1' AND A(16)='0' )then
          cVar1S1S38P019P069P015P006(0) <='1';
          else
          cVar1S1S38P019P069P015P006(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='1' AND A(16)='1' )then
          cVar1S2S38P019P069P015P006(0) <='1';
          else
          cVar1S2S38P019P069P015P006(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='1' AND A(16)='1' )then
          cVar1S3S38P019P069P015P006(0) <='1';
          else
          cVar1S3S38P019P069P015P006(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='1' )then
          cVar1S4S38P019P069N015P009(0) <='1';
          else
          cVar1S4S38P019P069N015P009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='1' )then
          cVar1S5S38P019P069N015P009(0) <='1';
          else
          cVar1S5S38P019P069N015P009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='0' )then
          cVar1S6S38P019P069N015N009(0) <='1';
          else
          cVar1S6S38P019P069N015N009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='0' )then
          cVar1S7S38P019P069N015N009(0) <='1';
          else
          cVar1S7S38P019P069N015N009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='0' )then
          cVar1S8S38P019P069N015N009(0) <='1';
          else
          cVar1S8S38P019P069N015N009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 2)='0' AND A( 5)='0' )then
          cVar1S9S38P019P069N015N009(0) <='1';
          else
          cVar1S9S38P019P069N015N009(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='1' AND B(10)='0' )then
          cVar1S10S38P019N069P008P034(0) <='1';
          else
          cVar1S10S38P019N069P008P034(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='1' AND B(10)='0' )then
          cVar1S11S38P019N069P008P034(0) <='1';
          else
          cVar1S11S38P019N069P008P034(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='1' AND B(10)='0' )then
          cVar1S12S38P019N069P008P034(0) <='1';
          else
          cVar1S12S38P019N069P008P034(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='1' AND B(10)='0' )then
          cVar1S13S38P019N069P008P034(0) <='1';
          else
          cVar1S13S38P019N069P008P034(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='1' AND B(10)='1' )then
          cVar1S14S38P019N069P008P034(0) <='1';
          else
          cVar1S14S38P019N069P008P034(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='1' )then
          cVar1S15S38P019N069N008P016(0) <='1';
          else
          cVar1S15S38P019N069N008P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='1' )then
          cVar1S16S38P019N069N008P016(0) <='1';
          else
          cVar1S16S38P019N069N008P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='1' )then
          cVar1S17S38P019N069N008P016(0) <='1';
          else
          cVar1S17S38P019N069N008P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='0' )then
          cVar1S18S38P019N069N008N016(0) <='1';
          else
          cVar1S18S38P019N069N008N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='0' )then
          cVar1S19S38P019N069N008N016(0) <='1';
          else
          cVar1S19S38P019N069N008N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND A(15)='0' AND A(11)='0' )then
          cVar1S20S38P019N069N008N016(0) <='1';
          else
          cVar1S20S38P019N069N008N016(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S21S38N019P069P033P003(0) <='1';
          else
          cVar1S21S38N019P069P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S22S38N019P069P033P003(0) <='1';
          else
          cVar1S22S38N019P069P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S23S38N019P069P033P003(0) <='1';
          else
          cVar1S23S38N019P069P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S24S38N019P069P033P003(0) <='1';
          else
          cVar1S24S38N019P069P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='1' AND A( 8)='1' )then
          cVar1S25S38N019P069P033P003(0) <='1';
          else
          cVar1S25S38N019P069P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='1' )then
          cVar1S26S38N019P069N033P041(0) <='1';
          else
          cVar1S26S38N019P069N033P041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='1' )then
          cVar1S27S38N019P069N033P041(0) <='1';
          else
          cVar1S27S38N019P069N033P041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='1' )then
          cVar1S28S38N019P069N033P041(0) <='1';
          else
          cVar1S28S38N019P069N033P041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='0' )then
          cVar1S29S38N019P069N033N041(0) <='1';
          else
          cVar1S29S38N019P069N033N041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='0' )then
          cVar1S30S38N019P069N033N041(0) <='1';
          else
          cVar1S30S38N019P069N033N041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='0' AND B( 2)='0' AND E(15)='0' )then
          cVar1S31S38N019P069N033N041(0) <='1';
          else
          cVar1S31S38N019P069N033N041(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='1' AND D( 3)='0' )then
          cVar1S32S38N019P069P058P054(0) <='1';
          else
          cVar1S32S38N019P069P058P054(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='1' AND D( 3)='0' )then
          cVar1S33S38N019P069P058P054(0) <='1';
          else
          cVar1S33S38N019P069P058P054(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='1' AND D( 3)='0' )then
          cVar1S34S38N019P069P058P054(0) <='1';
          else
          cVar1S34S38N019P069P058P054(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S35S38N019P069N058P011(0) <='1';
          else
          cVar1S35S38N019P069N058P011(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S36S38N019P069N058P011(0) <='1';
          else
          cVar1S36S38N019P069N058P011(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S37S38N019P069N058P011(0) <='1';
          else
          cVar1S37S38N019P069N058P011(0) <='0';
          end if;
        if(A( 0)='0' AND E( 8)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S38S38N019P069N058P011(0) <='1';
          else
          cVar1S38S38N019P069N058P011(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='0' )then
          cVar1S0S39P011P069P058P067(0) <='1';
          else
          cVar1S0S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='0' )then
          cVar1S1S39P011P069P058P067(0) <='1';
          else
          cVar1S1S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='0' )then
          cVar1S2S39P011P069P058P067(0) <='1';
          else
          cVar1S2S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='0' )then
          cVar1S3S39P011P069P058P067(0) <='1';
          else
          cVar1S3S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='1' )then
          cVar1S4S39P011P069P058P067(0) <='1';
          else
          cVar1S4S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='1' )then
          cVar1S5S39P011P069P058P067(0) <='1';
          else
          cVar1S5S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='1' )then
          cVar1S6S39P011P069P058P067(0) <='1';
          else
          cVar1S6S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='0' AND D( 8)='1' )then
          cVar1S7S39P011P069P058P067(0) <='1';
          else
          cVar1S7S39P011P069P058P067(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='1' AND D( 1)='0' )then
          cVar1S8S39P011P069P058P062(0) <='1';
          else
          cVar1S8S39P011P069P058P062(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='1' AND D( 1)='0' )then
          cVar1S9S39P011P069P058P062(0) <='1';
          else
          cVar1S9S39P011P069P058P062(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='1' AND D( 1)='0' )then
          cVar1S10S39P011P069P058P062(0) <='1';
          else
          cVar1S10S39P011P069P058P062(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='1' AND D( 1)='1' )then
          cVar1S11S39P011P069P058P062(0) <='1';
          else
          cVar1S11S39P011P069P058P062(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='0' AND D( 2)='1' AND D( 1)='1' )then
          cVar1S12S39P011P069P058P062(0) <='1';
          else
          cVar1S12S39P011P069P058P062(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='1' )then
          cVar1S13S39P011P069P017P068(0) <='1';
          else
          cVar1S13S39P011P069P017P068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='1' )then
          cVar1S14S39P011P069P017P068(0) <='1';
          else
          cVar1S14S39P011P069P017P068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='1' )then
          cVar1S15S39P011P069P017P068(0) <='1';
          else
          cVar1S15S39P011P069P017P068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='1' )then
          cVar1S16S39P011P069P017P068(0) <='1';
          else
          cVar1S16S39P011P069P017P068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='0' )then
          cVar1S17S39P011P069P017N068(0) <='1';
          else
          cVar1S17S39P011P069P017N068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='1' AND E( 0)='0' )then
          cVar1S18S39P011P069P017N068(0) <='1';
          else
          cVar1S18S39P011P069P017N068(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='0' AND D(13)='1' )then
          cVar1S19S39P011P069N017P047(0) <='1';
          else
          cVar1S19S39P011P069N017P047(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='0' AND D(13)='0' )then
          cVar1S20S39P011P069N017N047(0) <='1';
          else
          cVar1S20S39P011P069N017N047(0) <='0';
          end if;
        if(A( 4)='0' AND E( 8)='1' AND A( 1)='0' AND D(13)='0' )then
          cVar1S21S39P011P069N017N047(0) <='1';
          else
          cVar1S21S39P011P069N017N047(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='0' )then
          cVar1S22S39P011P019P062P015(0) <='1';
          else
          cVar1S22S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='0' )then
          cVar1S23S39P011P019P062P015(0) <='1';
          else
          cVar1S23S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='0' )then
          cVar1S24S39P011P019P062P015(0) <='1';
          else
          cVar1S24S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='1' )then
          cVar1S25S39P011P019P062P015(0) <='1';
          else
          cVar1S25S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='1' )then
          cVar1S26S39P011P019P062P015(0) <='1';
          else
          cVar1S26S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='1' AND A( 2)='1' )then
          cVar1S27S39P011P019P062P015(0) <='1';
          else
          cVar1S27S39P011P019P062P015(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='0' AND E( 1)='0' )then
          cVar1S28S39P011P019N062P064(0) <='1';
          else
          cVar1S28S39P011P019N062P064(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='0' AND E( 1)='0' )then
          cVar1S29S39P011P019N062P064(0) <='1';
          else
          cVar1S29S39P011P019N062P064(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='0' AND E( 1)='0' )then
          cVar1S30S39P011P019N062P064(0) <='1';
          else
          cVar1S30S39P011P019N062P064(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='1' AND D( 1)='0' AND E( 1)='1' )then
          cVar1S31S39P011P019N062P064(0) <='1';
          else
          cVar1S31S39P011P019N062P064(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='1' AND E(10)='1' )then
          cVar1S32S39P011N019P060P061(0) <='1';
          else
          cVar1S32S39P011N019P060P061(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='1' AND E(10)='1' )then
          cVar1S33S39P011N019P060P061(0) <='1';
          else
          cVar1S33S39P011N019P060P061(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='1' AND E(10)='1' )then
          cVar1S34S39P011N019P060P061(0) <='1';
          else
          cVar1S34S39P011N019P060P061(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='1' AND E(10)='0' )then
          cVar1S35S39P011N019P060N061(0) <='1';
          else
          cVar1S35S39P011N019P060N061(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='1' AND E(10)='0' )then
          cVar1S36S39P011N019P060N061(0) <='1';
          else
          cVar1S36S39P011N019P060N061(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='0' AND E(13)='1' )then
          cVar1S37S39P011N019N060P049(0) <='1';
          else
          cVar1S37S39P011N019N060P049(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='0' AND E(13)='1' )then
          cVar1S38S39P011N019N060P049(0) <='1';
          else
          cVar1S38S39P011N019N060P049(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='0' AND E(13)='0' )then
          cVar1S39S39P011N019N060N049(0) <='1';
          else
          cVar1S39S39P011N019N060N049(0) <='0';
          end if;
        if(A( 4)='1' AND A( 0)='0' AND E( 2)='0' AND E(13)='0' )then
          cVar1S40S39P011N019N060N049(0) <='1';
          else
          cVar1S40S39P011N019N060N049(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='1' AND A( 4)='0' )then
          cVar1S0S40P069P053P067P011(0) <='1';
          else
          cVar1S0S40P069P053P067P011(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='1' AND A( 4)='0' )then
          cVar1S1S40P069P053P067P011(0) <='1';
          else
          cVar1S1S40P069P053P067P011(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='1' AND A( 4)='0' )then
          cVar1S2S40P069P053P067P011(0) <='1';
          else
          cVar1S2S40P069P053P067P011(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='1' AND A( 4)='1' )then
          cVar1S3S40P069P053P067P011(0) <='1';
          else
          cVar1S3S40P069P053P067P011(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='1' AND A( 4)='1' )then
          cVar1S4S40P069P053P067P011(0) <='1';
          else
          cVar1S4S40P069P053P067P011(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='1' )then
          cVar1S5S40P069P053N067P064(0) <='1';
          else
          cVar1S5S40P069P053N067P064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='1' )then
          cVar1S6S40P069P053N067P064(0) <='1';
          else
          cVar1S6S40P069P053N067P064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='1' )then
          cVar1S7S40P069P053N067P064(0) <='1';
          else
          cVar1S7S40P069P053N067P064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='0' )then
          cVar1S8S40P069P053N067N064(0) <='1';
          else
          cVar1S8S40P069P053N067N064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='0' )then
          cVar1S9S40P069P053N067N064(0) <='1';
          else
          cVar1S9S40P069P053N067N064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='0' )then
          cVar1S10S40P069P053N067N064(0) <='1';
          else
          cVar1S10S40P069P053N067N064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='0' AND D( 8)='0' AND E( 1)='0' )then
          cVar1S11S40P069P053N067N064(0) <='1';
          else
          cVar1S11S40P069P053N067N064(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='1' AND D(10)='0' AND E( 2)='1' )then
          cVar1S12S40P069P053P059P060nsss(0) <='1';
          else
          cVar1S12S40P069P053P059P060nsss(0) <='0';
          end if;
        if(E( 8)='1' AND E(12)='1' AND D(10)='0' AND E( 2)='0' )then
          cVar1S13S40P069P053P059N060(0) <='1';
          else
          cVar1S13S40P069P053P059N060(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='0' )then
          cVar1S14S40N069P031P013P065(0) <='1';
          else
          cVar1S14S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='0' )then
          cVar1S15S40N069P031P013P065(0) <='1';
          else
          cVar1S15S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='0' )then
          cVar1S16S40N069P031P013P065(0) <='1';
          else
          cVar1S16S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='1' )then
          cVar1S17S40N069P031P013P065(0) <='1';
          else
          cVar1S17S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='1' )then
          cVar1S18S40N069P031P013P065(0) <='1';
          else
          cVar1S18S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='1' AND E( 9)='1' )then
          cVar1S19S40N069P031P013P065(0) <='1';
          else
          cVar1S19S40N069P031P013P065(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='0' AND D( 2)='1' )then
          cVar1S20S40N069P031N013P058(0) <='1';
          else
          cVar1S20S40N069P031N013P058(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='0' AND D( 2)='1' )then
          cVar1S21S40N069P031N013P058(0) <='1';
          else
          cVar1S21S40N069P031N013P058(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='0' AND D( 2)='0' )then
          cVar1S22S40N069P031N013N058(0) <='1';
          else
          cVar1S22S40N069P031N013N058(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='0' AND D( 2)='0' )then
          cVar1S23S40N069P031N013N058(0) <='1';
          else
          cVar1S23S40N069P031N013N058(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='1' AND A( 3)='0' AND D( 2)='0' )then
          cVar1S24S40N069P031N013N058(0) <='1';
          else
          cVar1S24S40N069P031N013N058(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='1' AND E(10)='1' )then
          cVar1S25S40N069N031P030P061(0) <='1';
          else
          cVar1S25S40N069N031P030P061(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='1' AND E(10)='1' )then
          cVar1S26S40N069N031P030P061(0) <='1';
          else
          cVar1S26S40N069N031P030P061(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='1' AND E(10)='0' )then
          cVar1S27S40N069N031P030N061(0) <='1';
          else
          cVar1S27S40N069N031P030N061(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='1' AND E(10)='0' )then
          cVar1S28S40N069N031P030N061(0) <='1';
          else
          cVar1S28S40N069N031P030N061(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='1' AND E(10)='0' )then
          cVar1S29S40N069N031P030N061(0) <='1';
          else
          cVar1S29S40N069N031P030N061(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='0' )then
          cVar1S30S40N069N031N030P000(0) <='1';
          else
          cVar1S30S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='0' )then
          cVar1S31S40N069N031N030P000(0) <='1';
          else
          cVar1S31S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='0' )then
          cVar1S32S40N069N031N030P000(0) <='1';
          else
          cVar1S32S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='1' )then
          cVar1S33S40N069N031N030P000(0) <='1';
          else
          cVar1S33S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='1' )then
          cVar1S34S40N069N031N030P000(0) <='1';
          else
          cVar1S34S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='1' )then
          cVar1S35S40N069N031N030P000(0) <='1';
          else
          cVar1S35S40N069N031N030P000(0) <='0';
          end if;
        if(E( 8)='0' AND B( 3)='0' AND B(12)='0' AND A(19)='1' )then
          cVar1S36S40N069N031N030P000(0) <='1';
          else
          cVar1S36S40N069N031N030P000(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='1' AND E( 5)='1' )then
          cVar1S0S41P025P004P048nsss(0) <='1';
          else
          cVar1S0S41P025P004P048nsss(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='1' AND E( 5)='0' AND A(15)='0' )then
          cVar1S1S41P025P004N048P008nsss(0) <='1';
          else
          cVar1S1S41P025P004N048P008nsss(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='1' AND D( 8)='0' )then
          cVar1S2S41P025N004P007P067(0) <='1';
          else
          cVar1S2S41P025N004P007P067(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='1' AND D( 8)='0' )then
          cVar1S3S41P025N004P007P067(0) <='1';
          else
          cVar1S3S41P025N004P007P067(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='1' AND D( 8)='1' )then
          cVar1S4S41P025N004P007P067(0) <='1';
          else
          cVar1S4S41P025N004P007P067(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='0' AND B( 0)='1' )then
          cVar1S5S41P025N004N007P037(0) <='1';
          else
          cVar1S5S41P025N004N007P037(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='0' AND B( 0)='1' )then
          cVar1S6S41P025N004N007P037(0) <='1';
          else
          cVar1S6S41P025N004N007P037(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S7S41P025N004N007N037(0) <='1';
          else
          cVar1S7S41P025N004N007N037(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S8S41P025N004N007N037(0) <='1';
          else
          cVar1S8S41P025N004N007N037(0) <='0';
          end if;
        if(B( 6)='1' AND A(17)='0' AND A( 6)='0' AND B( 0)='0' )then
          cVar1S9S41P025N004N007N037(0) <='1';
          else
          cVar1S9S41P025N004N007N037(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='0' )then
          cVar1S10S41N025P062P058P055(0) <='1';
          else
          cVar1S10S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='0' )then
          cVar1S11S41N025P062P058P055(0) <='1';
          else
          cVar1S11S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='0' )then
          cVar1S12S41N025P062P058P055(0) <='1';
          else
          cVar1S12S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='1' )then
          cVar1S13S41N025P062P058P055(0) <='1';
          else
          cVar1S13S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='1' )then
          cVar1S14S41N025P062P058P055(0) <='1';
          else
          cVar1S14S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='1' )then
          cVar1S15S41N025P062P058P055(0) <='1';
          else
          cVar1S15S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='0' AND D(11)='1' )then
          cVar1S16S41N025P062P058P055(0) <='1';
          else
          cVar1S16S41N025P062P058P055(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='1' AND E(13)='0' )then
          cVar1S17S41N025P062P058P049(0) <='1';
          else
          cVar1S17S41N025P062P058P049(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='1' AND D( 2)='1' AND E(13)='0' )then
          cVar1S18S41N025P062P058P049(0) <='1';
          else
          cVar1S18S41N025P062P058P049(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S19S41N025N062P027P026(0) <='1';
          else
          cVar1S19S41N025N062P027P026(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S20S41N025N062P027P026(0) <='1';
          else
          cVar1S20S41N025N062P027P026(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S21S41N025N062P027P026(0) <='1';
          else
          cVar1S21S41N025N062P027P026(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='1' AND B(14)='0' )then
          cVar1S22S41N025N062P027P026(0) <='1';
          else
          cVar1S22S41N025N062P027P026(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='1' AND B(14)='1' )then
          cVar1S23S41N025N062P027P026(0) <='1';
          else
          cVar1S23S41N025N062P027P026(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S24S41N025N062N027P048(0) <='1';
          else
          cVar1S24S41N025N062N027P048(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S25S41N025N062N027P048(0) <='1';
          else
          cVar1S25S41N025N062N027P048(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S26S41N025N062N027P048(0) <='1';
          else
          cVar1S26S41N025N062N027P048(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S27S41N025N062N027P048(0) <='1';
          else
          cVar1S27S41N025N062N027P048(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='1' )then
          cVar1S28S41N025N062N027P048(0) <='1';
          else
          cVar1S28S41N025N062N027P048(0) <='0';
          end if;
        if(B( 6)='0' AND D( 1)='0' AND B( 5)='0' AND E( 5)='1' )then
          cVar1S29S41N025N062N027P048(0) <='1';
          else
          cVar1S29S41N025N062N027P048(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='1' AND E( 5)='1' )then
          cVar1S0S42P068P004P025P048nsss(0) <='1';
          else
          cVar1S0S42P068P004P025P048nsss(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='1' AND E( 5)='0' )then
          cVar1S1S42P068P004P025N048(0) <='1';
          else
          cVar1S1S42P068P004P025N048(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S2S42P068P004N025P040(0) <='1';
          else
          cVar1S2S42P068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S3S42P068P004N025P040(0) <='1';
          else
          cVar1S3S42P068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S4S42P068P004N025P040(0) <='1';
          else
          cVar1S4S42P068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='0' )then
          cVar1S5S42P068P004N025N040(0) <='1';
          else
          cVar1S5S42P068P004N025N040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='0' )then
          cVar1S6S42P068P004N025N040(0) <='1';
          else
          cVar1S6S42P068P004N025N040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='0' AND A( 3)='0' )then
          cVar1S7S42P068N004P055P013(0) <='1';
          else
          cVar1S7S42P068N004P055P013(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='0' AND A( 3)='0' )then
          cVar1S8S42P068N004P055P013(0) <='1';
          else
          cVar1S8S42P068N004P055P013(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='0' AND A( 3)='1' )then
          cVar1S9S42P068N004P055P013(0) <='1';
          else
          cVar1S9S42P068N004P055P013(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='0' AND A( 3)='1' )then
          cVar1S10S42P068N004P055P013(0) <='1';
          else
          cVar1S10S42P068N004P055P013(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='0' AND A( 3)='1' )then
          cVar1S11S42P068N004P055P013(0) <='1';
          else
          cVar1S11S42P068N004P055P013(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='1' AND D( 0)='0' )then
          cVar1S12S42P068N004P055P066(0) <='1';
          else
          cVar1S12S42P068N004P055P066(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='1' AND D( 0)='0' )then
          cVar1S13S42P068N004P055P066(0) <='1';
          else
          cVar1S13S42P068N004P055P066(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='1' AND D( 0)='0' )then
          cVar1S14S42P068N004P055P066(0) <='1';
          else
          cVar1S14S42P068N004P055P066(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='1' AND D( 0)='0' )then
          cVar1S15S42P068N004P055P066(0) <='1';
          else
          cVar1S15S42P068N004P055P066(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND D(11)='1' AND D( 0)='1' )then
          cVar1S16S42P068N004P055P066(0) <='1';
          else
          cVar1S16S42P068N004P055P066(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S17S42P068P015P061P069(0) <='1';
          else
          cVar1S17S42P068P015P061P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S18S42P068P015P061P069(0) <='1';
          else
          cVar1S18S42P068P015P061P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S19S42P068P015P061P069(0) <='1';
          else
          cVar1S19S42P068P015P061P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='1' AND E( 8)='1' )then
          cVar1S20S42P068P015P061P069(0) <='1';
          else
          cVar1S20S42P068P015P061P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='1' AND E( 8)='1' )then
          cVar1S21S42P068P015P061P069(0) <='1';
          else
          cVar1S21S42P068P015P061P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='0' AND B( 6)='1' )then
          cVar1S22S42P068P015N061P025nsss(0) <='1';
          else
          cVar1S22S42P068P015N061P025nsss(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='0' AND B( 6)='0' )then
          cVar1S23S42P068P015N061N025(0) <='1';
          else
          cVar1S23S42P068P015N061N025(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='0' AND B( 6)='0' )then
          cVar1S24S42P068P015N061N025(0) <='1';
          else
          cVar1S24S42P068P015N061N025(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='1' AND E(10)='0' AND B( 6)='0' )then
          cVar1S25S42P068P015N061N025(0) <='1';
          else
          cVar1S25S42P068P015N061N025(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='0' AND E( 8)='0' )then
          cVar1S26S42P068N015P059P069(0) <='1';
          else
          cVar1S26S42P068N015P059P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='0' AND E( 8)='0' )then
          cVar1S27S42P068N015P059P069(0) <='1';
          else
          cVar1S27S42P068N015P059P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='0' AND E( 8)='1' )then
          cVar1S28S42P068N015P059P069(0) <='1';
          else
          cVar1S28S42P068N015P059P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='0' AND E( 8)='1' )then
          cVar1S29S42P068N015P059P069(0) <='1';
          else
          cVar1S29S42P068N015P059P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='0' AND E( 8)='1' )then
          cVar1S30S42P068N015P059P069(0) <='1';
          else
          cVar1S30S42P068N015P059P069(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S31S42P068N015P059P032(0) <='1';
          else
          cVar1S31S42P068N015P059P032(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S32S42P068N015P059P032(0) <='1';
          else
          cVar1S32S42P068N015P059P032(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S33S42P068N015P059P032(0) <='1';
          else
          cVar1S33S42P068N015P059P032(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S34S42P068N015P059P032(0) <='1';
          else
          cVar1S34S42P068N015P059P032(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S35S42P068N015P059N032(0) <='1';
          else
          cVar1S35S42P068N015P059N032(0) <='0';
          end if;
        if(E( 0)='1' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S36S42P068N015P059N032(0) <='1';
          else
          cVar1S36S42P068N015P059N032(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S0S43P068P069P000P047(0) <='1';
          else
          cVar1S0S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S1S43P068P069P000P047(0) <='1';
          else
          cVar1S1S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S2S43P068P069P000P047(0) <='1';
          else
          cVar1S2S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S3S43P068P069P000P047(0) <='1';
          else
          cVar1S3S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S4S43P068P069P000P047(0) <='1';
          else
          cVar1S4S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S5S43P068P069P000P047(0) <='1';
          else
          cVar1S5S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S6S43P068P069P000P047(0) <='1';
          else
          cVar1S6S43P068P069P000P047(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='1' AND E( 1)='1' )then
          cVar1S7S43P068P069P000P064(0) <='1';
          else
          cVar1S7S43P068P069P000P064(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='1' AND E( 1)='0' )then
          cVar1S8S43P068P069P000N064(0) <='1';
          else
          cVar1S8S43P068P069P000N064(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='0' AND A(19)='1' AND E( 1)='0' )then
          cVar1S9S43P068P069P000N064(0) <='1';
          else
          cVar1S9S43P068P069P000N064(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='1' AND B( 7)='0' AND A( 0)='0' )then
          cVar1S10S43P068P069P023P019(0) <='1';
          else
          cVar1S10S43P068P069P023P019(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='1' AND B( 7)='0' AND A( 0)='0' )then
          cVar1S11S43P068P069P023P019(0) <='1';
          else
          cVar1S11S43P068P069P023P019(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='1' AND B( 7)='0' AND A( 0)='1' )then
          cVar1S12S43P068P069P023P019(0) <='1';
          else
          cVar1S12S43P068P069P023P019(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='1' AND B( 7)='0' AND A( 0)='1' )then
          cVar1S13S43P068P069P023P019(0) <='1';
          else
          cVar1S13S43P068P069P023P019(0) <='0';
          end if;
        if(E( 0)='1' AND E( 8)='1' AND B( 7)='0' AND A( 0)='1' )then
          cVar1S14S43P068P069P023P019(0) <='1';
          else
          cVar1S14S43P068P069P023P019(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='1' AND E( 5)='1' )then
          cVar1S15S43N068P004P025P048nsss(0) <='1';
          else
          cVar1S15S43N068P004P025P048nsss(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='1' AND E( 5)='0' )then
          cVar1S16S43N068P004P025N048(0) <='1';
          else
          cVar1S16S43N068P004P025N048(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S17S43N068P004N025P040(0) <='1';
          else
          cVar1S17S43N068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S18S43N068P004N025P040(0) <='1';
          else
          cVar1S18S43N068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='1' )then
          cVar1S19S43N068P004N025P040(0) <='1';
          else
          cVar1S19S43N068P004N025P040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='0' )then
          cVar1S20S43N068P004N025N040(0) <='1';
          else
          cVar1S20S43N068P004N025N040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='0' )then
          cVar1S21S43N068P004N025N040(0) <='1';
          else
          cVar1S21S43N068P004N025N040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='1' AND B( 6)='0' AND E( 7)='0' )then
          cVar1S22S43N068P004N025N040(0) <='1';
          else
          cVar1S22S43N068P004N025N040(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='1' AND E( 1)='1' )then
          cVar1S23S43N068N004P013P064(0) <='1';
          else
          cVar1S23S43N068N004P013P064(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='1' AND E( 1)='1' )then
          cVar1S24S43N068N004P013P064(0) <='1';
          else
          cVar1S24S43N068N004P013P064(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S25S43N068N004P013N064(0) <='1';
          else
          cVar1S25S43N068N004P013N064(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S26S43N068N004P013N064(0) <='1';
          else
          cVar1S26S43N068N004P013N064(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S27S43N068N004P013N064(0) <='1';
          else
          cVar1S27S43N068N004P013N064(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='1' )then
          cVar1S28S43N068N004N013P032(0) <='1';
          else
          cVar1S28S43N068N004N013P032(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='1' )then
          cVar1S29S43N068N004N013P032(0) <='1';
          else
          cVar1S29S43N068N004N013P032(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='1' )then
          cVar1S30S43N068N004N013P032(0) <='1';
          else
          cVar1S30S43N068N004N013P032(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='1' )then
          cVar1S31S43N068N004N013P032(0) <='1';
          else
          cVar1S31S43N068N004N013P032(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='0' )then
          cVar1S32S43N068N004N013N032(0) <='1';
          else
          cVar1S32S43N068N004N013N032(0) <='0';
          end if;
        if(E( 0)='0' AND A(17)='0' AND A( 3)='0' AND B(11)='0' )then
          cVar1S33S43N068N004N013N032(0) <='1';
          else
          cVar1S33S43N068N004N013N032(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar1S0S44P068P001P018P065(0) <='1';
          else
          cVar1S0S44P068P001P018P065(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S1S44P068P001P018N065(0) <='1';
          else
          cVar1S1S44P068P001P018N065(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S2S44P068P001P018N065(0) <='1';
          else
          cVar1S2S44P068P001P018N065(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S3S44P068P001P018N065(0) <='1';
          else
          cVar1S3S44P068P001P018N065(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S4S44P068P001P018N065(0) <='1';
          else
          cVar1S4S44P068P001P018N065(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='1' )then
          cVar1S5S44P068P001N018P046(0) <='1';
          else
          cVar1S5S44P068P001N018P046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='1' )then
          cVar1S6S44P068P001N018P046(0) <='1';
          else
          cVar1S6S44P068P001N018P046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='0' )then
          cVar1S7S44P068P001N018N046(0) <='1';
          else
          cVar1S7S44P068P001N018N046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='0' )then
          cVar1S8S44P068P001N018N046(0) <='1';
          else
          cVar1S8S44P068P001N018N046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='0' )then
          cVar1S9S44P068P001N018N046(0) <='1';
          else
          cVar1S9S44P068P001N018N046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='0' AND A(10)='0' AND D( 5)='0' )then
          cVar1S10S44P068P001N018N046(0) <='1';
          else
          cVar1S10S44P068P001N018N046(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='1' AND D( 3)='0' AND B( 9)='0' )then
          cVar1S11S44P068P001P054P036(0) <='1';
          else
          cVar1S11S44P068P001P054P036(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='1' AND D( 3)='0' AND B( 9)='0' )then
          cVar1S12S44P068P001P054P036(0) <='1';
          else
          cVar1S12S44P068P001P054P036(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='1' AND D( 3)='0' AND B( 9)='0' )then
          cVar1S13S44P068P001P054P036(0) <='1';
          else
          cVar1S13S44P068P001P054P036(0) <='0';
          end if;
        if(E( 0)='0' AND A( 9)='1' AND D( 3)='0' AND B( 9)='1' )then
          cVar1S14S44P068P001P054P036(0) <='1';
          else
          cVar1S14S44P068P001P054P036(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND E(11)='0' AND B( 7)='0' )then
          cVar1S15S44P068P067P057P023(0) <='1';
          else
          cVar1S15S44P068P067P057P023(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND E(11)='1' AND B(11)='1' )then
          cVar1S16S44P068P067P057P032nsss(0) <='1';
          else
          cVar1S16S44P068P067P057P032nsss(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND E(11)='1' AND B(11)='0' )then
          cVar1S17S44P068P067P057N032(0) <='1';
          else
          cVar1S17S44P068P067P057N032(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='1' AND E(11)='1' AND B(11)='0' )then
          cVar1S18S44P068P067P057N032(0) <='1';
          else
          cVar1S18S44P068P067P057N032(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='1' AND A(11)='0' )then
          cVar1S19S44P068N067P025P016(0) <='1';
          else
          cVar1S19S44P068N067P025P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='1' AND A(11)='0' )then
          cVar1S20S44P068N067P025P016(0) <='1';
          else
          cVar1S20S44P068N067P025P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='1' AND A(11)='0' )then
          cVar1S21S44P068N067P025P016(0) <='1';
          else
          cVar1S21S44P068N067P025P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='1' AND A(11)='1' )then
          cVar1S22S44P068N067P025P016(0) <='1';
          else
          cVar1S22S44P068N067P025P016(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='0' AND D( 0)='1' )then
          cVar1S23S44P068N067N025P066(0) <='1';
          else
          cVar1S23S44P068N067N025P066(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='0' AND D( 0)='0' )then
          cVar1S24S44P068N067N025N066(0) <='1';
          else
          cVar1S24S44P068N067N025N066(0) <='0';
          end if;
        if(E( 0)='1' AND D( 8)='0' AND B( 6)='0' AND D( 0)='0' )then
          cVar1S25S44P068N067N025N066(0) <='1';
          else
          cVar1S25S44P068N067N025N066(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='1' AND D( 8)='0' )then
          cVar1S0S45P014P068P016P067(0) <='1';
          else
          cVar1S0S45P014P068P016P067(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='1' AND D( 8)='0' )then
          cVar1S1S45P014P068P016P067(0) <='1';
          else
          cVar1S1S45P014P068P016P067(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='1' AND D( 8)='0' )then
          cVar1S2S45P014P068P016P067(0) <='1';
          else
          cVar1S2S45P014P068P016P067(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='1' AND D( 8)='1' )then
          cVar1S3S45P014P068P016P067(0) <='1';
          else
          cVar1S3S45P014P068P016P067(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='1' AND D( 8)='1' )then
          cVar1S4S45P014P068P016P067(0) <='1';
          else
          cVar1S4S45P014P068P016P067(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='0' )then
          cVar1S5S45P014P068N016P036(0) <='1';
          else
          cVar1S5S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='0' )then
          cVar1S6S45P014P068N016P036(0) <='1';
          else
          cVar1S6S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='0' )then
          cVar1S7S45P014P068N016P036(0) <='1';
          else
          cVar1S7S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='0' )then
          cVar1S8S45P014P068N016P036(0) <='1';
          else
          cVar1S8S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='1' )then
          cVar1S9S45P014P068N016P036(0) <='1';
          else
          cVar1S9S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='1' )then
          cVar1S10S45P014P068N016P036(0) <='1';
          else
          cVar1S10S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='0' AND A(11)='0' AND B( 9)='1' )then
          cVar1S11S45P014P068N016P036(0) <='1';
          else
          cVar1S11S45P014P068N016P036(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='0' AND E(14)='1' )then
          cVar1S12S45P014P068P067P045(0) <='1';
          else
          cVar1S12S45P014P068P067P045(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='0' AND E(14)='1' )then
          cVar1S13S45P014P068P067P045(0) <='1';
          else
          cVar1S13S45P014P068P067P045(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='0' AND E(14)='0' )then
          cVar1S14S45P014P068P067N045(0) <='1';
          else
          cVar1S14S45P014P068P067N045(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='0' AND E(14)='0' )then
          cVar1S15S45P014P068P067N045(0) <='1';
          else
          cVar1S15S45P014P068P067N045(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='0' AND E(14)='0' )then
          cVar1S16S45P014P068P067N045(0) <='1';
          else
          cVar1S16S45P014P068P067N045(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='1' AND B( 1)='1' )then
          cVar1S17S45P014P068P067P035(0) <='1';
          else
          cVar1S17S45P014P068P067P035(0) <='0';
          end if;
        if(A(12)='0' AND E( 0)='1' AND D( 8)='1' AND B( 1)='1' )then
          cVar1S18S45P014P068P067P035(0) <='1';
          else
          cVar1S18S45P014P068P067P035(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='0' AND B(10)='1' )then
          cVar1S19S45P014P015P021P034(0) <='1';
          else
          cVar1S19S45P014P015P021P034(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='0' AND B(10)='1' )then
          cVar1S20S45P014P015P021P034(0) <='1';
          else
          cVar1S20S45P014P015P021P034(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='0' AND B(10)='0' )then
          cVar1S21S45P014P015P021N034(0) <='1';
          else
          cVar1S21S45P014P015P021N034(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='0' AND B(10)='0' )then
          cVar1S22S45P014P015P021N034(0) <='1';
          else
          cVar1S22S45P014P015P021N034(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='0' AND B(10)='0' )then
          cVar1S23S45P014P015P021N034(0) <='1';
          else
          cVar1S23S45P014P015P021N034(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='1' AND B( 0)='1' )then
          cVar1S24S45P014P015P021P037(0) <='1';
          else
          cVar1S24S45P014P015P021P037(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='0' AND B( 8)='1' AND B( 0)='0' )then
          cVar1S25S45P014P015P021N037(0) <='1';
          else
          cVar1S25S45P014P015P021N037(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='1' AND A(10)='1' AND E(10)='1' )then
          cVar1S26S45P014P015P018P061(0) <='1';
          else
          cVar1S26S45P014P015P018P061(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='1' AND A(10)='1' AND E(10)='1' )then
          cVar1S27S45P014P015P018P061(0) <='1';
          else
          cVar1S27S45P014P015P018P061(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='1' AND A(10)='1' AND E(10)='0' )then
          cVar1S28S45P014P015P018N061(0) <='1';
          else
          cVar1S28S45P014P015P018N061(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='1' AND A(10)='1' AND E(10)='0' )then
          cVar1S29S45P014P015P018N061(0) <='1';
          else
          cVar1S29S45P014P015P018N061(0) <='0';
          end if;
        if(A(12)='1' AND A( 2)='1' AND A(10)='0' AND B(10)='1' )then
          cVar1S30S45P014P015N018P034(0) <='1';
          else
          cVar1S30S45P014P015N018P034(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='1' AND B( 8)='1' )then
          cVar1S0S46P016P038P021nsss(0) <='1';
          else
          cVar1S0S46P016P038P021nsss(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='1' AND B( 8)='0' AND A( 0)='0' )then
          cVar1S1S46P016P038N021P019(0) <='1';
          else
          cVar1S1S46P016P038N021P019(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='1' AND B( 8)='0' AND A( 0)='0' )then
          cVar1S2S46P016P038N021P019(0) <='1';
          else
          cVar1S2S46P016P038N021P019(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='1' AND B( 8)='0' AND A( 0)='0' )then
          cVar1S3S46P016P038N021P019(0) <='1';
          else
          cVar1S3S46P016P038N021P019(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='1' AND B( 8)='0' AND A( 0)='1' )then
          cVar1S4S46P016P038N021P019(0) <='1';
          else
          cVar1S4S46P016P038N021P019(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='0' )then
          cVar1S5S46P016N038P010P036(0) <='1';
          else
          cVar1S5S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='0' )then
          cVar1S6S46P016N038P010P036(0) <='1';
          else
          cVar1S6S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='0' )then
          cVar1S7S46P016N038P010P036(0) <='1';
          else
          cVar1S7S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='0' )then
          cVar1S8S46P016N038P010P036(0) <='1';
          else
          cVar1S8S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='1' )then
          cVar1S9S46P016N038P010P036(0) <='1';
          else
          cVar1S9S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='1' AND B( 9)='1' )then
          cVar1S10S46P016N038P010P036(0) <='1';
          else
          cVar1S10S46P016N038P010P036(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='1' )then
          cVar1S11S46P016N038N010P008(0) <='1';
          else
          cVar1S11S46P016N038N010P008(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='1' )then
          cVar1S12S46P016N038N010P008(0) <='1';
          else
          cVar1S12S46P016N038N010P008(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='1' )then
          cVar1S13S46P016N038N010P008(0) <='1';
          else
          cVar1S13S46P016N038N010P008(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='0' )then
          cVar1S14S46P016N038N010N008(0) <='1';
          else
          cVar1S14S46P016N038N010N008(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='0' )then
          cVar1S15S46P016N038N010N008(0) <='1';
          else
          cVar1S15S46P016N038N010N008(0) <='0';
          end if;
        if(A(11)='0' AND D( 7)='0' AND A(14)='0' AND A(15)='0' )then
          cVar1S16S46P016N038N010N008(0) <='1';
          else
          cVar1S16S46P016N038N010N008(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='1' AND E(13)='0' AND E( 3)='0' )then
          cVar1S17S46P016P032P049P056(0) <='1';
          else
          cVar1S17S46P016P032P049P056(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='1' AND E(13)='0' AND E( 3)='0' )then
          cVar1S18S46P016P032P049P056(0) <='1';
          else
          cVar1S18S46P016P032P049P056(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='1' AND E(13)='0' AND E( 3)='1' )then
          cVar1S19S46P016P032P049P056(0) <='1';
          else
          cVar1S19S46P016P032P049P056(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='0' )then
          cVar1S20S46P016N032P018P035(0) <='1';
          else
          cVar1S20S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='0' )then
          cVar1S21S46P016N032P018P035(0) <='1';
          else
          cVar1S21S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='0' )then
          cVar1S22S46P016N032P018P035(0) <='1';
          else
          cVar1S22S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='0' )then
          cVar1S23S46P016N032P018P035(0) <='1';
          else
          cVar1S23S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='1' )then
          cVar1S24S46P016N032P018P035(0) <='1';
          else
          cVar1S24S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='0' AND B( 1)='1' )then
          cVar1S25S46P016N032P018P035(0) <='1';
          else
          cVar1S25S46P016N032P018P035(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S26S46P016N032P018P058(0) <='1';
          else
          cVar1S26S46P016N032P018P058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S27S46P016N032P018P058(0) <='1';
          else
          cVar1S27S46P016N032P018P058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S28S46P016N032P018P058(0) <='1';
          else
          cVar1S28S46P016N032P018P058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S29S46P016N032P018N058(0) <='1';
          else
          cVar1S29S46P016N032P018N058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S30S46P016N032P018N058(0) <='1';
          else
          cVar1S30S46P016N032P018N058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S31S46P016N032P018N058(0) <='1';
          else
          cVar1S31S46P016N032P018N058(0) <='0';
          end if;
        if(A(11)='1' AND B(11)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S32S46P016N032P018N058(0) <='1';
          else
          cVar1S32S46P016N032P018N058(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='1' )then
          cVar1S0S47P067P016P064P047(0) <='1';
          else
          cVar1S0S47P067P016P064P047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='1' )then
          cVar1S1S47P067P016P064P047(0) <='1';
          else
          cVar1S1S47P067P016P064P047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='1' )then
          cVar1S2S47P067P016P064P047(0) <='1';
          else
          cVar1S2S47P067P016P064P047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='0' )then
          cVar1S3S47P067P016P064N047(0) <='1';
          else
          cVar1S3S47P067P016P064N047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='0' )then
          cVar1S4S47P067P016P064N047(0) <='1';
          else
          cVar1S4S47P067P016P064N047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='0' )then
          cVar1S5S47P067P016P064N047(0) <='1';
          else
          cVar1S5S47P067P016P064N047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='0' AND D(13)='0' )then
          cVar1S6S47P067P016P064N047(0) <='1';
          else
          cVar1S6S47P067P016P064N047(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S7S47P067P016P064P048(0) <='1';
          else
          cVar1S7S47P067P016P064P048(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S8S47P067P016P064P048(0) <='1';
          else
          cVar1S8S47P067P016P064P048(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S9S47P067P016P064P048(0) <='1';
          else
          cVar1S9S47P067P016P064P048(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='1' )then
          cVar1S10S47P067P016P064P048(0) <='1';
          else
          cVar1S10S47P067P016P064P048(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='1' )then
          cVar1S11S47P067P016P064P048(0) <='1';
          else
          cVar1S11S47P067P016P064P048(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='0' AND A(16)='0' )then
          cVar1S12S47P067P016P002P006(0) <='1';
          else
          cVar1S12S47P067P016P002P006(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='0' AND A(16)='0' )then
          cVar1S13S47P067P016P002P006(0) <='1';
          else
          cVar1S13S47P067P016P002P006(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='0' AND A(16)='1' )then
          cVar1S14S47P067P016P002P006(0) <='1';
          else
          cVar1S14S47P067P016P002P006(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='0' AND A(16)='1' )then
          cVar1S15S47P067P016P002P006(0) <='1';
          else
          cVar1S15S47P067P016P002P006(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='0' AND A(16)='1' )then
          cVar1S16S47P067P016P002P006(0) <='1';
          else
          cVar1S16S47P067P016P002P006(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='1' AND D( 4)='0' )then
          cVar1S17S47P067P016P002P050(0) <='1';
          else
          cVar1S17S47P067P016P002P050(0) <='0';
          end if;
        if(D( 8)='0' AND A(11)='1' AND A(18)='1' AND D( 4)='0' )then
          cVar1S18S47P067P016P002P050(0) <='1';
          else
          cVar1S18S47P067P016P002P050(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar1S19S47P067P062P058P033(0) <='1';
          else
          cVar1S19S47P067P062P058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar1S20S47P067P062P058P033(0) <='1';
          else
          cVar1S20S47P067P062P058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar1S21S47P067P062P058P033(0) <='1';
          else
          cVar1S21S47P067P062P058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='0' )then
          cVar1S22S47P067P062P058N033(0) <='1';
          else
          cVar1S22S47P067P062P058N033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='0' )then
          cVar1S23S47P067P062P058N033(0) <='1';
          else
          cVar1S23S47P067P062P058N033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='1' AND B( 2)='0' )then
          cVar1S24S47P067P062P058N033(0) <='1';
          else
          cVar1S24S47P067P062P058N033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S25S47P067P062N058P033(0) <='1';
          else
          cVar1S25S47P067P062N058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S26S47P067P062N058P033(0) <='1';
          else
          cVar1S26S47P067P062N058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S27S47P067P062N058P033(0) <='1';
          else
          cVar1S27S47P067P062N058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='0' AND B( 2)='1' )then
          cVar1S28S47P067P062N058P033(0) <='1';
          else
          cVar1S28S47P067P062N058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND D( 2)='0' AND B( 2)='1' )then
          cVar1S29S47P067P062N058P033(0) <='1';
          else
          cVar1S29S47P067P062N058P033(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='1' AND E( 6)='0' AND B( 1)='1' )then
          cVar1S30S47P067P062P044P035(0) <='1';
          else
          cVar1S30S47P067P062P044P035(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='1' AND E( 6)='0' AND B( 1)='1' )then
          cVar1S31S47P067P062P044P035(0) <='1';
          else
          cVar1S31S47P067P062P044P035(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='1' AND E( 6)='0' AND B( 1)='0' )then
          cVar1S32S47P067P062P044N035(0) <='1';
          else
          cVar1S32S47P067P062P044N035(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='1' AND E( 6)='0' AND B( 1)='0' )then
          cVar1S33S47P067P062P044N035(0) <='1';
          else
          cVar1S33S47P067P062P044N035(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='0' AND E(13)='1' )then
          cVar1S0S48P067P062P057P049(0) <='1';
          else
          cVar1S0S48P067P062P057P049(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='0' AND E(13)='1' )then
          cVar1S1S48P067P062P057P049(0) <='1';
          else
          cVar1S1S48P067P062P057P049(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='0' AND E(13)='0' )then
          cVar1S2S48P067P062P057N049(0) <='1';
          else
          cVar1S2S48P067P062P057N049(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='0' AND E(13)='0' )then
          cVar1S3S48P067P062P057N049(0) <='1';
          else
          cVar1S3S48P067P062P057N049(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='0' AND E(13)='0' )then
          cVar1S4S48P067P062P057N049(0) <='1';
          else
          cVar1S4S48P067P062P057N049(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='1' AND D(12)='0' )then
          cVar1S5S48P067P062P057P051(0) <='1';
          else
          cVar1S5S48P067P062P057P051(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='1' AND D(12)='0' )then
          cVar1S6S48P067P062P057P051(0) <='1';
          else
          cVar1S6S48P067P062P057P051(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='1' AND D(12)='0' )then
          cVar1S7S48P067P062P057P051(0) <='1';
          else
          cVar1S7S48P067P062P057P051(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='0' AND E(11)='1' AND D(12)='0' )then
          cVar1S8S48P067P062P057P051(0) <='1';
          else
          cVar1S8S48P067P062P057P051(0) <='0';
          end if;
        if(D( 8)='1' AND D( 1)='1' AND E( 6)='0' AND D( 6)='0' )then
          cVar1S9S48P067P062P044P042(0) <='1';
          else
          cVar1S9S48P067P062P044P042(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='1' AND D( 4)='1' )then
          cVar1S10S48N067P036P027P050(0) <='1';
          else
          cVar1S10S48N067P036P027P050(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='1' AND D( 4)='1' )then
          cVar1S11S48N067P036P027P050(0) <='1';
          else
          cVar1S11S48N067P036P027P050(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='1' AND D( 4)='1' )then
          cVar1S12S48N067P036P027P050(0) <='1';
          else
          cVar1S12S48N067P036P027P050(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='1' AND D( 4)='0' )then
          cVar1S13S48N067P036P027N050(0) <='1';
          else
          cVar1S13S48N067P036P027N050(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='1' AND D( 4)='0' )then
          cVar1S14S48N067P036P027N050(0) <='1';
          else
          cVar1S14S48N067P036P027N050(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='1' )then
          cVar1S15S48N067P036N027P016(0) <='1';
          else
          cVar1S15S48N067P036N027P016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='1' )then
          cVar1S16S48N067P036N027P016(0) <='1';
          else
          cVar1S16S48N067P036N027P016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='1' )then
          cVar1S17S48N067P036N027P016(0) <='1';
          else
          cVar1S17S48N067P036N027P016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='0' )then
          cVar1S18S48N067P036N027N016(0) <='1';
          else
          cVar1S18S48N067P036N027N016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='0' )then
          cVar1S19S48N067P036N027N016(0) <='1';
          else
          cVar1S19S48N067P036N027N016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='0' )then
          cVar1S20S48N067P036N027N016(0) <='1';
          else
          cVar1S20S48N067P036N027N016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='0' AND B( 5)='0' AND A(11)='0' )then
          cVar1S21S48N067P036N027N016(0) <='1';
          else
          cVar1S21S48N067P036N027N016(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='0' AND D(14)='1' )then
          cVar1S22S48N067P036P005P043(0) <='1';
          else
          cVar1S22S48N067P036P005P043(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='0' AND D(14)='1' )then
          cVar1S23S48N067P036P005P043(0) <='1';
          else
          cVar1S23S48N067P036P005P043(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='0' AND D(14)='0' )then
          cVar1S24S48N067P036P005N043(0) <='1';
          else
          cVar1S24S48N067P036P005N043(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='1' AND B(11)='1' )then
          cVar1S25S48N067P036P005P032nsss(0) <='1';
          else
          cVar1S25S48N067P036P005P032nsss(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='1' AND B(11)='0' )then
          cVar1S26S48N067P036P005N032(0) <='1';
          else
          cVar1S26S48N067P036P005N032(0) <='0';
          end if;
        if(D( 8)='0' AND B( 9)='1' AND A( 7)='1' AND B(11)='0' )then
          cVar1S27S48N067P036P005N032(0) <='1';
          else
          cVar1S27S48N067P036P005N032(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S0S49P036P011P010P013(0) <='1';
          else
          cVar1S0S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S1S49P036P011P010P013(0) <='1';
          else
          cVar1S1S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S2S49P036P011P010P013(0) <='1';
          else
          cVar1S2S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar1S3S49P036P011P010P013(0) <='1';
          else
          cVar1S3S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar1S4S49P036P011P010P013(0) <='1';
          else
          cVar1S4S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar1S5S49P036P011P010P013(0) <='1';
          else
          cVar1S5S49P036P011P010P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='1' AND D( 6)='1' )then
          cVar1S6S49P036P011P010P042nsss(0) <='1';
          else
          cVar1S6S49P036P011P010P042nsss(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='1' AND D( 6)='0' )then
          cVar1S7S49P036P011P010N042(0) <='1';
          else
          cVar1S7S49P036P011P010N042(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND A(14)='1' AND D( 6)='0' )then
          cVar1S8S49P036P011P010N042(0) <='1';
          else
          cVar1S8S49P036P011P010N042(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='1' AND D(15)='1' )then
          cVar1S9S49P036N011P005P039(0) <='1';
          else
          cVar1S9S49P036N011P005P039(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='1' AND D(15)='1' )then
          cVar1S10S49P036N011P005P039(0) <='1';
          else
          cVar1S10S49P036N011P005P039(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='1' AND D(15)='1' )then
          cVar1S11S49P036N011P005P039(0) <='1';
          else
          cVar1S11S49P036N011P005P039(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='1' AND D(15)='0' )then
          cVar1S12S49P036N011P005N039(0) <='1';
          else
          cVar1S12S49P036N011P005N039(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='1' AND D(15)='0' )then
          cVar1S13S49P036N011P005N039(0) <='1';
          else
          cVar1S13S49P036N011P005N039(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='0' )then
          cVar1S14S49P036N011N005P016(0) <='1';
          else
          cVar1S14S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='0' )then
          cVar1S15S49P036N011N005P016(0) <='1';
          else
          cVar1S15S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='0' )then
          cVar1S16S49P036N011N005P016(0) <='1';
          else
          cVar1S16S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='0' )then
          cVar1S17S49P036N011N005P016(0) <='1';
          else
          cVar1S17S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='1' )then
          cVar1S18S49P036N011N005P016(0) <='1';
          else
          cVar1S18S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='1' )then
          cVar1S19S49P036N011N005P016(0) <='1';
          else
          cVar1S19S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A( 7)='0' AND A(11)='1' )then
          cVar1S20S49P036N011N005P016(0) <='1';
          else
          cVar1S20S49P036N011N005P016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='1' )then
          cVar1S21S49P036P043P022nsss(0) <='1';
          else
          cVar1S21S49P036P043P022nsss(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND A( 2)='0' )then
          cVar1S22S49P036P043N022P015(0) <='1';
          else
          cVar1S22S49P036P043N022P015(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND A( 2)='0' )then
          cVar1S23S49P036P043N022P015(0) <='1';
          else
          cVar1S23S49P036P043N022P015(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND A( 2)='0' )then
          cVar1S24S49P036P043N022P015(0) <='1';
          else
          cVar1S24S49P036P043N022P015(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND A(11)='1' )then
          cVar1S25S49P036N043P045P016(0) <='1';
          else
          cVar1S25S49P036N043P045P016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND A(11)='1' )then
          cVar1S26S49P036N043P045P016(0) <='1';
          else
          cVar1S26S49P036N043P045P016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND A(11)='0' )then
          cVar1S27S49P036N043P045N016(0) <='1';
          else
          cVar1S27S49P036N043P045N016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND A(11)='0' )then
          cVar1S28S49P036N043P045N016(0) <='1';
          else
          cVar1S28S49P036N043P045N016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND A(11)='0' )then
          cVar1S29S49P036N043P045N016(0) <='1';
          else
          cVar1S29S49P036N043P045N016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='1' AND A(11)='1' )then
          cVar1S30S49P036N043P045P016(0) <='1';
          else
          cVar1S30S49P036N043P045P016(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='1' )then
          cVar1S0S50P036P033P015P038(0) <='1';
          else
          cVar1S0S50P036P033P015P038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='1' )then
          cVar1S1S50P036P033P015P038(0) <='1';
          else
          cVar1S1S50P036P033P015P038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='1' )then
          cVar1S2S50P036P033P015P038(0) <='1';
          else
          cVar1S2S50P036P033P015P038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='0' )then
          cVar1S3S50P036P033P015N038(0) <='1';
          else
          cVar1S3S50P036P033P015N038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='0' )then
          cVar1S4S50P036P033P015N038(0) <='1';
          else
          cVar1S4S50P036P033P015N038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='0' )then
          cVar1S5S50P036P033P015N038(0) <='1';
          else
          cVar1S5S50P036P033P015N038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='0' AND D( 7)='0' )then
          cVar1S6S50P036P033P015N038(0) <='1';
          else
          cVar1S6S50P036P033P015N038(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='0' )then
          cVar1S7S50P036P033P015P049(0) <='1';
          else
          cVar1S7S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='0' )then
          cVar1S8S50P036P033P015P049(0) <='1';
          else
          cVar1S8S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='0' )then
          cVar1S9S50P036P033P015P049(0) <='1';
          else
          cVar1S9S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='0' )then
          cVar1S10S50P036P033P015P049(0) <='1';
          else
          cVar1S10S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='1' )then
          cVar1S11S50P036P033P015P049(0) <='1';
          else
          cVar1S11S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='0' AND A( 2)='1' AND E(13)='1' )then
          cVar1S12S50P036P033P015P049(0) <='1';
          else
          cVar1S12S50P036P033P015P049(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='0' AND A( 9)='0' )then
          cVar1S13S50P036P033P026P001(0) <='1';
          else
          cVar1S13S50P036P033P026P001(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='0' AND A( 9)='0' )then
          cVar1S14S50P036P033P026P001(0) <='1';
          else
          cVar1S14S50P036P033P026P001(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='0' AND A( 9)='0' )then
          cVar1S15S50P036P033P026P001(0) <='1';
          else
          cVar1S15S50P036P033P026P001(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='0' AND A( 9)='1' )then
          cVar1S16S50P036P033P026P001(0) <='1';
          else
          cVar1S16S50P036P033P026P001(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='1' AND D(13)='1' )then
          cVar1S17S50P036P033P026P047nsss(0) <='1';
          else
          cVar1S17S50P036P033P026P047nsss(0) <='0';
          end if;
        if(B( 9)='0' AND B( 2)='1' AND B(14)='1' AND D(13)='0' )then
          cVar1S18S50P036P033P026N047(0) <='1';
          else
          cVar1S18S50P036P033P026N047(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='1' AND A(10)='1' )then
          cVar1S19S50P036P068P065P018(0) <='1';
          else
          cVar1S19S50P036P068P065P018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='1' AND A(10)='0' )then
          cVar1S20S50P036P068P065N018(0) <='1';
          else
          cVar1S20S50P036P068P065N018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='1' AND A(10)='0' )then
          cVar1S21S50P036P068P065N018(0) <='1';
          else
          cVar1S21S50P036P068P065N018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='1' AND A(10)='0' )then
          cVar1S22S50P036P068P065N018(0) <='1';
          else
          cVar1S22S50P036P068P065N018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='0' AND A(10)='0' )then
          cVar1S23S50P036P068N065P018(0) <='1';
          else
          cVar1S23S50P036P068N065P018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='0' AND A(10)='0' )then
          cVar1S24S50P036P068N065P018(0) <='1';
          else
          cVar1S24S50P036P068N065P018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='0' AND A(10)='1' )then
          cVar1S25S50P036P068N065P018(0) <='1';
          else
          cVar1S25S50P036P068N065P018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='0' AND E( 9)='0' AND A(10)='1' )then
          cVar1S26S50P036P068N065P018(0) <='1';
          else
          cVar1S26S50P036P068N065P018(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='1' AND B( 6)='1' )then
          cVar1S27S50P036P068P019P025nsss(0) <='1';
          else
          cVar1S27S50P036P068P019P025nsss(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='1' AND B( 6)='0' )then
          cVar1S28S50P036P068P019N025(0) <='1';
          else
          cVar1S28S50P036P068P019N025(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='1' AND B( 6)='0' )then
          cVar1S29S50P036P068P019N025(0) <='1';
          else
          cVar1S29S50P036P068P019N025(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S30S50P036P068N019P066(0) <='1';
          else
          cVar1S30S50P036P068N019P066(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S31S50P036P068N019P066(0) <='1';
          else
          cVar1S31S50P036P068N019P066(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S32S50P036P068N019P066(0) <='1';
          else
          cVar1S32S50P036P068N019P066(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S33S50P036P068N019P066(0) <='1';
          else
          cVar1S33S50P036P068N019P066(0) <='0';
          end if;
        if(B( 9)='1' AND E( 0)='1' AND A( 0)='0' AND D( 0)='0' )then
          cVar1S34S50P036P068N019N066(0) <='1';
          else
          cVar1S34S50P036P068N019N066(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='1' AND B( 1)='0' )then
          cVar1S0S51P033P015P032P035(0) <='1';
          else
          cVar1S0S51P033P015P032P035(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='1' AND B( 1)='0' )then
          cVar1S1S51P033P015P032P035(0) <='1';
          else
          cVar1S1S51P033P015P032P035(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='1' AND B( 1)='1' )then
          cVar1S2S51P033P015P032P035(0) <='1';
          else
          cVar1S2S51P033P015P032P035(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='1' AND B( 1)='1' )then
          cVar1S3S51P033P015P032P035(0) <='1';
          else
          cVar1S3S51P033P015P032P035(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='1' AND B( 1)='1' )then
          cVar1S4S51P033P015P032P035(0) <='1';
          else
          cVar1S4S51P033P015P032P035(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='0' AND A( 1)='0' )then
          cVar1S5S51P033P015N032P017(0) <='1';
          else
          cVar1S5S51P033P015N032P017(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='0' AND A( 1)='0' )then
          cVar1S6S51P033P015N032P017(0) <='1';
          else
          cVar1S6S51P033P015N032P017(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='0' AND A( 1)='1' )then
          cVar1S7S51P033P015N032P017(0) <='1';
          else
          cVar1S7S51P033P015N032P017(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='0' AND A( 1)='1' )then
          cVar1S8S51P033P015N032P017(0) <='1';
          else
          cVar1S8S51P033P015N032P017(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='1' AND B(11)='0' AND A( 1)='1' )then
          cVar1S9S51P033P015N032P017(0) <='1';
          else
          cVar1S9S51P033P015N032P017(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S10S51P033N015P059P049(0) <='1';
          else
          cVar1S10S51P033N015P059P049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S11S51P033N015P059P049(0) <='1';
          else
          cVar1S11S51P033N015P059P049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S12S51P033N015P059P049(0) <='1';
          else
          cVar1S12S51P033N015P059P049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S13S51P033N015P059P049(0) <='1';
          else
          cVar1S13S51P033N015P059P049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='0' )then
          cVar1S14S51P033N015P059N049(0) <='1';
          else
          cVar1S14S51P033N015P059N049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='0' )then
          cVar1S15S51P033N015P059N049(0) <='1';
          else
          cVar1S15S51P033N015P059N049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='0' AND E(13)='0' )then
          cVar1S16S51P033N015P059N049(0) <='1';
          else
          cVar1S16S51P033N015P059N049(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S17S51P033N015P059P032(0) <='1';
          else
          cVar1S17S51P033N015P059P032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S18S51P033N015P059P032(0) <='1';
          else
          cVar1S18S51P033N015P059P032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='1' )then
          cVar1S19S51P033N015P059P032(0) <='1';
          else
          cVar1S19S51P033N015P059P032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S20S51P033N015P059N032(0) <='1';
          else
          cVar1S20S51P033N015P059N032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S21S51P033N015P059N032(0) <='1';
          else
          cVar1S21S51P033N015P059N032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S22S51P033N015P059N032(0) <='1';
          else
          cVar1S22S51P033N015P059N032(0) <='0';
          end if;
        if(B( 2)='0' AND A( 2)='0' AND D(10)='1' AND B(11)='0' )then
          cVar1S23S51P033N015P059N032(0) <='1';
          else
          cVar1S23S51P033N015P059N032(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='1' AND A(11)='0' AND E( 2)='0' )then
          cVar1S24S51P033P056P016P060(0) <='1';
          else
          cVar1S24S51P033P056P016P060(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='1' AND A(11)='0' AND E( 2)='0' )then
          cVar1S25S51P033P056P016P060(0) <='1';
          else
          cVar1S25S51P033P056P016P060(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='1' AND A(11)='0' AND E( 2)='1' )then
          cVar1S26S51P033P056P016P060(0) <='1';
          else
          cVar1S26S51P033P056P016P060(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='1' AND A(11)='0' AND E( 2)='1' )then
          cVar1S27S51P033P056P016P060(0) <='1';
          else
          cVar1S27S51P033P056P016P060(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='1' AND A(11)='1' AND D( 2)='1' )then
          cVar1S28S51P033P056P016P058(0) <='1';
          else
          cVar1S28S51P033P056P016P058(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='0' AND A(16)='1' AND D( 6)='1' )then
          cVar1S29S51P033N056P006P042nsss(0) <='1';
          else
          cVar1S29S51P033N056P006P042nsss(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='0' AND A(16)='1' AND D( 6)='0' )then
          cVar1S30S51P033N056P006N042(0) <='1';
          else
          cVar1S30S51P033N056P006N042(0) <='0';
          end if;
        if(B( 2)='1' AND E( 3)='0' AND A(16)='1' AND D( 6)='0' )then
          cVar1S31S51P033N056P006N042(0) <='1';
          else
          cVar1S31S51P033N056P006N042(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='1' AND B( 0)='1' )then
          cVar1S0S52P006P017P064P037(0) <='1';
          else
          cVar1S0S52P006P017P064P037(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='1' AND B( 0)='1' )then
          cVar1S1S52P006P017P064P037(0) <='1';
          else
          cVar1S1S52P006P017P064P037(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='1' AND B( 0)='0' )then
          cVar1S2S52P006P017P064N037(0) <='1';
          else
          cVar1S2S52P006P017P064N037(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='1' AND B( 0)='0' )then
          cVar1S3S52P006P017P064N037(0) <='1';
          else
          cVar1S3S52P006P017P064N037(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='1' AND B( 0)='0' )then
          cVar1S4S52P006P017P064N037(0) <='1';
          else
          cVar1S4S52P006P017P064N037(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='0' AND A( 7)='0' )then
          cVar1S5S52P006P017N064P005(0) <='1';
          else
          cVar1S5S52P006P017N064P005(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='0' AND A( 7)='0' )then
          cVar1S6S52P006P017N064P005(0) <='1';
          else
          cVar1S6S52P006P017N064P005(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='0' AND A( 7)='0' )then
          cVar1S7S52P006P017N064P005(0) <='1';
          else
          cVar1S7S52P006P017N064P005(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='0' AND A( 7)='1' )then
          cVar1S8S52P006P017N064P005(0) <='1';
          else
          cVar1S8S52P006P017N064P005(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='1' AND E( 1)='0' AND A( 7)='1' )then
          cVar1S9S52P006P017N064P005(0) <='1';
          else
          cVar1S9S52P006P017N064P005(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='0' )then
          cVar1S10S52P006N017P059P044(0) <='1';
          else
          cVar1S10S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='0' )then
          cVar1S11S52P006N017P059P044(0) <='1';
          else
          cVar1S11S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='0' )then
          cVar1S12S52P006N017P059P044(0) <='1';
          else
          cVar1S12S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='0' )then
          cVar1S13S52P006N017P059P044(0) <='1';
          else
          cVar1S13S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='1' )then
          cVar1S14S52P006N017P059P044(0) <='1';
          else
          cVar1S14S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='0' AND E( 6)='1' )then
          cVar1S15S52P006N017P059P044(0) <='1';
          else
          cVar1S15S52P006N017P059P044(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='1' AND E( 2)='0' )then
          cVar1S16S52P006N017P059P060(0) <='1';
          else
          cVar1S16S52P006N017P059P060(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='1' AND E( 2)='0' )then
          cVar1S17S52P006N017P059P060(0) <='1';
          else
          cVar1S17S52P006N017P059P060(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='1' AND E( 2)='1' )then
          cVar1S18S52P006N017P059P060(0) <='1';
          else
          cVar1S18S52P006N017P059P060(0) <='0';
          end if;
        if(A(16)='0' AND A( 1)='0' AND D(10)='1' AND E( 2)='1' )then
          cVar1S19S52P006N017P059P060(0) <='1';
          else
          cVar1S19S52P006N017P059P060(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='1' AND E( 6)='1' )then
          cVar1S20S52P006P042P044nsss(0) <='1';
          else
          cVar1S20S52P006P042P044nsss(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='1' AND E( 6)='0' AND A( 0)='1' )then
          cVar1S21S52P006P042N044P019nsss(0) <='1';
          else
          cVar1S21S52P006P042N044P019nsss(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='1' AND E( 1)='0' )then
          cVar1S22S52P006N042P047P064(0) <='1';
          else
          cVar1S22S52P006N042P047P064(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='1' AND E( 1)='0' )then
          cVar1S23S52P006N042P047P064(0) <='1';
          else
          cVar1S23S52P006N042P047P064(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='1' AND E( 1)='0' )then
          cVar1S24S52P006N042P047P064(0) <='1';
          else
          cVar1S24S52P006N042P047P064(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='0' AND D(14)='1' )then
          cVar1S25S52P006N042N047P043(0) <='1';
          else
          cVar1S25S52P006N042N047P043(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='0' AND D(14)='0' )then
          cVar1S26S52P006N042N047N043(0) <='1';
          else
          cVar1S26S52P006N042N047N043(0) <='0';
          end if;
        if(A(16)='1' AND D( 6)='0' AND D(13)='0' AND D(14)='0' )then
          cVar1S27S52P006N042N047N043(0) <='1';
          else
          cVar1S27S52P006N042N047N043(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='0' )then
          cVar1S0S53P016P059P017P061(0) <='1';
          else
          cVar1S0S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='0' )then
          cVar1S1S53P016P059P017P061(0) <='1';
          else
          cVar1S1S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='0' )then
          cVar1S2S53P016P059P017P061(0) <='1';
          else
          cVar1S2S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='0' )then
          cVar1S3S53P016P059P017P061(0) <='1';
          else
          cVar1S3S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='1' )then
          cVar1S4S53P016P059P017P061(0) <='1';
          else
          cVar1S4S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='1' )then
          cVar1S5S53P016P059P017P061(0) <='1';
          else
          cVar1S5S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='0' AND E(10)='1' )then
          cVar1S6S53P016P059P017P061(0) <='1';
          else
          cVar1S6S53P016P059P017P061(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar1S7S53P016P059P017P015(0) <='1';
          else
          cVar1S7S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar1S8S53P016P059P017P015(0) <='1';
          else
          cVar1S8S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar1S9S53P016P059P017P015(0) <='1';
          else
          cVar1S9S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar1S10S53P016P059P017P015(0) <='1';
          else
          cVar1S10S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='1' )then
          cVar1S11S53P016P059P017P015(0) <='1';
          else
          cVar1S11S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='1' )then
          cVar1S12S53P016P059P017P015(0) <='1';
          else
          cVar1S12S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='1' )then
          cVar1S13S53P016P059P017P015(0) <='1';
          else
          cVar1S13S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='0' AND A( 1)='1' AND A( 2)='1' )then
          cVar1S14S53P016P059P017P015(0) <='1';
          else
          cVar1S14S53P016P059P017P015(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='1' )then
          cVar1S15S53P016P059P015P019(0) <='1';
          else
          cVar1S15S53P016P059P015P019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='1' )then
          cVar1S16S53P016P059P015P019(0) <='1';
          else
          cVar1S16S53P016P059P015P019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='1' )then
          cVar1S17S53P016P059P015P019(0) <='1';
          else
          cVar1S17S53P016P059P015P019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='0' )then
          cVar1S18S53P016P059P015N019(0) <='1';
          else
          cVar1S18S53P016P059P015N019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='0' )then
          cVar1S19S53P016P059P015N019(0) <='1';
          else
          cVar1S19S53P016P059P015N019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='1' AND A( 0)='0' )then
          cVar1S20S53P016P059P015N019(0) <='1';
          else
          cVar1S20S53P016P059P015N019(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='0' AND D( 0)='0' )then
          cVar1S21S53P016P059N015P066(0) <='1';
          else
          cVar1S21S53P016P059N015P066(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='0' AND D( 0)='0' )then
          cVar1S22S53P016P059N015P066(0) <='1';
          else
          cVar1S22S53P016P059N015P066(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='0' AND D( 0)='0' )then
          cVar1S23S53P016P059N015P066(0) <='1';
          else
          cVar1S23S53P016P059N015P066(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='0' AND D( 0)='0' )then
          cVar1S24S53P016P059N015P066(0) <='1';
          else
          cVar1S24S53P016P059N015P066(0) <='0';
          end if;
        if(A(11)='0' AND D(10)='1' AND A( 2)='0' AND D( 0)='1' )then
          cVar1S25S53P016P059N015P066(0) <='1';
          else
          cVar1S25S53P016P059N015P066(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='0' AND B( 8)='0' )then
          cVar1S26S53P016P038P002P021(0) <='1';
          else
          cVar1S26S53P016P038P002P021(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='0' AND B( 8)='0' )then
          cVar1S27S53P016P038P002P021(0) <='1';
          else
          cVar1S27S53P016P038P002P021(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='0' AND B( 8)='0' )then
          cVar1S28S53P016P038P002P021(0) <='1';
          else
          cVar1S28S53P016P038P002P021(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='0' AND B( 8)='0' )then
          cVar1S29S53P016P038P002P021(0) <='1';
          else
          cVar1S29S53P016P038P002P021(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='0' AND B( 8)='1' )then
          cVar1S30S53P016P038P002P021(0) <='1';
          else
          cVar1S30S53P016P038P002P021(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='1' AND A( 0)='1' )then
          cVar1S31S53P016P038P002P019(0) <='1';
          else
          cVar1S31S53P016P038P002P019(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='1' AND A( 0)='1' )then
          cVar1S32S53P016P038P002P019(0) <='1';
          else
          cVar1S32S53P016P038P002P019(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='1' AND A( 0)='0' )then
          cVar1S33S53P016P038P002N019(0) <='1';
          else
          cVar1S33S53P016P038P002N019(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND A(18)='1' AND A( 0)='0' )then
          cVar1S34S53P016P038P002N019(0) <='1';
          else
          cVar1S34S53P016P038P002N019(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='1' AND B( 2)='0' AND E( 1)='0' )then
          cVar1S35S53P016P038P033P064(0) <='1';
          else
          cVar1S35S53P016P038P033P064(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='1' AND B( 2)='0' AND E( 1)='0' )then
          cVar1S36S53P016P038P033P064(0) <='1';
          else
          cVar1S36S53P016P038P033P064(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='1' AND B( 2)='0' AND E( 1)='0' )then
          cVar1S37S53P016P038P033P064(0) <='1';
          else
          cVar1S37S53P016P038P033P064(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='0' AND A(18)='0' )then
          cVar1S0S54P037P016P038P002(0) <='1';
          else
          cVar1S0S54P037P016P038P002(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='0' AND A(18)='0' )then
          cVar1S1S54P037P016P038P002(0) <='1';
          else
          cVar1S1S54P037P016P038P002(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='0' AND A(18)='0' )then
          cVar1S2S54P037P016P038P002(0) <='1';
          else
          cVar1S2S54P037P016P038P002(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='0' AND A(18)='1' )then
          cVar1S3S54P037P016P038P002(0) <='1';
          else
          cVar1S3S54P037P016P038P002(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='0' AND A(18)='1' )then
          cVar1S4S54P037P016P038P002(0) <='1';
          else
          cVar1S4S54P037P016P038P002(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='1' AND B( 2)='0' )then
          cVar1S5S54P037P016P038P033(0) <='1';
          else
          cVar1S5S54P037P016P038P033(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='1' AND D( 7)='1' AND B( 2)='0' )then
          cVar1S6S54P037P016P038P033(0) <='1';
          else
          cVar1S6S54P037P016P038P033(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='1' AND D( 5)='0' )then
          cVar1S7S54P037N016P050P046(0) <='1';
          else
          cVar1S7S54P037N016P050P046(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='1' AND D( 5)='0' )then
          cVar1S8S54P037N016P050P046(0) <='1';
          else
          cVar1S8S54P037N016P050P046(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='1' AND D( 5)='1' )then
          cVar1S9S54P037N016P050P046(0) <='1';
          else
          cVar1S9S54P037N016P050P046(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='0' AND D(15)='1' )then
          cVar1S10S54P037N016N050P039(0) <='1';
          else
          cVar1S10S54P037N016N050P039(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='0' AND D(15)='1' )then
          cVar1S11S54P037N016N050P039(0) <='1';
          else
          cVar1S11S54P037N016N050P039(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='0' AND D(15)='1' )then
          cVar1S12S54P037N016N050P039(0) <='1';
          else
          cVar1S12S54P037N016N050P039(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='0' AND D(15)='0' )then
          cVar1S13S54P037N016N050N039(0) <='1';
          else
          cVar1S13S54P037N016N050N039(0) <='0';
          end if;
        if(B( 0)='0' AND A(11)='0' AND D( 4)='0' AND D(15)='0' )then
          cVar1S14S54P037N016N050N039(0) <='1';
          else
          cVar1S14S54P037N016N050N039(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='0' )then
          cVar1S15S54P037P018P060P031(0) <='1';
          else
          cVar1S15S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='0' )then
          cVar1S16S54P037P018P060P031(0) <='1';
          else
          cVar1S16S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='0' )then
          cVar1S17S54P037P018P060P031(0) <='1';
          else
          cVar1S17S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='1' )then
          cVar1S18S54P037P018P060P031(0) <='1';
          else
          cVar1S18S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='1' )then
          cVar1S19S54P037P018P060P031(0) <='1';
          else
          cVar1S19S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='0' AND B( 3)='1' )then
          cVar1S20S54P037P018P060P031(0) <='1';
          else
          cVar1S20S54P037P018P060P031(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='1' AND D( 0)='1' )then
          cVar1S21S54P037P018P060P066(0) <='1';
          else
          cVar1S21S54P037P018P060P066(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='1' AND D( 0)='1' )then
          cVar1S22S54P037P018P060P066(0) <='1';
          else
          cVar1S22S54P037P018P060P066(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='1' AND D( 0)='1' )then
          cVar1S23S54P037P018P060P066(0) <='1';
          else
          cVar1S23S54P037P018P060P066(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='1' AND E( 2)='1' AND D( 0)='0' )then
          cVar1S24S54P037P018P060N066(0) <='1';
          else
          cVar1S24S54P037P018P060N066(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='0' )then
          cVar1S25S54P037N018P017P065(0) <='1';
          else
          cVar1S25S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='0' )then
          cVar1S26S54P037N018P017P065(0) <='1';
          else
          cVar1S26S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='0' )then
          cVar1S27S54P037N018P017P065(0) <='1';
          else
          cVar1S27S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='1' )then
          cVar1S28S54P037N018P017P065(0) <='1';
          else
          cVar1S28S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='1' )then
          cVar1S29S54P037N018P017P065(0) <='1';
          else
          cVar1S29S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='1' )then
          cVar1S30S54P037N018P017P065(0) <='1';
          else
          cVar1S30S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='1' AND E( 9)='1' )then
          cVar1S31S54P037N018P017P065(0) <='1';
          else
          cVar1S31S54P037N018P017P065(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='0' AND E( 1)='0' )then
          cVar1S32S54P037N018N017P064(0) <='1';
          else
          cVar1S32S54P037N018N017P064(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='0' AND E( 1)='0' )then
          cVar1S33S54P037N018N017P064(0) <='1';
          else
          cVar1S33S54P037N018N017P064(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='0' AND E( 1)='1' )then
          cVar1S34S54P037N018N017P064(0) <='1';
          else
          cVar1S34S54P037N018N017P064(0) <='0';
          end if;
        if(B( 0)='1' AND A(10)='0' AND A( 1)='0' AND E( 1)='1' )then
          cVar1S35S54P037N018N017P064(0) <='1';
          else
          cVar1S35S54P037N018N017P064(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='0' AND A( 9)='0' )then
          cVar1S0S55P016P037P062P001(0) <='1';
          else
          cVar1S0S55P016P037P062P001(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='0' AND A( 9)='0' )then
          cVar1S1S55P016P037P062P001(0) <='1';
          else
          cVar1S1S55P016P037P062P001(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='0' AND A( 9)='0' )then
          cVar1S2S55P016P037P062P001(0) <='1';
          else
          cVar1S2S55P016P037P062P001(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='0' AND A( 9)='0' )then
          cVar1S3S55P016P037P062P001(0) <='1';
          else
          cVar1S3S55P016P037P062P001(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='0' AND A( 9)='1' )then
          cVar1S4S55P016P037P062P001(0) <='1';
          else
          cVar1S4S55P016P037P062P001(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='1' AND D(13)='0' )then
          cVar1S5S55P016P037P062P047(0) <='1';
          else
          cVar1S5S55P016P037P062P047(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='1' AND D(13)='0' )then
          cVar1S6S55P016P037P062P047(0) <='1';
          else
          cVar1S6S55P016P037P062P047(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='0' AND D( 1)='1' AND D(13)='1' )then
          cVar1S7S55P016P037P062P047(0) <='1';
          else
          cVar1S7S55P016P037P062P047(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='1' AND A(15)='1' )then
          cVar1S8S55P016P037P017P008nsss(0) <='1';
          else
          cVar1S8S55P016P037P017P008nsss(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='1' AND A(15)='0' )then
          cVar1S9S55P016P037P017N008(0) <='1';
          else
          cVar1S9S55P016P037P017N008(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='1' AND A(15)='0' )then
          cVar1S10S55P016P037P017N008(0) <='1';
          else
          cVar1S10S55P016P037P017N008(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='1' AND A(15)='0' )then
          cVar1S11S55P016P037P017N008(0) <='1';
          else
          cVar1S11S55P016P037P017N008(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='1' AND A(15)='0' )then
          cVar1S12S55P016P037P017N008(0) <='1';
          else
          cVar1S12S55P016P037P017N008(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='0' AND D( 8)='1' )then
          cVar1S13S55P016P037N017P067(0) <='1';
          else
          cVar1S13S55P016P037N017P067(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='0' AND D( 8)='1' )then
          cVar1S14S55P016P037N017P067(0) <='1';
          else
          cVar1S14S55P016P037N017P067(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='0' AND D( 8)='0' )then
          cVar1S15S55P016P037N017N067(0) <='1';
          else
          cVar1S15S55P016P037N017N067(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='0' AND D( 8)='0' )then
          cVar1S16S55P016P037N017N067(0) <='1';
          else
          cVar1S16S55P016P037N017N067(0) <='0';
          end if;
        if(A(11)='0' AND B( 0)='1' AND A( 1)='0' AND D( 8)='0' )then
          cVar1S17S55P016P037N017N067(0) <='1';
          else
          cVar1S17S55P016P037N017N067(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='0' )then
          cVar1S18S55P016P036P038P037(0) <='1';
          else
          cVar1S18S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='0' )then
          cVar1S19S55P016P036P038P037(0) <='1';
          else
          cVar1S19S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='0' )then
          cVar1S20S55P016P036P038P037(0) <='1';
          else
          cVar1S20S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='1' )then
          cVar1S21S55P016P036P038P037(0) <='1';
          else
          cVar1S21S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='1' )then
          cVar1S22S55P016P036P038P037(0) <='1';
          else
          cVar1S22S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 7)='0' AND B( 0)='1' )then
          cVar1S23S55P016P036P038P037(0) <='1';
          else
          cVar1S23S55P016P036P038P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='1' AND B(15)='1' )then
          cVar1S24S55P016N036P046P024nsss(0) <='1';
          else
          cVar1S24S55P016N036P046P024nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='1' AND B(15)='0' )then
          cVar1S25S55P016N036P046N024(0) <='1';
          else
          cVar1S25S55P016N036P046N024(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='1' AND B(15)='0' )then
          cVar1S26S55P016N036P046N024(0) <='1';
          else
          cVar1S26S55P016N036P046N024(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='0' AND B( 6)='0' )then
          cVar1S27S55P016N036N046P025(0) <='1';
          else
          cVar1S27S55P016N036N046P025(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='0' AND B( 6)='0' )then
          cVar1S28S55P016N036N046P025(0) <='1';
          else
          cVar1S28S55P016N036N046P025(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='0' AND B( 6)='0' )then
          cVar1S29S55P016N036N046P025(0) <='1';
          else
          cVar1S29S55P016N036N046P025(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='0' AND B( 6)='1' )then
          cVar1S30S55P016N036N046P025(0) <='1';
          else
          cVar1S30S55P016N036N046P025(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 5)='0' AND B( 6)='1' )then
          cVar1S31S55P016N036N046P025(0) <='1';
          else
          cVar1S31S55P016N036N046P025(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='0' AND A(19)='0' )then
          cVar1S0S56P016P036P054P000(0) <='1';
          else
          cVar1S0S56P016P036P054P000(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='0' AND A(19)='0' )then
          cVar1S1S56P016P036P054P000(0) <='1';
          else
          cVar1S1S56P016P036P054P000(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='0' AND A(19)='0' )then
          cVar1S2S56P016P036P054P000(0) <='1';
          else
          cVar1S2S56P016P036P054P000(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='0' AND A(19)='1' )then
          cVar1S3S56P016P036P054P000(0) <='1';
          else
          cVar1S3S56P016P036P054P000(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='0' AND A(19)='1' )then
          cVar1S4S56P016P036P054P000(0) <='1';
          else
          cVar1S4S56P016P036P054P000(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='1' AND E( 4)='0' )then
          cVar1S5S56P016P036P054P052(0) <='1';
          else
          cVar1S5S56P016P036P054P052(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='1' AND E( 4)='0' )then
          cVar1S6S56P016P036P054P052(0) <='1';
          else
          cVar1S6S56P016P036P054P052(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='1' AND E( 4)='0' )then
          cVar1S7S56P016P036P054P052(0) <='1';
          else
          cVar1S7S56P016P036P054P052(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='1' AND E( 4)='1' )then
          cVar1S8S56P016P036P054P052(0) <='1';
          else
          cVar1S8S56P016P036P054P052(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND D( 3)='1' AND E( 4)='1' )then
          cVar1S9S56P016P036P054P052(0) <='1';
          else
          cVar1S9S56P016P036P054P052(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D(14)='1' AND A( 2)='0' )then
          cVar1S10S56P016P036P043P015nsss(0) <='1';
          else
          cVar1S10S56P016P036P043P015nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D(14)='0' AND A( 7)='0' )then
          cVar1S11S56P016P036N043P005(0) <='1';
          else
          cVar1S11S56P016P036N043P005(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D(14)='0' AND A( 7)='1' )then
          cVar1S12S56P016P036N043P005(0) <='1';
          else
          cVar1S12S56P016P036N043P005(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D(14)='0' AND A( 7)='1' )then
          cVar1S13S56P016P036N043P005(0) <='1';
          else
          cVar1S13S56P016P036N043P005(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='0' AND E(11)='1' )then
          cVar1S14S56N016P053P051P057(0) <='1';
          else
          cVar1S14S56N016P053P051P057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='0' AND E(11)='1' )then
          cVar1S15S56N016P053P051P057(0) <='1';
          else
          cVar1S15S56N016P053P051P057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='0' AND E(11)='0' )then
          cVar1S16S56N016P053P051N057(0) <='1';
          else
          cVar1S16S56N016P053P051N057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='0' AND E(11)='0' )then
          cVar1S17S56N016P053P051N057(0) <='1';
          else
          cVar1S17S56N016P053P051N057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='1' AND E(11)='0' )then
          cVar1S18S56N016P053P051P057(0) <='1';
          else
          cVar1S18S56N016P053P051P057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND D(12)='1' AND E(11)='0' )then
          cVar1S19S56N016P053P051P057(0) <='1';
          else
          cVar1S19S56N016P053P051P057(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='1' AND D( 0)='0' )then
          cVar1S20S56N016P053P028P066(0) <='1';
          else
          cVar1S20S56N016P053P028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='1' AND D( 0)='0' )then
          cVar1S21S56N016P053P028P066(0) <='1';
          else
          cVar1S21S56N016P053P028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='1' AND D( 0)='0' )then
          cVar1S22S56N016P053P028P066(0) <='1';
          else
          cVar1S22S56N016P053P028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='1' AND D( 0)='1' )then
          cVar1S23S56N016P053P028P066(0) <='1';
          else
          cVar1S23S56N016P053P028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='1' AND D( 0)='1' )then
          cVar1S24S56N016P053P028P066(0) <='1';
          else
          cVar1S24S56N016P053P028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='0' AND D( 0)='1' )then
          cVar1S25S56N016P053N028P066(0) <='1';
          else
          cVar1S25S56N016P053N028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='0' AND D( 0)='1' )then
          cVar1S26S56N016P053N028P066(0) <='1';
          else
          cVar1S26S56N016P053N028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='0' AND D( 0)='1' )then
          cVar1S27S56N016P053N028P066(0) <='1';
          else
          cVar1S27S56N016P053N028P066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='0' AND D( 0)='0' )then
          cVar1S28S56N016P053N028N066(0) <='1';
          else
          cVar1S28S56N016P053N028N066(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(13)='0' AND D( 0)='0' )then
          cVar1S29S56N016P053N028N066(0) <='1';
          else
          cVar1S29S56N016P053N028N066(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='0' )then
          cVar1S0S57P056P051P016P053(0) <='1';
          else
          cVar1S0S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='0' )then
          cVar1S1S57P056P051P016P053(0) <='1';
          else
          cVar1S1S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='0' )then
          cVar1S2S57P056P051P016P053(0) <='1';
          else
          cVar1S2S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='0' )then
          cVar1S3S57P056P051P016P053(0) <='1';
          else
          cVar1S3S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='1' )then
          cVar1S4S57P056P051P016P053(0) <='1';
          else
          cVar1S4S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='0' AND E(12)='1' )then
          cVar1S5S57P056P051P016P053(0) <='1';
          else
          cVar1S5S57P056P051P016P053(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='1' )then
          cVar1S6S57P056P051P016P036(0) <='1';
          else
          cVar1S6S57P056P051P016P036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='1' )then
          cVar1S7S57P056P051P016P036(0) <='1';
          else
          cVar1S7S57P056P051P016P036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='1' )then
          cVar1S8S57P056P051P016P036(0) <='1';
          else
          cVar1S8S57P056P051P016P036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='0' )then
          cVar1S9S57P056P051P016N036(0) <='1';
          else
          cVar1S9S57P056P051P016N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='0' )then
          cVar1S10S57P056P051P016N036(0) <='1';
          else
          cVar1S10S57P056P051P016N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='0' )then
          cVar1S11S57P056P051P016N036(0) <='1';
          else
          cVar1S11S57P056P051P016N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='0' AND A(11)='1' AND B( 9)='0' )then
          cVar1S12S57P056P051P016N036(0) <='1';
          else
          cVar1S12S57P056P051P016N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='1' AND B( 9)='1' )then
          cVar1S13S57P056P051P008P036(0) <='1';
          else
          cVar1S13S57P056P051P008P036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='1' AND B( 9)='1' )then
          cVar1S14S57P056P051P008P036(0) <='1';
          else
          cVar1S14S57P056P051P008P036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='1' AND B( 9)='0' )then
          cVar1S15S57P056P051P008N036(0) <='1';
          else
          cVar1S15S57P056P051P008N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='1' AND B( 9)='0' )then
          cVar1S16S57P056P051P008N036(0) <='1';
          else
          cVar1S16S57P056P051P008N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='1' AND B( 9)='0' )then
          cVar1S17S57P056P051P008N036(0) <='1';
          else
          cVar1S17S57P056P051P008N036(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='0' AND E( 1)='0' )then
          cVar1S18S57P056P051N008P064(0) <='1';
          else
          cVar1S18S57P056P051N008P064(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='0' AND E( 1)='0' )then
          cVar1S19S57P056P051N008P064(0) <='1';
          else
          cVar1S19S57P056P051N008P064(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='0' AND E( 1)='1' )then
          cVar1S20S57P056P051N008P064(0) <='1';
          else
          cVar1S20S57P056P051N008P064(0) <='0';
          end if;
        if(E( 3)='0' AND D(12)='1' AND A(15)='0' AND E( 1)='1' )then
          cVar1S21S57P056P051N008P064(0) <='1';
          else
          cVar1S21S57P056P051N008P064(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='0' AND B( 5)='0' AND D( 4)='0' )then
          cVar1S22S57P056P052P027P050(0) <='1';
          else
          cVar1S22S57P056P052P027P050(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='0' AND B( 5)='0' AND D( 4)='0' )then
          cVar1S23S57P056P052P027P050(0) <='1';
          else
          cVar1S23S57P056P052P027P050(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='0' AND B( 5)='0' AND D( 4)='0' )then
          cVar1S24S57P056P052P027P050(0) <='1';
          else
          cVar1S24S57P056P052P027P050(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='0' AND B( 5)='0' AND D( 4)='1' )then
          cVar1S25S57P056P052P027P050(0) <='1';
          else
          cVar1S25S57P056P052P027P050(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='1' AND A( 5)='1' )then
          cVar1S26S57P056P052P009nsss(0) <='1';
          else
          cVar1S26S57P056P052P009nsss(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='1' AND A( 5)='0' AND A(15)='1' )then
          cVar1S27S57P056P052N009P008nsss(0) <='1';
          else
          cVar1S27S57P056P052N009P008nsss(0) <='0';
          end if;
        if(E( 3)='1' AND E( 4)='1' AND A( 5)='0' AND A(15)='0' )then
          cVar1S28S57P056P052N009N008(0) <='1';
          else
          cVar1S28S57P056P052N009N008(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='1' AND D( 1)='0' )then
          cVar1S0S58P017P065P041P062(0) <='1';
          else
          cVar1S0S58P017P065P041P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='1' AND D( 1)='0' )then
          cVar1S1S58P017P065P041P062(0) <='1';
          else
          cVar1S1S58P017P065P041P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='1' AND D( 1)='0' )then
          cVar1S2S58P017P065P041P062(0) <='1';
          else
          cVar1S2S58P017P065P041P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='1' AND D( 1)='1' )then
          cVar1S3S58P017P065P041P062(0) <='1';
          else
          cVar1S3S58P017P065P041P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='0' AND D( 7)='1' )then
          cVar1S4S58P017P065N041P038(0) <='1';
          else
          cVar1S4S58P017P065N041P038(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='0' AND D( 7)='1' )then
          cVar1S5S58P017P065N041P038(0) <='1';
          else
          cVar1S5S58P017P065N041P038(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='0' AND D( 7)='0' )then
          cVar1S6S58P017P065N041N038(0) <='1';
          else
          cVar1S6S58P017P065N041N038(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='0' AND D( 7)='0' )then
          cVar1S7S58P017P065N041N038(0) <='1';
          else
          cVar1S7S58P017P065N041N038(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='0' AND E(15)='0' AND D( 7)='0' )then
          cVar1S8S58P017P065N041N038(0) <='1';
          else
          cVar1S8S58P017P065N041N038(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='0' )then
          cVar1S9S58P017P065P063P056(0) <='1';
          else
          cVar1S9S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='0' )then
          cVar1S10S58P017P065P063P056(0) <='1';
          else
          cVar1S10S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='0' )then
          cVar1S11S58P017P065P063P056(0) <='1';
          else
          cVar1S11S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='0' )then
          cVar1S12S58P017P065P063P056(0) <='1';
          else
          cVar1S12S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='1' )then
          cVar1S13S58P017P065P063P056(0) <='1';
          else
          cVar1S13S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='1' )then
          cVar1S14S58P017P065P063P056(0) <='1';
          else
          cVar1S14S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='1' AND E( 3)='1' )then
          cVar1S15S58P017P065P063P056(0) <='1';
          else
          cVar1S15S58P017P065P063P056(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='0' AND A(19)='1' )then
          cVar1S16S58P017P065N063P000(0) <='1';
          else
          cVar1S16S58P017P065N063P000(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='0' AND A(19)='0' )then
          cVar1S17S58P017P065N063N000(0) <='1';
          else
          cVar1S17S58P017P065N063N000(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='0' AND A(19)='0' )then
          cVar1S18S58P017P065N063N000(0) <='1';
          else
          cVar1S18S58P017P065N063N000(0) <='0';
          end if;
        if(A( 1)='0' AND E( 9)='1' AND D( 9)='0' AND A(19)='0' )then
          cVar1S19S58P017P065N063N000(0) <='1';
          else
          cVar1S19S58P017P065N063N000(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='1' AND B(14)='0' )then
          cVar1S20S58P017P064P037P026(0) <='1';
          else
          cVar1S20S58P017P064P037P026(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='1' AND B(14)='0' )then
          cVar1S21S58P017P064P037P026(0) <='1';
          else
          cVar1S21S58P017P064P037P026(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='1' AND B(14)='0' )then
          cVar1S22S58P017P064P037P026(0) <='1';
          else
          cVar1S22S58P017P064P037P026(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='1' AND B(14)='0' )then
          cVar1S23S58P017P064P037P026(0) <='1';
          else
          cVar1S23S58P017P064P037P026(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='0' AND A( 8)='1' )then
          cVar1S24S58P017P064N037P003(0) <='1';
          else
          cVar1S24S58P017P064N037P003(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='0' AND A( 8)='1' )then
          cVar1S25S58P017P064N037P003(0) <='1';
          else
          cVar1S25S58P017P064N037P003(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='0' AND A( 8)='1' )then
          cVar1S26S58P017P064N037P003(0) <='1';
          else
          cVar1S26S58P017P064N037P003(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='1' AND B( 0)='0' AND A( 8)='0' )then
          cVar1S27S58P017P064N037N003(0) <='1';
          else
          cVar1S27S58P017P064N037N003(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='1' AND E( 0)='0' )then
          cVar1S28S58P017N064P063P068(0) <='1';
          else
          cVar1S28S58P017N064P063P068(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='1' AND E( 0)='0' )then
          cVar1S29S58P017N064P063P068(0) <='1';
          else
          cVar1S29S58P017N064P063P068(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='1' AND E( 0)='0' )then
          cVar1S30S58P017N064P063P068(0) <='1';
          else
          cVar1S30S58P017N064P063P068(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='1' AND E( 0)='1' )then
          cVar1S31S58P017N064P063P068(0) <='1';
          else
          cVar1S31S58P017N064P063P068(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='1' AND E( 0)='1' )then
          cVar1S32S58P017N064P063P068(0) <='1';
          else
          cVar1S32S58P017N064P063P068(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='0' AND B( 9)='1' )then
          cVar1S33S58P017N064N063P036(0) <='1';
          else
          cVar1S33S58P017N064N063P036(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='0' AND B( 9)='1' )then
          cVar1S34S58P017N064N063P036(0) <='1';
          else
          cVar1S34S58P017N064N063P036(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='0' AND B( 9)='0' )then
          cVar1S35S58P017N064N063N036(0) <='1';
          else
          cVar1S35S58P017N064N063N036(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='0' AND B( 9)='0' )then
          cVar1S36S58P017N064N063N036(0) <='1';
          else
          cVar1S36S58P017N064N063N036(0) <='0';
          end if;
        if(A( 1)='1' AND E( 1)='0' AND D( 9)='0' AND B( 9)='0' )then
          cVar1S37S58P017N064N063N036(0) <='1';
          else
          cVar1S37S58P017N064N063N036(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='1' AND A( 2)='0' )then
          cVar1S0S59P063P001P035P015(0) <='1';
          else
          cVar1S0S59P063P001P035P015(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='1' AND A( 2)='0' )then
          cVar1S1S59P063P001P035P015(0) <='1';
          else
          cVar1S1S59P063P001P035P015(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='1' AND A( 2)='0' )then
          cVar1S2S59P063P001P035P015(0) <='1';
          else
          cVar1S2S59P063P001P035P015(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='1' AND A( 2)='1' )then
          cVar1S3S59P063P001P035P015(0) <='1';
          else
          cVar1S3S59P063P001P035P015(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='1' AND A( 2)='1' )then
          cVar1S4S59P063P001P035P015(0) <='1';
          else
          cVar1S4S59P063P001P035P015(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='0' AND E(11)='0' )then
          cVar1S5S59P063P001N035P057(0) <='1';
          else
          cVar1S5S59P063P001N035P057(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='0' AND E(11)='0' )then
          cVar1S6S59P063P001N035P057(0) <='1';
          else
          cVar1S6S59P063P001N035P057(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='0' AND E(11)='0' )then
          cVar1S7S59P063P001N035P057(0) <='1';
          else
          cVar1S7S59P063P001N035P057(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='0' AND E(11)='0' )then
          cVar1S8S59P063P001N035P057(0) <='1';
          else
          cVar1S8S59P063P001N035P057(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='0' AND B( 1)='0' AND E(11)='1' )then
          cVar1S9S59P063P001N035P057(0) <='1';
          else
          cVar1S9S59P063P001N035P057(0) <='0';
          end if;
        if(D( 9)='1' AND A( 9)='1' AND B(10)='1' AND E( 0)='0' )then
          cVar1S10S59P063P001P034P068(0) <='1';
          else
          cVar1S10S59P063P001P034P068(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='0' AND E( 1)='0' )then
          cVar1S11S59N063P060P054P064(0) <='1';
          else
          cVar1S11S59N063P060P054P064(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='0' AND E( 1)='0' )then
          cVar1S12S59N063P060P054P064(0) <='1';
          else
          cVar1S12S59N063P060P054P064(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='0' AND E( 1)='0' )then
          cVar1S13S59N063P060P054P064(0) <='1';
          else
          cVar1S13S59N063P060P054P064(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='0' AND E( 1)='0' )then
          cVar1S14S59N063P060P054P064(0) <='1';
          else
          cVar1S14S59N063P060P054P064(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='0' AND E( 1)='1' )then
          cVar1S15S59N063P060P054P064(0) <='1';
          else
          cVar1S15S59N063P060P054P064(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='1' AND D( 3)='1' AND E( 3)='1' )then
          cVar1S16S59N063P060P054P056(0) <='1';
          else
          cVar1S16S59N063P060P054P056(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='1' AND E( 9)='1' )then
          cVar1S17S59N063N060P064P065(0) <='1';
          else
          cVar1S17S59N063N060P064P065(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='1' AND E( 9)='0' )then
          cVar1S18S59N063N060P064N065(0) <='1';
          else
          cVar1S18S59N063N060P064N065(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S19S59N063N060N064P062(0) <='1';
          else
          cVar1S19S59N063N060N064P062(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S20S59N063N060N064P062(0) <='1';
          else
          cVar1S20S59N063N060N064P062(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S21S59N063N060N064P062(0) <='1';
          else
          cVar1S21S59N063N060N064P062(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S22S59N063N060N064P062(0) <='1';
          else
          cVar1S22S59N063N060N064P062(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S23S59N063N060N064P062(0) <='1';
          else
          cVar1S23S59N063N060N064P062(0) <='0';
          end if;
        if(D( 9)='0' AND E( 2)='0' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S24S59N063N060N064P062(0) <='1';
          else
          cVar1S24S59N063N060N064P062(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='1' )then
          cVar1S0S60P037P063P033P017(0) <='1';
          else
          cVar1S0S60P037P063P033P017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='1' )then
          cVar1S1S60P037P063P033P017(0) <='1';
          else
          cVar1S1S60P037P063P033P017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='1' )then
          cVar1S2S60P037P063P033P017(0) <='1';
          else
          cVar1S2S60P037P063P033P017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='0' )then
          cVar1S3S60P037P063P033N017(0) <='1';
          else
          cVar1S3S60P037P063P033N017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='0' )then
          cVar1S4S60P037P063P033N017(0) <='1';
          else
          cVar1S4S60P037P063P033N017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='0' AND A( 1)='0' )then
          cVar1S5S60P037P063P033N017(0) <='1';
          else
          cVar1S5S60P037P063P033N017(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='1' AND D(10)='1' )then
          cVar1S6S60P037P063P033P059(0) <='1';
          else
          cVar1S6S60P037P063P033P059(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='1' AND D(10)='1' )then
          cVar1S7S60P037P063P033P059(0) <='1';
          else
          cVar1S7S60P037P063P033P059(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='1' AND D(10)='0' )then
          cVar1S8S60P037P063P033N059(0) <='1';
          else
          cVar1S8S60P037P063P033N059(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='1' AND D(10)='0' )then
          cVar1S9S60P037P063P033N059(0) <='1';
          else
          cVar1S9S60P037P063P033N059(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='0' AND B( 2)='1' AND D(10)='0' )then
          cVar1S10S60P037P063P033N059(0) <='1';
          else
          cVar1S10S60P037P063P033N059(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='1' )then
          cVar1S11S60P037P063P068P013(0) <='1';
          else
          cVar1S11S60P037P063P068P013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='1' )then
          cVar1S12S60P037P063P068P013(0) <='1';
          else
          cVar1S12S60P037P063P068P013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='1' )then
          cVar1S13S60P037P063P068P013(0) <='1';
          else
          cVar1S13S60P037P063P068P013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='0' )then
          cVar1S14S60P037P063P068N013(0) <='1';
          else
          cVar1S14S60P037P063P068N013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='0' )then
          cVar1S15S60P037P063P068N013(0) <='1';
          else
          cVar1S15S60P037P063P068N013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='0' AND A( 3)='0' )then
          cVar1S16S60P037P063P068N013(0) <='1';
          else
          cVar1S16S60P037P063P068N013(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='1' AND E( 4)='1' )then
          cVar1S17S60P037P063P068P052nsss(0) <='1';
          else
          cVar1S17S60P037P063P068P052nsss(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='1' AND E( 4)='0' )then
          cVar1S18S60P037P063P068N052(0) <='1';
          else
          cVar1S18S60P037P063P068N052(0) <='0';
          end if;
        if(B( 0)='1' AND D( 9)='1' AND E( 0)='1' AND E( 4)='0' )then
          cVar1S19S60P037P063P068N052(0) <='1';
          else
          cVar1S19S60P037P063P068N052(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='0' AND B(16)='1' )then
          cVar1S20S60N037P035P065P022(0) <='1';
          else
          cVar1S20S60N037P035P065P022(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='0' AND B(16)='1' )then
          cVar1S21S60N037P035P065P022(0) <='1';
          else
          cVar1S21S60N037P035P065P022(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='0' AND B(16)='0' )then
          cVar1S22S60N037P035P065N022(0) <='1';
          else
          cVar1S22S60N037P035P065N022(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='0' AND B(16)='0' )then
          cVar1S23S60N037P035P065N022(0) <='1';
          else
          cVar1S23S60N037P035P065N022(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='0' AND B(16)='0' )then
          cVar1S24S60N037P035P065N022(0) <='1';
          else
          cVar1S24S60N037P035P065N022(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='1' AND A(18)='0' )then
          cVar1S25S60N037P035P065P002(0) <='1';
          else
          cVar1S25S60N037P035P065P002(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='1' AND A(18)='0' )then
          cVar1S26S60N037P035P065P002(0) <='1';
          else
          cVar1S26S60N037P035P065P002(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='0' AND E( 9)='1' AND A(18)='1' )then
          cVar1S27S60N037P035P065P002(0) <='1';
          else
          cVar1S27S60N037P035P065P002(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='1' AND E(15)='0' )then
          cVar1S28S60N037P035P065P041(0) <='1';
          else
          cVar1S28S60N037P035P065P041(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='1' AND E(15)='0' )then
          cVar1S29S60N037P035P065P041(0) <='1';
          else
          cVar1S29S60N037P035P065P041(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='1' AND E(15)='0' )then
          cVar1S30S60N037P035P065P041(0) <='1';
          else
          cVar1S30S60N037P035P065P041(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='1' )then
          cVar1S31S60N037P035N065P054(0) <='1';
          else
          cVar1S31S60N037P035N065P054(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='1' )then
          cVar1S32S60N037P035N065P054(0) <='1';
          else
          cVar1S32S60N037P035N065P054(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='1' )then
          cVar1S33S60N037P035N065P054(0) <='1';
          else
          cVar1S33S60N037P035N065P054(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='0' )then
          cVar1S34S60N037P035N065N054(0) <='1';
          else
          cVar1S34S60N037P035N065N054(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='0' )then
          cVar1S35S60N037P035N065N054(0) <='1';
          else
          cVar1S35S60N037P035N065N054(0) <='0';
          end if;
        if(B( 0)='0' AND B( 1)='1' AND E( 9)='0' AND D( 3)='0' )then
          cVar1S36S60N037P035N065N054(0) <='1';
          else
          cVar1S36S60N037P035N065N054(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S0S61P063P035P015P017(0) <='1';
          else
          cVar1S0S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S1S61P063P035P015P017(0) <='1';
          else
          cVar1S1S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S2S61P063P035P015P017(0) <='1';
          else
          cVar1S2S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S3S61P063P035P015P017(0) <='1';
          else
          cVar1S3S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S4S61P063P035P015P017(0) <='1';
          else
          cVar1S4S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S5S61P063P035P015P017(0) <='1';
          else
          cVar1S5S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S6S61P063P035P015P017(0) <='1';
          else
          cVar1S6S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S7S61P063P035P015P017(0) <='1';
          else
          cVar1S7S61P063P035P015P017(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='1' AND B( 6)='1' )then
          cVar1S8S61P063P035P015P025(0) <='1';
          else
          cVar1S8S61P063P035P015P025(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='1' AND B( 6)='1' )then
          cVar1S9S61P063P035P015P025(0) <='1';
          else
          cVar1S9S61P063P035P015P025(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='1' AND B( 6)='0' )then
          cVar1S10S61P063P035P015N025(0) <='1';
          else
          cVar1S10S61P063P035P015N025(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='1' AND B( 6)='0' )then
          cVar1S11S61P063P035P015N025(0) <='1';
          else
          cVar1S11S61P063P035P015N025(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='0' AND A( 2)='1' AND B( 6)='0' )then
          cVar1S12S61P063P035P015N025(0) <='1';
          else
          cVar1S12S61P063P035P015N025(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='1' AND D(13)='0' )then
          cVar1S13S61P063P035P014P047(0) <='1';
          else
          cVar1S13S61P063P035P014P047(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='1' AND D(13)='0' )then
          cVar1S14S61P063P035P014P047(0) <='1';
          else
          cVar1S14S61P063P035P014P047(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='1' AND D(13)='0' )then
          cVar1S15S61P063P035P014P047(0) <='1';
          else
          cVar1S15S61P063P035P014P047(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='1' )then
          cVar1S16S61P063P035N014P061(0) <='1';
          else
          cVar1S16S61P063P035N014P061(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='1' )then
          cVar1S17S61P063P035N014P061(0) <='1';
          else
          cVar1S17S61P063P035N014P061(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='1' )then
          cVar1S18S61P063P035N014P061(0) <='1';
          else
          cVar1S18S61P063P035N014P061(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='0' )then
          cVar1S19S61P063P035N014N061(0) <='1';
          else
          cVar1S19S61P063P035N014N061(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='0' )then
          cVar1S20S61P063P035N014N061(0) <='1';
          else
          cVar1S20S61P063P035N014N061(0) <='0';
          end if;
        if(D( 9)='0' AND B( 1)='1' AND A(12)='0' AND E(10)='0' )then
          cVar1S21S61P063P035N014N061(0) <='1';
          else
          cVar1S21S61P063P035N014N061(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='1' AND E( 2)='1' )then
          cVar1S22S61P063P062P068P060nsss(0) <='1';
          else
          cVar1S22S61P063P062P068P060nsss(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='1' AND E( 2)='0' )then
          cVar1S23S61P063P062P068N060(0) <='1';
          else
          cVar1S23S61P063P062P068N060(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='1' AND E( 2)='0' )then
          cVar1S24S61P063P062P068N060(0) <='1';
          else
          cVar1S24S61P063P062P068N060(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='1' AND E( 2)='0' )then
          cVar1S25S61P063P062P068N060(0) <='1';
          else
          cVar1S25S61P063P062P068N060(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='0' AND B(16)='0' )then
          cVar1S26S61P063P062N068P022(0) <='1';
          else
          cVar1S26S61P063P062N068P022(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='0' AND B(16)='0' )then
          cVar1S27S61P063P062N068P022(0) <='1';
          else
          cVar1S27S61P063P062N068P022(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='0' AND B(16)='0' )then
          cVar1S28S61P063P062N068P022(0) <='1';
          else
          cVar1S28S61P063P062N068P022(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='1' AND E( 0)='0' AND B(16)='0' )then
          cVar1S29S61P063P062N068P022(0) <='1';
          else
          cVar1S29S61P063P062N068P022(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND A(18)='0' AND B( 1)='1' )then
          cVar1S30S61P063N062P002P035(0) <='1';
          else
          cVar1S30S61P063N062P002P035(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND A(18)='0' AND B( 1)='0' )then
          cVar1S31S61P063N062P002N035(0) <='1';
          else
          cVar1S31S61P063N062P002N035(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND A(18)='0' AND B( 1)='0' )then
          cVar1S32S61P063N062P002N035(0) <='1';
          else
          cVar1S32S61P063N062P002N035(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND A(18)='1' AND B( 0)='1' )then
          cVar1S33S61P063N062P002P037(0) <='1';
          else
          cVar1S33S61P063N062P002P037(0) <='0';
          end if;
        if(D( 9)='1' AND D( 1)='0' AND A(18)='1' AND B( 0)='0' )then
          cVar1S34S61P063N062P002N037(0) <='1';
          else
          cVar1S34S61P063N062P002N037(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='0' AND B(16)='0' )then
          cVar1S0S62P062P017P048P022(0) <='1';
          else
          cVar1S0S62P062P017P048P022(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='0' AND B(16)='0' )then
          cVar1S1S62P062P017P048P022(0) <='1';
          else
          cVar1S1S62P062P017P048P022(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='0' AND B(16)='0' )then
          cVar1S2S62P062P017P048P022(0) <='1';
          else
          cVar1S2S62P062P017P048P022(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='0' AND B(16)='0' )then
          cVar1S3S62P062P017P048P022(0) <='1';
          else
          cVar1S3S62P062P017P048P022(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='1' AND D( 5)='1' )then
          cVar1S4S62P062P017P048P046nsss(0) <='1';
          else
          cVar1S4S62P062P017P048P046nsss(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='1' AND E( 5)='1' AND D( 5)='0' )then
          cVar1S5S62P062P017P048N046(0) <='1';
          else
          cVar1S5S62P062P017P048N046(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='0' AND A( 7)='0' )then
          cVar1S6S62P062N017P047P005(0) <='1';
          else
          cVar1S6S62P062N017P047P005(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='0' AND A( 7)='0' )then
          cVar1S7S62P062N017P047P005(0) <='1';
          else
          cVar1S7S62P062N017P047P005(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='0' AND A( 7)='0' )then
          cVar1S8S62P062N017P047P005(0) <='1';
          else
          cVar1S8S62P062N017P047P005(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='0' AND A( 7)='1' )then
          cVar1S9S62P062N017P047P005(0) <='1';
          else
          cVar1S9S62P062N017P047P005(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='0' AND A( 7)='1' )then
          cVar1S10S62P062N017P047P005(0) <='1';
          else
          cVar1S10S62P062N017P047P005(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='1' AND B(14)='1' )then
          cVar1S11S62P062N017P047P026nsss(0) <='1';
          else
          cVar1S11S62P062N017P047P026nsss(0) <='0';
          end if;
        if(D( 1)='1' AND A( 1)='0' AND D(13)='1' AND B(14)='0' )then
          cVar1S12S62P062N017P047N026(0) <='1';
          else
          cVar1S12S62P062N017P047N026(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='0' )then
          cVar1S13S62N062P066P067P059(0) <='1';
          else
          cVar1S13S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='0' )then
          cVar1S14S62N062P066P067P059(0) <='1';
          else
          cVar1S14S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='0' )then
          cVar1S15S62N062P066P067P059(0) <='1';
          else
          cVar1S15S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='1' )then
          cVar1S16S62N062P066P067P059(0) <='1';
          else
          cVar1S16S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='1' )then
          cVar1S17S62N062P066P067P059(0) <='1';
          else
          cVar1S17S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='1' )then
          cVar1S18S62N062P066P067P059(0) <='1';
          else
          cVar1S18S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='0' AND D(10)='1' )then
          cVar1S19S62N062P066P067P059(0) <='1';
          else
          cVar1S19S62N062P066P067P059(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='1' )then
          cVar1S20S62N062P066P067P016(0) <='1';
          else
          cVar1S20S62N062P066P067P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='1' )then
          cVar1S21S62N062P066P067P016(0) <='1';
          else
          cVar1S21S62N062P066P067P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='1' )then
          cVar1S22S62N062P066P067P016(0) <='1';
          else
          cVar1S22S62N062P066P067P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='0' )then
          cVar1S23S62N062P066P067N016(0) <='1';
          else
          cVar1S23S62N062P066P067N016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='0' )then
          cVar1S24S62N062P066P067N016(0) <='1';
          else
          cVar1S24S62N062P066P067N016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='1' AND D( 8)='1' AND A(11)='0' )then
          cVar1S25S62N062P066P067N016(0) <='1';
          else
          cVar1S25S62N062P066P067N016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='1' )then
          cVar1S26S62N062N066P034P010(0) <='1';
          else
          cVar1S26S62N062N066P034P010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='1' )then
          cVar1S27S62N062N066P034P010(0) <='1';
          else
          cVar1S27S62N062N066P034P010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='1' )then
          cVar1S28S62N062N066P034P010(0) <='1';
          else
          cVar1S28S62N062N066P034P010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='0' )then
          cVar1S29S62N062N066P034N010(0) <='1';
          else
          cVar1S29S62N062N066P034N010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='0' )then
          cVar1S30S62N062N066P034N010(0) <='1';
          else
          cVar1S30S62N062N066P034N010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='0' AND A(14)='0' )then
          cVar1S31S62N062N066P034N010(0) <='1';
          else
          cVar1S31S62N062N066P034N010(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='1' )then
          cVar1S32S62N062N066P034P016(0) <='1';
          else
          cVar1S32S62N062N066P034P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='1' )then
          cVar1S33S62N062N066P034P016(0) <='1';
          else
          cVar1S33S62N062N066P034P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='1' )then
          cVar1S34S62N062N066P034P016(0) <='1';
          else
          cVar1S34S62N062N066P034P016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='0' )then
          cVar1S35S62N062N066P034N016(0) <='1';
          else
          cVar1S35S62N062N066P034N016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='0' )then
          cVar1S36S62N062N066P034N016(0) <='1';
          else
          cVar1S36S62N062N066P034N016(0) <='0';
          end if;
        if(D( 1)='0' AND D( 0)='0' AND B(10)='1' AND A(11)='0' )then
          cVar1S37S62N062N066P034N016(0) <='1';
          else
          cVar1S37S62N062N066P034N016(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='0' AND D( 1)='0' )then
          cVar1S0S63P067P018P050P062(0) <='1';
          else
          cVar1S0S63P067P018P050P062(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='0' AND D( 1)='0' )then
          cVar1S1S63P067P018P050P062(0) <='1';
          else
          cVar1S1S63P067P018P050P062(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='0' AND D( 1)='0' )then
          cVar1S2S63P067P018P050P062(0) <='1';
          else
          cVar1S2S63P067P018P050P062(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='0' AND D( 1)='1' )then
          cVar1S3S63P067P018P050P062(0) <='1';
          else
          cVar1S3S63P067P018P050P062(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='0' AND D( 1)='1' )then
          cVar1S4S63P067P018P050P062(0) <='1';
          else
          cVar1S4S63P067P018P050P062(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='1' AND A(14)='1' )then
          cVar1S5S63P067P018P050P010(0) <='1';
          else
          cVar1S5S63P067P018P050P010(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='1' AND A(14)='0' )then
          cVar1S6S63P067P018P050N010(0) <='1';
          else
          cVar1S6S63P067P018P050N010(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='1' AND D( 4)='1' AND A(14)='0' )then
          cVar1S7S63P067P018P050N010(0) <='1';
          else
          cVar1S7S63P067P018P050N010(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='1' AND E(13)='0' )then
          cVar1S8S63P067N018P068P049(0) <='1';
          else
          cVar1S8S63P067N018P068P049(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='1' AND E(13)='0' )then
          cVar1S9S63P067N018P068P049(0) <='1';
          else
          cVar1S9S63P067N018P068P049(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='1' )then
          cVar1S10S63P067N018N068P015(0) <='1';
          else
          cVar1S10S63P067N018N068P015(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='1' )then
          cVar1S11S63P067N018N068P015(0) <='1';
          else
          cVar1S11S63P067N018N068P015(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='1' )then
          cVar1S12S63P067N018N068P015(0) <='1';
          else
          cVar1S12S63P067N018N068P015(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='0' )then
          cVar1S13S63P067N018N068N015(0) <='1';
          else
          cVar1S13S63P067N018N068N015(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='0' )then
          cVar1S14S63P067N018N068N015(0) <='1';
          else
          cVar1S14S63P067N018N068N015(0) <='0';
          end if;
        if(D( 8)='1' AND A(10)='0' AND E( 0)='0' AND A( 2)='0' )then
          cVar1S15S63P067N018N068N015(0) <='1';
          else
          cVar1S15S63P067N018N068N015(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='1' )then
          cVar1S16S63N067P044P028nsss(0) <='1';
          else
          cVar1S16S63N067P044P028nsss(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='0' AND B( 7)='1' )then
          cVar1S17S63N067P044N028P023(0) <='1';
          else
          cVar1S17S63N067P044N028P023(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='0' AND B( 7)='0' )then
          cVar1S18S63N067P044N028N023(0) <='1';
          else
          cVar1S18S63N067P044N028N023(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='0' AND B( 7)='0' )then
          cVar1S19S63N067P044N028N023(0) <='1';
          else
          cVar1S19S63N067P044N028N023(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='0' AND B( 7)='0' )then
          cVar1S20S63N067P044N028N023(0) <='1';
          else
          cVar1S20S63N067P044N028N023(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='1' AND B(13)='0' AND B( 7)='0' )then
          cVar1S21S63N067P044N028N023(0) <='1';
          else
          cVar1S21S63N067P044N028N023(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='1' AND E(13)='0' )then
          cVar1S22S63N067N044P059P049(0) <='1';
          else
          cVar1S22S63N067N044P059P049(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='1' AND E(13)='0' )then
          cVar1S23S63N067N044P059P049(0) <='1';
          else
          cVar1S23S63N067N044P059P049(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='1' AND E(13)='0' )then
          cVar1S24S63N067N044P059P049(0) <='1';
          else
          cVar1S24S63N067N044P059P049(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='1' AND E(13)='1' )then
          cVar1S25S63N067N044P059P049(0) <='1';
          else
          cVar1S25S63N067N044P059P049(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='1' )then
          cVar1S26S63N067N044N059P031(0) <='1';
          else
          cVar1S26S63N067N044N059P031(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='1' )then
          cVar1S27S63N067N044N059P031(0) <='1';
          else
          cVar1S27S63N067N044N059P031(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='1' )then
          cVar1S28S63N067N044N059P031(0) <='1';
          else
          cVar1S28S63N067N044N059P031(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='0' )then
          cVar1S29S63N067N044N059N031(0) <='1';
          else
          cVar1S29S63N067N044N059N031(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='0' )then
          cVar1S30S63N067N044N059N031(0) <='1';
          else
          cVar1S30S63N067N044N059N031(0) <='0';
          end if;
        if(D( 8)='0' AND E( 6)='0' AND D(10)='0' AND B( 3)='0' )then
          cVar1S31S63N067N044N059N031(0) <='1';
          else
          cVar1S31S63N067N044N059N031(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='1' AND B(11)='1' )then
          cVar1S0S64P059P061P058P032(0) <='1';
          else
          cVar1S0S64P059P061P058P032(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='1' AND B(11)='1' )then
          cVar1S1S64P059P061P058P032(0) <='1';
          else
          cVar1S1S64P059P061P058P032(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='1' AND B(11)='0' )then
          cVar1S2S64P059P061P058N032(0) <='1';
          else
          cVar1S2S64P059P061P058N032(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='1' AND B(11)='0' )then
          cVar1S3S64P059P061P058N032(0) <='1';
          else
          cVar1S3S64P059P061P058N032(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='1' AND B(11)='0' )then
          cVar1S4S64P059P061P058N032(0) <='1';
          else
          cVar1S4S64P059P061P058N032(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S5S64P059P061N058P033(0) <='1';
          else
          cVar1S5S64P059P061N058P033(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S6S64P059P061N058P033(0) <='1';
          else
          cVar1S6S64P059P061N058P033(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='0' AND B( 2)='1' )then
          cVar1S7S64P059P061N058P033(0) <='1';
          else
          cVar1S7S64P059P061N058P033(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='0' AND D( 2)='0' AND B( 2)='1' )then
          cVar1S8S64P059P061N058P033(0) <='1';
          else
          cVar1S8S64P059P061N058P033(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='1' AND D( 8)='0' AND E( 8)='1' )then
          cVar1S9S64P059P061P067P069nsss(0) <='1';
          else
          cVar1S9S64P059P061P067P069nsss(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='1' AND D( 8)='0' AND E( 8)='0' )then
          cVar1S10S64P059P061P067N069(0) <='1';
          else
          cVar1S10S64P059P061P067N069(0) <='0';
          end if;
        if(D(10)='0' AND E(10)='1' AND D( 8)='1' AND B( 0)='1' )then
          cVar1S11S64P059P061P067P037(0) <='1';
          else
          cVar1S11S64P059P061P067P037(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='1' AND A(17)='0' )then
          cVar1S12S64P059P049P030P004(0) <='1';
          else
          cVar1S12S64P059P049P030P004(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='1' AND A(17)='0' )then
          cVar1S13S64P059P049P030P004(0) <='1';
          else
          cVar1S13S64P059P049P030P004(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='1' AND A(17)='0' )then
          cVar1S14S64P059P049P030P004(0) <='1';
          else
          cVar1S14S64P059P049P030P004(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='0' AND A( 7)='0' )then
          cVar1S15S64P059P049N030P005(0) <='1';
          else
          cVar1S15S64P059P049N030P005(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='0' AND A( 7)='0' )then
          cVar1S16S64P059P049N030P005(0) <='1';
          else
          cVar1S16S64P059P049N030P005(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='0' AND A( 7)='0' )then
          cVar1S17S64P059P049N030P005(0) <='1';
          else
          cVar1S17S64P059P049N030P005(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='0' AND A( 7)='1' )then
          cVar1S18S64P059P049N030P005(0) <='1';
          else
          cVar1S18S64P059P049N030P005(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='0' AND B(12)='0' AND A( 7)='1' )then
          cVar1S19S64P059P049N030P005(0) <='1';
          else
          cVar1S19S64P059P049N030P005(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='1' AND D(11)='0' AND D(12)='1' )then
          cVar1S20S64P059P049P055P051nsss(0) <='1';
          else
          cVar1S20S64P059P049P055P051nsss(0) <='0';
          end if;
        if(D(10)='1' AND E(13)='1' AND D(11)='0' AND D(12)='0' )then
          cVar1S21S64P059P049P055N051(0) <='1';
          else
          cVar1S21S64P059P049P055N051(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='1' AND B(14)='1' )then
          cVar1S0S65P058P054P047P026nsss(0) <='1';
          else
          cVar1S0S65P058P054P047P026nsss(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='1' AND B(14)='0' )then
          cVar1S1S65P058P054P047N026(0) <='1';
          else
          cVar1S1S65P058P054P047N026(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='1' )then
          cVar1S2S65P058P054N047P013(0) <='1';
          else
          cVar1S2S65P058P054N047P013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='1' )then
          cVar1S3S65P058P054N047P013(0) <='1';
          else
          cVar1S3S65P058P054N047P013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='1' )then
          cVar1S4S65P058P054N047P013(0) <='1';
          else
          cVar1S4S65P058P054N047P013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='0' )then
          cVar1S5S65P058P054N047N013(0) <='1';
          else
          cVar1S5S65P058P054N047N013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='0' )then
          cVar1S6S65P058P054N047N013(0) <='1';
          else
          cVar1S6S65P058P054N047N013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='0' AND D(13)='0' AND A( 3)='0' )then
          cVar1S7S65P058P054N047N013(0) <='1';
          else
          cVar1S7S65P058P054N047N013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='1' AND A( 2)='1' AND A( 3)='1' )then
          cVar1S8S65P058P054P015P013nsss(0) <='1';
          else
          cVar1S8S65P058P054P015P013nsss(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='1' AND A( 2)='1' AND A( 3)='0' )then
          cVar1S9S65P058P054P015N013(0) <='1';
          else
          cVar1S9S65P058P054P015N013(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='1' AND A( 2)='0' AND B( 2)='1' )then
          cVar1S10S65P058P054N015P033(0) <='1';
          else
          cVar1S10S65P058P054N015P033(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='1' AND A( 2)='0' AND B( 2)='1' )then
          cVar1S11S65P058P054N015P033(0) <='1';
          else
          cVar1S11S65P058P054N015P033(0) <='0';
          end if;
        if(D( 2)='1' AND D( 3)='1' AND A( 2)='0' AND B( 2)='0' )then
          cVar1S12S65P058P054N015N033(0) <='1';
          else
          cVar1S12S65P058P054N015N033(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='1' AND A( 8)='1' )then
          cVar1S13S65N058P043P022P003nsss(0) <='1';
          else
          cVar1S13S65N058P043P022P003nsss(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='1' AND A( 8)='0' )then
          cVar1S14S65N058P043P022N003(0) <='1';
          else
          cVar1S14S65N058P043P022N003(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='1' AND A( 8)='0' )then
          cVar1S15S65N058P043P022N003(0) <='1';
          else
          cVar1S15S65N058P043P022N003(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='0' AND D(13)='0' )then
          cVar1S16S65N058P043N022P047(0) <='1';
          else
          cVar1S16S65N058P043N022P047(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='0' AND D(13)='0' )then
          cVar1S17S65N058P043N022P047(0) <='1';
          else
          cVar1S17S65N058P043N022P047(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='1' AND B(16)='0' AND D(13)='0' )then
          cVar1S18S65N058P043N022P047(0) <='1';
          else
          cVar1S18S65N058P043N022P047(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='1' AND A(18)='1' )then
          cVar1S19S65N058N043P040P002(0) <='1';
          else
          cVar1S19S65N058N043P040P002(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='1' AND A(18)='1' )then
          cVar1S20S65N058N043P040P002(0) <='1';
          else
          cVar1S20S65N058N043P040P002(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='1' AND A(18)='1' )then
          cVar1S21S65N058N043P040P002(0) <='1';
          else
          cVar1S21S65N058N043P040P002(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='1' AND A(18)='0' )then
          cVar1S22S65N058N043P040N002(0) <='1';
          else
          cVar1S22S65N058N043P040N002(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='1' AND A(18)='0' )then
          cVar1S23S65N058N043P040N002(0) <='1';
          else
          cVar1S23S65N058N043P040N002(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='0' AND D( 7)='0' )then
          cVar1S24S65N058N043N040P038(0) <='1';
          else
          cVar1S24S65N058N043N040P038(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='0' AND D( 7)='0' )then
          cVar1S25S65N058N043N040P038(0) <='1';
          else
          cVar1S25S65N058N043N040P038(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='0' AND D( 7)='0' )then
          cVar1S26S65N058N043N040P038(0) <='1';
          else
          cVar1S26S65N058N043N040P038(0) <='0';
          end if;
        if(D( 2)='0' AND D(14)='0' AND E( 7)='0' AND D( 7)='1' )then
          cVar1S27S65N058N043N040P038(0) <='1';
          else
          cVar1S27S65N058N043N040P038(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 6)='1' )then
          cVar1S0S66P015P044P025nsss(0) <='1';
          else
          cVar1S0S66P015P044P025nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 6)='0' AND B( 7)='1' )then
          cVar1S1S66P015P044N025P023nsss(0) <='1';
          else
          cVar1S1S66P015P044N025P023nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 6)='0' AND B( 7)='0' )then
          cVar1S2S66P015P044N025N023(0) <='1';
          else
          cVar1S2S66P015P044N025N023(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 6)='0' AND B( 7)='0' )then
          cVar1S3S66P015P044N025N023(0) <='1';
          else
          cVar1S3S66P015P044N025N023(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='1' )then
          cVar1S4S66P015N044P003P055(0) <='1';
          else
          cVar1S4S66P015N044P003P055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S5S66P015N044P003N055(0) <='1';
          else
          cVar1S5S66P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S6S66P015N044P003N055(0) <='1';
          else
          cVar1S6S66P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S7S66P015N044P003N055(0) <='1';
          else
          cVar1S7S66P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='1' )then
          cVar1S8S66P015N044N003P027(0) <='1';
          else
          cVar1S8S66P015N044N003P027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S9S66P015N044N003N027(0) <='1';
          else
          cVar1S9S66P015N044N003N027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S10S66P015N044N003N027(0) <='1';
          else
          cVar1S10S66P015N044N003N027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S11S66P015N044N003N027(0) <='1';
          else
          cVar1S11S66P015N044N003N027(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='1' AND D( 8)='0' )then
          cVar1S12S66N015P063P037P067(0) <='1';
          else
          cVar1S12S66N015P063P037P067(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='1' AND D( 8)='0' )then
          cVar1S13S66N015P063P037P067(0) <='1';
          else
          cVar1S13S66N015P063P037P067(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='1' AND D( 8)='0' )then
          cVar1S14S66N015P063P037P067(0) <='1';
          else
          cVar1S14S66N015P063P037P067(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='1' AND D( 8)='1' )then
          cVar1S15S66N015P063P037P067(0) <='1';
          else
          cVar1S15S66N015P063P037P067(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='1' AND D( 8)='1' )then
          cVar1S16S66N015P063P037P067(0) <='1';
          else
          cVar1S16S66N015P063P037P067(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='1' )then
          cVar1S17S66N015P063N037P017(0) <='1';
          else
          cVar1S17S66N015P063N037P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='1' )then
          cVar1S18S66N015P063N037P017(0) <='1';
          else
          cVar1S18S66N015P063N037P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='1' )then
          cVar1S19S66N015P063N037P017(0) <='1';
          else
          cVar1S19S66N015P063N037P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='0' )then
          cVar1S20S66N015P063N037N017(0) <='1';
          else
          cVar1S20S66N015P063N037N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='0' )then
          cVar1S21S66N015P063N037N017(0) <='1';
          else
          cVar1S21S66N015P063N037N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='1' AND B( 0)='0' AND A( 1)='0' )then
          cVar1S22S66N015P063N037N017(0) <='1';
          else
          cVar1S22S66N015P063N037N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='1' AND D( 2)='0' )then
          cVar1S23S66N015N063P029P058(0) <='1';
          else
          cVar1S23S66N015N063P029P058(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='1' AND D( 2)='0' )then
          cVar1S24S66N015N063P029P058(0) <='1';
          else
          cVar1S24S66N015N063P029P058(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='1' AND D( 2)='0' )then
          cVar1S25S66N015N063P029P058(0) <='1';
          else
          cVar1S25S66N015N063P029P058(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='1' AND D( 2)='0' )then
          cVar1S26S66N015N063P029P058(0) <='1';
          else
          cVar1S26S66N015N063P029P058(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='1' AND D( 2)='1' )then
          cVar1S27S66N015N063P029P058(0) <='1';
          else
          cVar1S27S66N015N063P029P058(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='1' )then
          cVar1S28S66N015N063N029P028(0) <='1';
          else
          cVar1S28S66N015N063N029P028(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='1' )then
          cVar1S29S66N015N063N029P028(0) <='1';
          else
          cVar1S29S66N015N063N029P028(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S30S66N015N063N029N028(0) <='1';
          else
          cVar1S30S66N015N063N029N028(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S31S66N015N063N029N028(0) <='1';
          else
          cVar1S31S66N015N063N029N028(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S32S66N015N063N029N028(0) <='1';
          else
          cVar1S32S66N015N063N029N028(0) <='0';
          end if;
        if(A( 2)='0' AND D( 9)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S33S66N015N063N029N028(0) <='1';
          else
          cVar1S33S66N015N063N029N028(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='0' )then
          cVar1S0S67P015P014P050P061(0) <='1';
          else
          cVar1S0S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='0' )then
          cVar1S1S67P015P014P050P061(0) <='1';
          else
          cVar1S1S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='0' )then
          cVar1S2S67P015P014P050P061(0) <='1';
          else
          cVar1S2S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='0' )then
          cVar1S3S67P015P014P050P061(0) <='1';
          else
          cVar1S3S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='1' )then
          cVar1S4S67P015P014P050P061(0) <='1';
          else
          cVar1S4S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='1' )then
          cVar1S5S67P015P014P050P061(0) <='1';
          else
          cVar1S5S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='0' AND E(10)='1' )then
          cVar1S6S67P015P014P050P061(0) <='1';
          else
          cVar1S6S67P015P014P050P061(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='1' AND A( 4)='1' )then
          cVar1S7S67P015P014P050P011(0) <='1';
          else
          cVar1S7S67P015P014P050P011(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='1' AND A( 4)='1' )then
          cVar1S8S67P015P014P050P011(0) <='1';
          else
          cVar1S8S67P015P014P050P011(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='1' AND A( 4)='0' )then
          cVar1S9S67P015P014P050N011(0) <='1';
          else
          cVar1S9S67P015P014P050N011(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='1' AND A( 4)='0' )then
          cVar1S10S67P015P014P050N011(0) <='1';
          else
          cVar1S10S67P015P014P050N011(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='0' AND D( 4)='1' AND A( 4)='0' )then
          cVar1S11S67P015P014P050N011(0) <='1';
          else
          cVar1S11S67P015P014P050N011(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='0' )then
          cVar1S12S67P015P014P021P012(0) <='1';
          else
          cVar1S12S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='0' )then
          cVar1S13S67P015P014P021P012(0) <='1';
          else
          cVar1S13S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='0' )then
          cVar1S14S67P015P014P021P012(0) <='1';
          else
          cVar1S14S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='0' )then
          cVar1S15S67P015P014P021P012(0) <='1';
          else
          cVar1S15S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='1' )then
          cVar1S16S67P015P014P021P012(0) <='1';
          else
          cVar1S16S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='0' AND A(13)='1' )then
          cVar1S17S67P015P014P021P012(0) <='1';
          else
          cVar1S17S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='1' AND A(13)='0' )then
          cVar1S18S67P015P014P021P012(0) <='1';
          else
          cVar1S18S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='0' AND A(12)='1' AND B( 8)='1' AND A(13)='0' )then
          cVar1S19S67P015P014P021P012(0) <='1';
          else
          cVar1S19S67P015P014P021P012(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 3)='0' AND A(16)='1' )then
          cVar1S20S67P015P044P031P006nsss(0) <='1';
          else
          cVar1S20S67P015P044P031P006nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 3)='0' AND A(16)='0' )then
          cVar1S21S67P015P044P031N006(0) <='1';
          else
          cVar1S21S67P015P044P031N006(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='1' AND B( 3)='0' AND A(16)='0' )then
          cVar1S22S67P015P044P031N006(0) <='1';
          else
          cVar1S22S67P015P044P031N006(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='1' )then
          cVar1S23S67P015N044P003P055nsss(0) <='1';
          else
          cVar1S23S67P015N044P003P055nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S24S67P015N044P003N055(0) <='1';
          else
          cVar1S24S67P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S25S67P015N044P003N055(0) <='1';
          else
          cVar1S25S67P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='1' AND D(11)='0' )then
          cVar1S26S67P015N044P003N055(0) <='1';
          else
          cVar1S26S67P015N044P003N055(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='1' )then
          cVar1S27S67P015N044N003P027(0) <='1';
          else
          cVar1S27S67P015N044N003P027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='1' )then
          cVar1S28S67P015N044N003P027(0) <='1';
          else
          cVar1S28S67P015N044N003P027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S29S67P015N044N003N027(0) <='1';
          else
          cVar1S29S67P015N044N003N027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S30S67P015N044N003N027(0) <='1';
          else
          cVar1S30S67P015N044N003N027(0) <='0';
          end if;
        if(A( 2)='1' AND E( 6)='0' AND A( 8)='0' AND B( 5)='0' )then
          cVar1S31S67P015N044N003N027(0) <='1';
          else
          cVar1S31S67P015N044N003N027(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='1' )then
          cVar1S0S68P014P012P021P032(0) <='1';
          else
          cVar1S0S68P014P012P021P032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='1' )then
          cVar1S1S68P014P012P021P032(0) <='1';
          else
          cVar1S1S68P014P012P021P032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='1' )then
          cVar1S2S68P014P012P021P032(0) <='1';
          else
          cVar1S2S68P014P012P021P032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='0' )then
          cVar1S3S68P014P012P021N032(0) <='1';
          else
          cVar1S3S68P014P012P021N032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='0' )then
          cVar1S4S68P014P012P021N032(0) <='1';
          else
          cVar1S4S68P014P012P021N032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='0' )then
          cVar1S5S68P014P012P021N032(0) <='1';
          else
          cVar1S5S68P014P012P021N032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='0' AND B(11)='0' )then
          cVar1S6S68P014P012P021N032(0) <='1';
          else
          cVar1S6S68P014P012P021N032(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='0' AND B( 8)='1' AND B(14)='0' )then
          cVar1S7S68P014P012P021P026(0) <='1';
          else
          cVar1S7S68P014P012P021P026(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='1' AND A(14)='1' )then
          cVar1S8S68P014P012P001P010nsss(0) <='1';
          else
          cVar1S8S68P014P012P001P010nsss(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='1' AND A(14)='0' )then
          cVar1S9S68P014P012P001N010(0) <='1';
          else
          cVar1S9S68P014P012P001N010(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='1' AND A(14)='0' )then
          cVar1S10S68P014P012P001N010(0) <='1';
          else
          cVar1S10S68P014P012P001N010(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='0' AND A( 5)='0' )then
          cVar1S11S68P014P012N001P009(0) <='1';
          else
          cVar1S11S68P014P012N001P009(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='0' AND A( 5)='0' )then
          cVar1S12S68P014P012N001P009(0) <='1';
          else
          cVar1S12S68P014P012N001P009(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='0' AND A( 5)='0' )then
          cVar1S13S68P014P012N001P009(0) <='1';
          else
          cVar1S13S68P014P012N001P009(0) <='0';
          end if;
        if(A(12)='1' AND A(13)='1' AND A( 9)='0' AND A( 5)='1' )then
          cVar1S14S68P014P012N001P009(0) <='1';
          else
          cVar1S14S68P014P012N001P009(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='1' AND D( 9)='0' )then
          cVar1S15S68N014P027P009P063(0) <='1';
          else
          cVar1S15S68N014P027P009P063(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='1' AND D( 9)='0' )then
          cVar1S16S68N014P027P009P063(0) <='1';
          else
          cVar1S16S68N014P027P009P063(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='1' AND D( 9)='0' )then
          cVar1S17S68N014P027P009P063(0) <='1';
          else
          cVar1S17S68N014P027P009P063(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='1' AND D( 9)='1' )then
          cVar1S18S68N014P027P009P063(0) <='1';
          else
          cVar1S18S68N014P027P009P063(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='0' AND B(14)='0' )then
          cVar1S19S68N014P027N009P026(0) <='1';
          else
          cVar1S19S68N014P027N009P026(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='0' AND B(14)='0' )then
          cVar1S20S68N014P027N009P026(0) <='1';
          else
          cVar1S20S68N014P027N009P026(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='1' AND A( 5)='0' AND B(14)='1' )then
          cVar1S21S68N014P027N009P026(0) <='1';
          else
          cVar1S21S68N014P027N009P026(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S22S68N014N027P017P069(0) <='1';
          else
          cVar1S22S68N014N027P017P069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S23S68N014N027P017P069(0) <='1';
          else
          cVar1S23S68N014N027P017P069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S24S68N014N027P017P069(0) <='1';
          else
          cVar1S24S68N014N027P017P069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S25S68N014N027P017P069(0) <='1';
          else
          cVar1S25S68N014N027P017P069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S26S68N014N027P017N069(0) <='1';
          else
          cVar1S26S68N014N027P017N069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S27S68N014N027P017N069(0) <='1';
          else
          cVar1S27S68N014N027P017N069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S28S68N014N027P017N069(0) <='1';
          else
          cVar1S28S68N014N027P017N069(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='1' AND E(10)='1' )then
          cVar1S29S68N014N027P017P061(0) <='1';
          else
          cVar1S29S68N014N027P017P061(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='1' AND E(10)='1' )then
          cVar1S30S68N014N027P017P061(0) <='1';
          else
          cVar1S30S68N014N027P017P061(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='1' AND E(10)='0' )then
          cVar1S31S68N014N027P017N061(0) <='1';
          else
          cVar1S31S68N014N027P017N061(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='1' AND E(10)='0' )then
          cVar1S32S68N014N027P017N061(0) <='1';
          else
          cVar1S32S68N014N027P017N061(0) <='0';
          end if;
        if(A(12)='0' AND B( 5)='0' AND A( 1)='1' AND E(10)='0' )then
          cVar1S33S68N014N027P017N061(0) <='1';
          else
          cVar1S33S68N014N027P017N061(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='1' )then
          cVar1S0S69P017P062P034P064(0) <='1';
          else
          cVar1S0S69P017P062P034P064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='1' )then
          cVar1S1S69P017P062P034P064(0) <='1';
          else
          cVar1S1S69P017P062P034P064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='1' )then
          cVar1S2S69P017P062P034P064(0) <='1';
          else
          cVar1S2S69P017P062P034P064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='1' )then
          cVar1S3S69P017P062P034P064(0) <='1';
          else
          cVar1S3S69P017P062P034P064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='0' )then
          cVar1S4S69P017P062P034N064(0) <='1';
          else
          cVar1S4S69P017P062P034N064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='0' )then
          cVar1S5S69P017P062P034N064(0) <='1';
          else
          cVar1S5S69P017P062P034N064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='0' AND E( 1)='0' )then
          cVar1S6S69P017P062P034N064(0) <='1';
          else
          cVar1S6S69P017P062P034N064(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='1' )then
          cVar1S7S69P017P062P034P060(0) <='1';
          else
          cVar1S7S69P017P062P034P060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='1' )then
          cVar1S8S69P017P062P034P060(0) <='1';
          else
          cVar1S8S69P017P062P034P060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='0' )then
          cVar1S9S69P017P062P034N060(0) <='1';
          else
          cVar1S9S69P017P062P034N060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='0' )then
          cVar1S10S69P017P062P034N060(0) <='1';
          else
          cVar1S10S69P017P062P034N060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='0' )then
          cVar1S11S69P017P062P034N060(0) <='1';
          else
          cVar1S11S69P017P062P034N060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND B(10)='1' AND E( 2)='0' )then
          cVar1S12S69P017P062P034N060(0) <='1';
          else
          cVar1S12S69P017P062P034N060(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='1' )then
          cVar1S13S69P017N062P014P054(0) <='1';
          else
          cVar1S13S69P017N062P014P054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='1' )then
          cVar1S14S69P017N062P014P054(0) <='1';
          else
          cVar1S14S69P017N062P014P054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='1' )then
          cVar1S15S69P017N062P014P054(0) <='1';
          else
          cVar1S15S69P017N062P014P054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='0' )then
          cVar1S16S69P017N062P014N054(0) <='1';
          else
          cVar1S16S69P017N062P014N054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='0' )then
          cVar1S17S69P017N062P014N054(0) <='1';
          else
          cVar1S17S69P017N062P014N054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='0' AND D( 3)='0' )then
          cVar1S18S69P017N062P014N054(0) <='1';
          else
          cVar1S18S69P017N062P014N054(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='1' AND B( 1)='0' )then
          cVar1S19S69P017N062P014P035(0) <='1';
          else
          cVar1S19S69P017N062P014P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='1' AND B( 1)='0' )then
          cVar1S20S69P017N062P014P035(0) <='1';
          else
          cVar1S20S69P017N062P014P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='1' AND B( 1)='0' )then
          cVar1S21S69P017N062P014P035(0) <='1';
          else
          cVar1S21S69P017N062P014P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='1' AND B( 1)='1' )then
          cVar1S22S69P017N062P014P035(0) <='1';
          else
          cVar1S22S69P017N062P014P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A(12)='1' AND B( 1)='1' )then
          cVar1S23S69P017N062P014P035(0) <='1';
          else
          cVar1S23S69P017N062P014P035(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='0' )then
          cVar1S24S69N017P066P028P055(0) <='1';
          else
          cVar1S24S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='0' )then
          cVar1S25S69N017P066P028P055(0) <='1';
          else
          cVar1S25S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='0' )then
          cVar1S26S69N017P066P028P055(0) <='1';
          else
          cVar1S26S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='1' )then
          cVar1S27S69N017P066P028P055(0) <='1';
          else
          cVar1S27S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='1' )then
          cVar1S28S69N017P066P028P055(0) <='1';
          else
          cVar1S28S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='1' )then
          cVar1S29S69N017P066P028P055(0) <='1';
          else
          cVar1S29S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='0' AND D(11)='1' )then
          cVar1S30S69N017P066P028P055(0) <='1';
          else
          cVar1S30S69N017P066P028P055(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND B(13)='1' AND B(12)='0' )then
          cVar1S31S69N017P066P028P030(0) <='1';
          else
          cVar1S31S69N017P066P028P030(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='1' )then
          cVar1S32S69N017N066P047P049(0) <='1';
          else
          cVar1S32S69N017N066P047P049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='1' )then
          cVar1S33S69N017N066P047P049(0) <='1';
          else
          cVar1S33S69N017N066P047P049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='1' )then
          cVar1S34S69N017N066P047P049(0) <='1';
          else
          cVar1S34S69N017N066P047P049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='0' )then
          cVar1S35S69N017N066P047N049(0) <='1';
          else
          cVar1S35S69N017N066P047N049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='0' )then
          cVar1S36S69N017N066P047N049(0) <='1';
          else
          cVar1S36S69N017N066P047N049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='1' AND E(13)='0' )then
          cVar1S37S69N017N066P047N049(0) <='1';
          else
          cVar1S37S69N017N066P047N049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='1' )then
          cVar1S38S69N017N066N047P023(0) <='1';
          else
          cVar1S38S69N017N066N047P023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='1' )then
          cVar1S39S69N017N066N047P023(0) <='1';
          else
          cVar1S39S69N017N066N047P023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='0' )then
          cVar1S40S69N017N066N047N023(0) <='1';
          else
          cVar1S40S69N017N066N047N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='0' )then
          cVar1S41S69N017N066N047N023(0) <='1';
          else
          cVar1S41S69N017N066N047N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='0' )then
          cVar1S42S69N017N066N047N023(0) <='1';
          else
          cVar1S42S69N017N066N047N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND D(13)='0' AND B( 7)='0' )then
          cVar1S43S69N017N066N047N023(0) <='1';
          else
          cVar1S43S69N017N066N047N023(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='0' AND A(14)='1' )then
          cVar1S0S70P017P014P062P010(0) <='1';
          else
          cVar1S0S70P017P014P062P010(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='0' AND A(14)='1' )then
          cVar1S1S70P017P014P062P010(0) <='1';
          else
          cVar1S1S70P017P014P062P010(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='0' AND A(14)='0' )then
          cVar1S2S70P017P014P062N010(0) <='1';
          else
          cVar1S2S70P017P014P062N010(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='0' AND A(14)='0' )then
          cVar1S3S70P017P014P062N010(0) <='1';
          else
          cVar1S3S70P017P014P062N010(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='0' AND A(14)='0' )then
          cVar1S4S70P017P014P062N010(0) <='1';
          else
          cVar1S4S70P017P014P062N010(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='1' AND B( 2)='1' )then
          cVar1S5S70P017P014P062P033(0) <='1';
          else
          cVar1S5S70P017P014P062P033(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='1' AND B( 2)='0' )then
          cVar1S6S70P017P014P062N033(0) <='1';
          else
          cVar1S6S70P017P014P062N033(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND D( 1)='1' AND B( 2)='0' )then
          cVar1S7S70P017P014P062N033(0) <='1';
          else
          cVar1S7S70P017P014P062N033(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND A(13)='0' AND E(15)='1' )then
          cVar1S8S70P017P014P012P041nsss(0) <='1';
          else
          cVar1S8S70P017P014P012P041nsss(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND A(13)='0' AND E(15)='0' )then
          cVar1S9S70P017P014P012N041(0) <='1';
          else
          cVar1S9S70P017P014P012N041(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND A(13)='1' AND E(13)='0' )then
          cVar1S10S70P017P014P012P049(0) <='1';
          else
          cVar1S10S70P017P014P012P049(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND A(13)='1' AND E(13)='0' )then
          cVar1S11S70P017P014P012P049(0) <='1';
          else
          cVar1S11S70P017P014P012P049(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND A(13)='1' AND E(13)='0' )then
          cVar1S12S70P017P014P012P049(0) <='1';
          else
          cVar1S12S70P017P014P012P049(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='1' )then
          cVar1S13S70N017P066P044P032(0) <='1';
          else
          cVar1S13S70N017P066P044P032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='1' )then
          cVar1S14S70N017P066P044P032(0) <='1';
          else
          cVar1S14S70N017P066P044P032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='1' )then
          cVar1S15S70N017P066P044P032(0) <='1';
          else
          cVar1S15S70N017P066P044P032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='0' )then
          cVar1S16S70N017P066P044N032(0) <='1';
          else
          cVar1S16S70N017P066P044N032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='0' )then
          cVar1S17S70N017P066P044N032(0) <='1';
          else
          cVar1S17S70N017P066P044N032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='0' AND B(11)='0' )then
          cVar1S18S70N017P066P044N032(0) <='1';
          else
          cVar1S18S70N017P066P044N032(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='1' AND E(14)='0' )then
          cVar1S19S70N017P066P044P045(0) <='1';
          else
          cVar1S19S70N017P066P044P045(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='1' AND E(14)='0' )then
          cVar1S20S70N017P066P044P045(0) <='1';
          else
          cVar1S20S70N017P066P044P045(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='0' AND E( 6)='1' AND E(14)='0' )then
          cVar1S21S70N017P066P044P045(0) <='1';
          else
          cVar1S21S70N017P066P044P045(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='0' AND B(10)='1' )then
          cVar1S22S70N017P066P004P034(0) <='1';
          else
          cVar1S22S70N017P066P004P034(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='0' AND B(10)='0' )then
          cVar1S23S70N017P066P004N034(0) <='1';
          else
          cVar1S23S70N017P066P004N034(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='0' AND B(10)='0' )then
          cVar1S24S70N017P066P004N034(0) <='1';
          else
          cVar1S24S70N017P066P004N034(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='1' AND E(10)='1' )then
          cVar1S25S70N017P066P004P061nsss(0) <='1';
          else
          cVar1S25S70N017P066P004P061nsss(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='1' AND E(10)='0' )then
          cVar1S26S70N017P066P004N061(0) <='1';
          else
          cVar1S26S70N017P066P004N061(0) <='0';
          end if;
        if(A( 1)='0' AND D( 0)='1' AND A(17)='1' AND E(10)='0' )then
          cVar1S27S70N017P066P004N061(0) <='1';
          else
          cVar1S27S70N017P066P004N061(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='0' )then
          cVar1S0S71P067P015P018P069(0) <='1';
          else
          cVar1S0S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='0' )then
          cVar1S1S71P067P015P018P069(0) <='1';
          else
          cVar1S1S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='0' )then
          cVar1S2S71P067P015P018P069(0) <='1';
          else
          cVar1S2S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='0' )then
          cVar1S3S71P067P015P018P069(0) <='1';
          else
          cVar1S3S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='1' )then
          cVar1S4S71P067P015P018P069(0) <='1';
          else
          cVar1S4S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='1' AND E( 8)='1' )then
          cVar1S5S71P067P015P018P069(0) <='1';
          else
          cVar1S5S71P067P015P018P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='1' )then
          cVar1S6S71P067P015N018P002(0) <='1';
          else
          cVar1S6S71P067P015N018P002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='1' )then
          cVar1S7S71P067P015N018P002(0) <='1';
          else
          cVar1S7S71P067P015N018P002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='0' )then
          cVar1S8S71P067P015N018N002(0) <='1';
          else
          cVar1S8S71P067P015N018N002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='0' )then
          cVar1S9S71P067P015N018N002(0) <='1';
          else
          cVar1S9S71P067P015N018N002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='0' )then
          cVar1S10S71P067P015N018N002(0) <='1';
          else
          cVar1S10S71P067P015N018N002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='0' AND A(10)='0' AND A(18)='0' )then
          cVar1S11S71P067P015N018N002(0) <='1';
          else
          cVar1S11S71P067P015N018N002(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='1' )then
          cVar1S12S71P067P015P017P069(0) <='1';
          else
          cVar1S12S71P067P015P017P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='1' )then
          cVar1S13S71P067P015P017P069(0) <='1';
          else
          cVar1S13S71P067P015P017P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='1' )then
          cVar1S14S71P067P015P017P069(0) <='1';
          else
          cVar1S14S71P067P015P017P069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='0' )then
          cVar1S15S71P067P015P017N069(0) <='1';
          else
          cVar1S15S71P067P015P017N069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='0' )then
          cVar1S16S71P067P015P017N069(0) <='1';
          else
          cVar1S16S71P067P015P017N069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='0' )then
          cVar1S17S71P067P015P017N069(0) <='1';
          else
          cVar1S17S71P067P015P017N069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='1' AND E( 8)='0' )then
          cVar1S18S71P067P015P017N069(0) <='1';
          else
          cVar1S18S71P067P015P017N069(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='0' AND B(14)='0' )then
          cVar1S19S71P067P015N017P026(0) <='1';
          else
          cVar1S19S71P067P015N017P026(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='0' AND B(14)='0' )then
          cVar1S20S71P067P015N017P026(0) <='1';
          else
          cVar1S20S71P067P015N017P026(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='0' AND B(14)='0' )then
          cVar1S21S71P067P015N017P026(0) <='1';
          else
          cVar1S21S71P067P015N017P026(0) <='0';
          end if;
        if(D( 8)='0' AND A( 2)='1' AND A( 1)='0' AND B(14)='1' )then
          cVar1S22S71P067P015N017P026(0) <='1';
          else
          cVar1S22S71P067P015N017P026(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='1' AND E(11)='0' AND B( 0)='0' )then
          cVar1S23S71P067P001P057P037(0) <='1';
          else
          cVar1S23S71P067P001P057P037(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='1' AND E(11)='0' AND B( 0)='0' )then
          cVar1S24S71P067P001P057P037(0) <='1';
          else
          cVar1S24S71P067P001P057P037(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='1' AND E(11)='0' AND B( 0)='0' )then
          cVar1S25S71P067P001P057P037(0) <='1';
          else
          cVar1S25S71P067P001P057P037(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='1' AND E(11)='0' AND B( 0)='1' )then
          cVar1S26S71P067P001P057P037(0) <='1';
          else
          cVar1S26S71P067P001P057P037(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='1' AND D( 3)='0' )then
          cVar1S27S71P067N001P003P054(0) <='1';
          else
          cVar1S27S71P067N001P003P054(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='1' AND D( 3)='0' )then
          cVar1S28S71P067N001P003P054(0) <='1';
          else
          cVar1S28S71P067N001P003P054(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='0' AND E(14)='0' )then
          cVar1S29S71P067N001N003P045(0) <='1';
          else
          cVar1S29S71P067N001N003P045(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='0' AND E(14)='0' )then
          cVar1S30S71P067N001N003P045(0) <='1';
          else
          cVar1S30S71P067N001N003P045(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='0' AND E(14)='1' )then
          cVar1S31S71P067N001N003P045(0) <='1';
          else
          cVar1S31S71P067N001N003P045(0) <='0';
          end if;
        if(D( 8)='1' AND A( 9)='0' AND A( 8)='0' AND E(14)='1' )then
          cVar1S32S71P067N001N003P045(0) <='1';
          else
          cVar1S32S71P067N001N003P045(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='1' AND E( 3)='0' )then
          cVar1S0S72P069P045P052P056(0) <='1';
          else
          cVar1S0S72P069P045P052P056(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='0' )then
          cVar1S1S72P069P045N052P029(0) <='1';
          else
          cVar1S1S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='0' )then
          cVar1S2S72P069P045N052P029(0) <='1';
          else
          cVar1S2S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='0' )then
          cVar1S3S72P069P045N052P029(0) <='1';
          else
          cVar1S3S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='1' )then
          cVar1S4S72P069P045N052P029(0) <='1';
          else
          cVar1S4S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='1' )then
          cVar1S5S72P069P045N052P029(0) <='1';
          else
          cVar1S5S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='1' )then
          cVar1S6S72P069P045N052P029(0) <='1';
          else
          cVar1S6S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='0' AND E( 4)='0' AND B( 4)='1' )then
          cVar1S7S72P069P045N052P029(0) <='1';
          else
          cVar1S7S72P069P045N052P029(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='1' AND A(10)='0' AND A(16)='1' )then
          cVar1S8S72P069P045P018P006nsss(0) <='1';
          else
          cVar1S8S72P069P045P018P006nsss(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='1' AND A(10)='0' AND A(16)='0' )then
          cVar1S9S72P069P045P018N006(0) <='1';
          else
          cVar1S9S72P069P045P018N006(0) <='0';
          end if;
        if(E( 8)='1' AND E(14)='1' AND A(10)='1' AND D(13)='0' )then
          cVar1S10S72P069P045P018P047(0) <='1';
          else
          cVar1S10S72P069P045P018P047(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='1' AND A(15)='1' )then
          cVar1S11S72N069P015P027P008(0) <='1';
          else
          cVar1S11S72N069P015P027P008(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='1' AND A(15)='1' )then
          cVar1S12S72N069P015P027P008(0) <='1';
          else
          cVar1S12S72N069P015P027P008(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='1' AND A(15)='0' )then
          cVar1S13S72N069P015P027N008(0) <='1';
          else
          cVar1S13S72N069P015P027N008(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='1' AND A(15)='0' )then
          cVar1S14S72N069P015P027N008(0) <='1';
          else
          cVar1S14S72N069P015P027N008(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='0' AND A(19)='0' )then
          cVar1S15S72N069P015N027P000(0) <='1';
          else
          cVar1S15S72N069P015N027P000(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='0' AND A(19)='0' )then
          cVar1S16S72N069P015N027P000(0) <='1';
          else
          cVar1S16S72N069P015N027P000(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='0' AND A(19)='0' )then
          cVar1S17S72N069P015N027P000(0) <='1';
          else
          cVar1S17S72N069P015N027P000(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='0' AND A(19)='1' )then
          cVar1S18S72N069P015N027P000(0) <='1';
          else
          cVar1S18S72N069P015N027P000(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='0' AND B( 5)='0' AND A(19)='1' )then
          cVar1S19S72N069P015N027P000(0) <='1';
          else
          cVar1S19S72N069P015N027P000(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='1' AND B(14)='0' )then
          cVar1S20S72N069P015P028P026(0) <='1';
          else
          cVar1S20S72N069P015P028P026(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='1' AND B(14)='0' )then
          cVar1S21S72N069P015P028P026(0) <='1';
          else
          cVar1S21S72N069P015P028P026(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='1' AND B(14)='0' )then
          cVar1S22S72N069P015P028P026(0) <='1';
          else
          cVar1S22S72N069P015P028P026(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='0' AND B(17)='0' )then
          cVar1S23S72N069P015N028P020(0) <='1';
          else
          cVar1S23S72N069P015N028P020(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='0' AND B(17)='0' )then
          cVar1S24S72N069P015N028P020(0) <='1';
          else
          cVar1S24S72N069P015N028P020(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='0' AND B(17)='0' )then
          cVar1S25S72N069P015N028P020(0) <='1';
          else
          cVar1S25S72N069P015N028P020(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='0' AND B(17)='1' )then
          cVar1S26S72N069P015N028P020(0) <='1';
          else
          cVar1S26S72N069P015N028P020(0) <='0';
          end if;
        if(E( 8)='0' AND A( 2)='1' AND B(13)='0' AND B(17)='1' )then
          cVar1S27S72N069P015N028P020(0) <='1';
          else
          cVar1S27S72N069P015N028P020(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='1' AND E(14)='1' )then
          cVar1S0S73P016P038P043P045(0) <='1';
          else
          cVar1S0S73P016P038P043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='1' AND E(14)='0' )then
          cVar1S1S73P016P038P043N045(0) <='1';
          else
          cVar1S1S73P016P038P043N045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='1' AND E(14)='0' )then
          cVar1S2S73P016P038P043N045(0) <='1';
          else
          cVar1S2S73P016P038P043N045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='1' AND E(14)='0' )then
          cVar1S3S73P016P038P043N045(0) <='1';
          else
          cVar1S3S73P016P038P043N045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S4S73P016P038N043P045(0) <='1';
          else
          cVar1S4S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S5S73P016P038N043P045(0) <='1';
          else
          cVar1S5S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S6S73P016P038N043P045(0) <='1';
          else
          cVar1S6S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S7S73P016P038N043P045(0) <='1';
          else
          cVar1S7S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S8S73P016P038N043P045(0) <='1';
          else
          cVar1S8S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S9S73P016P038N043P045(0) <='1';
          else
          cVar1S9S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S10S73P016P038N043P045(0) <='1';
          else
          cVar1S10S73P016P038N043P045(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='1' AND B( 2)='0' AND A(10)='0' )then
          cVar1S11S73P016P038P033P018(0) <='1';
          else
          cVar1S11S73P016P038P033P018(0) <='0';
          end if;
        if(A(11)='1' AND D( 7)='1' AND B( 2)='0' AND A(10)='0' )then
          cVar1S12S73P016P038P033P018(0) <='1';
          else
          cVar1S12S73P016P038P033P018(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='0' )then
          cVar1S13S73N016P036P027P014(0) <='1';
          else
          cVar1S13S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='0' )then
          cVar1S14S73N016P036P027P014(0) <='1';
          else
          cVar1S14S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='0' )then
          cVar1S15S73N016P036P027P014(0) <='1';
          else
          cVar1S15S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='1' )then
          cVar1S16S73N016P036P027P014(0) <='1';
          else
          cVar1S16S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='1' )then
          cVar1S17S73N016P036P027P014(0) <='1';
          else
          cVar1S17S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='1' AND A(12)='1' )then
          cVar1S18S73N016P036P027P014(0) <='1';
          else
          cVar1S18S73N016P036P027P014(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='1' )then
          cVar1S19S73N016P036N027P038(0) <='1';
          else
          cVar1S19S73N016P036N027P038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='1' )then
          cVar1S20S73N016P036N027P038(0) <='1';
          else
          cVar1S20S73N016P036N027P038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='1' )then
          cVar1S21S73N016P036N027P038(0) <='1';
          else
          cVar1S21S73N016P036N027P038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='0' )then
          cVar1S22S73N016P036N027N038(0) <='1';
          else
          cVar1S22S73N016P036N027N038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='0' )then
          cVar1S23S73N016P036N027N038(0) <='1';
          else
          cVar1S23S73N016P036N027N038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='0' )then
          cVar1S24S73N016P036N027N038(0) <='1';
          else
          cVar1S24S73N016P036N027N038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='0' AND B( 5)='0' AND D( 7)='0' )then
          cVar1S25S73N016P036N027N038(0) <='1';
          else
          cVar1S25S73N016P036N027N038(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='1' AND E(14)='0' AND E( 0)='0' )then
          cVar1S26S73N016P036P045P068(0) <='1';
          else
          cVar1S26S73N016P036P045P068(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='1' AND E(14)='0' AND E( 0)='0' )then
          cVar1S27S73N016P036P045P068(0) <='1';
          else
          cVar1S27S73N016P036P045P068(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='1' AND E(14)='0' AND E( 0)='1' )then
          cVar1S28S73N016P036P045P068(0) <='1';
          else
          cVar1S28S73N016P036P045P068(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='1' AND E(14)='0' AND E( 0)='1' )then
          cVar1S29S73N016P036P045P068(0) <='1';
          else
          cVar1S29S73N016P036P045P068(0) <='0';
          end if;
        if(A(11)='0' AND B( 9)='1' AND E(14)='1' AND D(14)='1' )then
          cVar1S30S73N016P036P045P043(0) <='1';
          else
          cVar1S30S73N016P036P045P043(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar1S0S74P016P053P035P026(0) <='1';
          else
          cVar1S0S74P016P053P035P026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar1S1S74P016P053P035P026(0) <='1';
          else
          cVar1S1S74P016P053P035P026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar1S2S74P016P053P035P026(0) <='1';
          else
          cVar1S2S74P016P053P035P026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar1S3S74P016P053P035P026(0) <='1';
          else
          cVar1S3S74P016P053P035P026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='0' )then
          cVar1S4S74P016P053P035N026(0) <='1';
          else
          cVar1S4S74P016P053P035N026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='0' )then
          cVar1S5S74P016P053P035N026(0) <='1';
          else
          cVar1S5S74P016P053P035N026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='0' AND B(14)='0' )then
          cVar1S6S74P016P053P035N026(0) <='1';
          else
          cVar1S6S74P016P053P035N026(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='1' AND E( 4)='1' )then
          cVar1S7S74P016P053P035P052(0) <='1';
          else
          cVar1S7S74P016P053P035P052(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='1' AND E( 4)='1' )then
          cVar1S8S74P016P053P035P052(0) <='1';
          else
          cVar1S8S74P016P053P035P052(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='1' AND E( 4)='1' )then
          cVar1S9S74P016P053P035P052(0) <='1';
          else
          cVar1S9S74P016P053P035P052(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='0' AND B( 1)='1' AND E( 4)='0' )then
          cVar1S10S74P016P053P035N052(0) <='1';
          else
          cVar1S10S74P016P053P035N052(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='1' AND A( 0)='0' )then
          cVar1S11S74P016P053P030P019(0) <='1';
          else
          cVar1S11S74P016P053P030P019(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='1' AND A( 0)='0' )then
          cVar1S12S74P016P053P030P019(0) <='1';
          else
          cVar1S12S74P016P053P030P019(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='1' AND A( 0)='0' )then
          cVar1S13S74P016P053P030P019(0) <='1';
          else
          cVar1S13S74P016P053P030P019(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='0' AND D(10)='0' )then
          cVar1S14S74P016P053N030P059(0) <='1';
          else
          cVar1S14S74P016P053N030P059(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='0' AND D(10)='0' )then
          cVar1S15S74P016P053N030P059(0) <='1';
          else
          cVar1S15S74P016P053N030P059(0) <='0';
          end if;
        if(A(11)='0' AND E(12)='1' AND B(12)='0' AND D(10)='1' )then
          cVar1S16S74P016P053N030P059(0) <='1';
          else
          cVar1S16S74P016P053N030P059(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='1' AND D( 1)='1' )then
          cVar1S17S74P016P043P062nsss(0) <='1';
          else
          cVar1S17S74P016P043P062nsss(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='1' AND D( 1)='0' AND B(16)='1' )then
          cVar1S18S74P016P043N062P022nsss(0) <='1';
          else
          cVar1S18S74P016P043N062P022nsss(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='1' AND D( 1)='0' AND B(16)='0' )then
          cVar1S19S74P016P043N062N022(0) <='1';
          else
          cVar1S19S74P016P043N062N022(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='1' AND D( 1)='0' AND B(16)='0' )then
          cVar1S20S74P016P043N062N022(0) <='1';
          else
          cVar1S20S74P016P043N062N022(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='0' AND E( 3)='0' )then
          cVar1S21S74P016N043P038P056(0) <='1';
          else
          cVar1S21S74P016N043P038P056(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='0' AND E( 3)='0' )then
          cVar1S22S74P016N043P038P056(0) <='1';
          else
          cVar1S22S74P016N043P038P056(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='0' AND E( 3)='0' )then
          cVar1S23S74P016N043P038P056(0) <='1';
          else
          cVar1S23S74P016N043P038P056(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='0' AND E( 3)='1' )then
          cVar1S24S74P016N043P038P056(0) <='1';
          else
          cVar1S24S74P016N043P038P056(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='0' AND E( 3)='1' )then
          cVar1S25S74P016N043P038P056(0) <='1';
          else
          cVar1S25S74P016N043P038P056(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='1' AND B( 2)='0' )then
          cVar1S26S74P016N043P038P033(0) <='1';
          else
          cVar1S26S74P016N043P038P033(0) <='0';
          end if;
        if(A(11)='1' AND D(14)='0' AND D( 7)='1' AND B( 2)='0' )then
          cVar1S27S74P016N043P038P033(0) <='1';
          else
          cVar1S27S74P016N043P038P033(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='1' AND B(14)='0' AND A(16)='1' )then
          cVar1S0S75P064P027P026P006(0) <='1';
          else
          cVar1S0S75P064P027P026P006(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='1' AND B(14)='0' AND A(16)='1' )then
          cVar1S1S75P064P027P026P006(0) <='1';
          else
          cVar1S1S75P064P027P026P006(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='1' AND B(14)='0' AND A(16)='0' )then
          cVar1S2S75P064P027P026N006(0) <='1';
          else
          cVar1S2S75P064P027P026N006(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='1' AND B(14)='0' AND A(16)='0' )then
          cVar1S3S75P064P027P026N006(0) <='1';
          else
          cVar1S3S75P064P027P026N006(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='1' AND B(14)='1' AND A(14)='0' )then
          cVar1S4S75P064P027P026P010(0) <='1';
          else
          cVar1S4S75P064P027P026P010(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='0' )then
          cVar1S5S75P064N027P060P054(0) <='1';
          else
          cVar1S5S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='0' )then
          cVar1S6S75P064N027P060P054(0) <='1';
          else
          cVar1S6S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='0' )then
          cVar1S7S75P064N027P060P054(0) <='1';
          else
          cVar1S7S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='0' )then
          cVar1S8S75P064N027P060P054(0) <='1';
          else
          cVar1S8S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='1' )then
          cVar1S9S75P064N027P060P054(0) <='1';
          else
          cVar1S9S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='1' AND D( 3)='1' )then
          cVar1S10S75P064N027P060P054(0) <='1';
          else
          cVar1S10S75P064N027P060P054(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='0' )then
          cVar1S11S75P064N027N060P062(0) <='1';
          else
          cVar1S11S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='0' )then
          cVar1S12S75P064N027N060P062(0) <='1';
          else
          cVar1S12S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='1' )then
          cVar1S13S75P064N027N060P062(0) <='1';
          else
          cVar1S13S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='1' )then
          cVar1S14S75P064N027N060P062(0) <='1';
          else
          cVar1S14S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='1' )then
          cVar1S15S75P064N027N060P062(0) <='1';
          else
          cVar1S15S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='0' AND B( 5)='0' AND E( 2)='0' AND D( 1)='1' )then
          cVar1S16S75P064N027N060P062(0) <='1';
          else
          cVar1S16S75P064N027N060P062(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='1' AND D( 5)='0' AND D( 2)='1' )then
          cVar1S17S75P064P003P046P058(0) <='1';
          else
          cVar1S17S75P064P003P046P058(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='1' AND D( 5)='0' AND D( 2)='0' )then
          cVar1S18S75P064P003P046N058(0) <='1';
          else
          cVar1S18S75P064P003P046N058(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='1' AND D( 5)='0' AND D( 2)='0' )then
          cVar1S19S75P064P003P046N058(0) <='1';
          else
          cVar1S19S75P064P003P046N058(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='1' AND D( 5)='0' AND D( 2)='0' )then
          cVar1S20S75P064P003P046N058(0) <='1';
          else
          cVar1S20S75P064P003P046N058(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar1S21S75P064N003P018P065(0) <='1';
          else
          cVar1S21S75P064N003P018P065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar1S22S75P064N003P018P065(0) <='1';
          else
          cVar1S22S75P064N003P018P065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar1S23S75P064N003P018P065(0) <='1';
          else
          cVar1S23S75P064N003P018P065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar1S24S75P064N003P018P065(0) <='1';
          else
          cVar1S24S75P064N003P018P065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S25S75P064N003P018N065(0) <='1';
          else
          cVar1S25S75P064N003P018N065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S26S75P064N003P018N065(0) <='1';
          else
          cVar1S26S75P064N003P018N065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='1' AND E( 9)='0' )then
          cVar1S27S75P064N003P018N065(0) <='1';
          else
          cVar1S27S75P064N003P018N065(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S28S75P064N003N018P013(0) <='1';
          else
          cVar1S28S75P064N003N018P013(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S29S75P064N003N018P013(0) <='1';
          else
          cVar1S29S75P064N003N018P013(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S30S75P064N003N018P013(0) <='1';
          else
          cVar1S30S75P064N003N018P013(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar1S31S75P064N003N018N013(0) <='1';
          else
          cVar1S31S75P064N003N018N013(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar1S32S75P064N003N018N013(0) <='1';
          else
          cVar1S32S75P064N003N018N013(0) <='0';
          end if;
        if(E( 1)='1' AND A( 8)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar1S33S75P064N003N018N013(0) <='1';
          else
          cVar1S33S75P064N003N018N013(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='0' )then
          cVar1S0S76P016P060P056P067(0) <='1';
          else
          cVar1S0S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='0' )then
          cVar1S1S76P016P060P056P067(0) <='1';
          else
          cVar1S1S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='0' )then
          cVar1S2S76P016P060P056P067(0) <='1';
          else
          cVar1S2S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='1' )then
          cVar1S3S76P016P060P056P067(0) <='1';
          else
          cVar1S3S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='1' )then
          cVar1S4S76P016P060P056P067(0) <='1';
          else
          cVar1S4S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='0' AND D( 8)='1' )then
          cVar1S5S76P016P060P056P067(0) <='1';
          else
          cVar1S5S76P016P060P056P067(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='1' AND A( 4)='0' )then
          cVar1S6S76P016P060P056P011(0) <='1';
          else
          cVar1S6S76P016P060P056P011(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='1' AND A( 4)='0' )then
          cVar1S7S76P016P060P056P011(0) <='1';
          else
          cVar1S7S76P016P060P056P011(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='0' AND E( 3)='1' AND A( 4)='1' )then
          cVar1S8S76P016P060P056P011(0) <='1';
          else
          cVar1S8S76P016P060P056P011(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='0' AND E( 1)='0' )then
          cVar1S9S76P016P060P015P064(0) <='1';
          else
          cVar1S9S76P016P060P015P064(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='0' AND E( 1)='0' )then
          cVar1S10S76P016P060P015P064(0) <='1';
          else
          cVar1S10S76P016P060P015P064(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='0' AND E( 1)='0' )then
          cVar1S11S76P016P060P015P064(0) <='1';
          else
          cVar1S11S76P016P060P015P064(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='0' AND E( 1)='1' )then
          cVar1S12S76P016P060P015P064(0) <='1';
          else
          cVar1S12S76P016P060P015P064(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='0' AND E( 1)='1' )then
          cVar1S13S76P016P060P015P064(0) <='1';
          else
          cVar1S13S76P016P060P015P064(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='1' AND B(17)='0' )then
          cVar1S14S76P016P060P015P020(0) <='1';
          else
          cVar1S14S76P016P060P015P020(0) <='0';
          end if;
        if(A(11)='1' AND E( 2)='1' AND A( 2)='1' AND B(17)='0' )then
          cVar1S15S76P016P060P015P020(0) <='1';
          else
          cVar1S15S76P016P060P015P020(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='1' )then
          cVar1S16S76N016P064P048P062(0) <='1';
          else
          cVar1S16S76N016P064P048P062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='1' )then
          cVar1S17S76N016P064P048P062(0) <='1';
          else
          cVar1S17S76N016P064P048P062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='1' )then
          cVar1S18S76N016P064P048P062(0) <='1';
          else
          cVar1S18S76N016P064P048P062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='0' )then
          cVar1S19S76N016P064P048N062(0) <='1';
          else
          cVar1S19S76N016P064P048N062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='0' )then
          cVar1S20S76N016P064P048N062(0) <='1';
          else
          cVar1S20S76N016P064P048N062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='0' AND D( 1)='0' )then
          cVar1S21S76N016P064P048N062(0) <='1';
          else
          cVar1S21S76N016P064P048N062(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='1' AND D( 2)='0' )then
          cVar1S22S76N016P064P048P058(0) <='1';
          else
          cVar1S22S76N016P064P048P058(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='1' AND E( 5)='1' AND D( 2)='0' )then
          cVar1S23S76N016P064P048P058(0) <='1';
          else
          cVar1S23S76N016P064P048P058(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='1' AND A(16)='1' )then
          cVar1S24S76N016N064P027P006(0) <='1';
          else
          cVar1S24S76N016N064P027P006(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='1' AND A(16)='0' )then
          cVar1S25S76N016N064P027N006(0) <='1';
          else
          cVar1S25S76N016N064P027N006(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='1' AND A(16)='0' )then
          cVar1S26S76N016N064P027N006(0) <='1';
          else
          cVar1S26S76N016N064P027N006(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='0' )then
          cVar1S27S76N016N064N027P057(0) <='1';
          else
          cVar1S27S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='0' )then
          cVar1S28S76N016N064N027P057(0) <='1';
          else
          cVar1S28S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='0' )then
          cVar1S29S76N016N064N027P057(0) <='1';
          else
          cVar1S29S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='1' )then
          cVar1S30S76N016N064N027P057(0) <='1';
          else
          cVar1S30S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='1' )then
          cVar1S31S76N016N064N027P057(0) <='1';
          else
          cVar1S31S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='1' )then
          cVar1S32S76N016N064N027P057(0) <='1';
          else
          cVar1S32S76N016N064N027P057(0) <='0';
          end if;
        if(A(11)='0' AND E( 1)='0' AND B( 5)='0' AND E(11)='1' )then
          cVar1S33S76N016N064N027P057(0) <='1';
          else
          cVar1S33S76N016N064N027P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='0' )then
          cVar1S0S77P035P053P016P057(0) <='1';
          else
          cVar1S0S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='0' )then
          cVar1S1S77P035P053P016P057(0) <='1';
          else
          cVar1S1S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='0' )then
          cVar1S2S77P035P053P016P057(0) <='1';
          else
          cVar1S2S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='0' )then
          cVar1S3S77P035P053P016P057(0) <='1';
          else
          cVar1S3S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='1' )then
          cVar1S4S77P035P053P016P057(0) <='1';
          else
          cVar1S4S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='0' AND E(11)='1' )then
          cVar1S5S77P035P053P016P057(0) <='1';
          else
          cVar1S5S77P035P053P016P057(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='1' AND B(13)='0' )then
          cVar1S6S77P035P053P016P028(0) <='1';
          else
          cVar1S6S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='1' AND B(13)='0' )then
          cVar1S7S77P035P053P016P028(0) <='1';
          else
          cVar1S7S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='1' AND B(13)='0' )then
          cVar1S8S77P035P053P016P028(0) <='1';
          else
          cVar1S8S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='1' AND B(13)='0' )then
          cVar1S9S77P035P053P016P028(0) <='1';
          else
          cVar1S9S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='0' AND A(11)='1' AND B(13)='1' )then
          cVar1S10S77P035P053P016P028(0) <='1';
          else
          cVar1S10S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='1' AND B(13)='1' )then
          cVar1S11S77P035P053P016P028(0) <='1';
          else
          cVar1S11S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='1' AND B(13)='1' )then
          cVar1S12S77P035P053P016P028(0) <='1';
          else
          cVar1S12S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='1' AND B(13)='1' )then
          cVar1S13S77P035P053P016P028(0) <='1';
          else
          cVar1S13S77P035P053P016P028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='1' AND B(13)='0' )then
          cVar1S14S77P035P053P016N028(0) <='1';
          else
          cVar1S14S77P035P053P016N028(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='0' AND D(10)='0' )then
          cVar1S15S77P035P053N016P059(0) <='1';
          else
          cVar1S15S77P035P053N016P059(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='0' AND D(10)='0' )then
          cVar1S16S77P035P053N016P059(0) <='1';
          else
          cVar1S16S77P035P053N016P059(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='0' AND D(10)='0' )then
          cVar1S17S77P035P053N016P059(0) <='1';
          else
          cVar1S17S77P035P053N016P059(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='0' AND D(10)='0' )then
          cVar1S18S77P035P053N016P059(0) <='1';
          else
          cVar1S18S77P035P053N016P059(0) <='0';
          end if;
        if(B( 1)='0' AND E(12)='1' AND A(11)='0' AND D(10)='1' )then
          cVar1S19S77P035P053N016P059(0) <='1';
          else
          cVar1S19S77P035P053N016P059(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='1' AND A(13)='0' AND B( 4)='1' )then
          cVar1S20S77P035P052P012P029nsss(0) <='1';
          else
          cVar1S20S77P035P052P012P029nsss(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='1' AND A(13)='0' AND B( 4)='0' )then
          cVar1S21S77P035P052P012N029(0) <='1';
          else
          cVar1S21S77P035P052P012N029(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='1' AND A(13)='0' AND B( 4)='0' )then
          cVar1S22S77P035P052P012N029(0) <='1';
          else
          cVar1S22S77P035P052P012N029(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='1' AND A(13)='1' AND E( 1)='1' )then
          cVar1S23S77P035P052P012P064nsss(0) <='1';
          else
          cVar1S23S77P035P052P012P064nsss(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='1' AND B( 2)='0' )then
          cVar1S24S77P035N052P046P033(0) <='1';
          else
          cVar1S24S77P035N052P046P033(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='1' AND B( 2)='0' )then
          cVar1S25S77P035N052P046P033(0) <='1';
          else
          cVar1S25S77P035N052P046P033(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='0' AND D(12)='1' )then
          cVar1S26S77P035N052N046P051(0) <='1';
          else
          cVar1S26S77P035N052N046P051(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='0' AND D(12)='1' )then
          cVar1S27S77P035N052N046P051(0) <='1';
          else
          cVar1S27S77P035N052N046P051(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='0' AND D(12)='0' )then
          cVar1S28S77P035N052N046N051(0) <='1';
          else
          cVar1S28S77P035N052N046N051(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='0' AND D(12)='0' )then
          cVar1S29S77P035N052N046N051(0) <='1';
          else
          cVar1S29S77P035N052N046N051(0) <='0';
          end if;
        if(B( 1)='1' AND E( 4)='0' AND D( 5)='0' AND D(12)='0' )then
          cVar1S30S77P035N052N046N051(0) <='1';
          else
          cVar1S30S77P035N052N046N051(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='1' AND B( 9)='1' )then
          cVar1S0S78P035P064P052P036nsss(0) <='1';
          else
          cVar1S0S78P035P064P052P036nsss(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='1' AND B( 9)='0' )then
          cVar1S1S78P035P064P052N036(0) <='1';
          else
          cVar1S1S78P035P064P052N036(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='1' AND B( 9)='0' )then
          cVar1S2S78P035P064P052N036(0) <='1';
          else
          cVar1S2S78P035P064P052N036(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='1' AND B( 9)='0' )then
          cVar1S3S78P035P064P052N036(0) <='1';
          else
          cVar1S3S78P035P064P052N036(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='1' )then
          cVar1S4S78P035P064N052P037(0) <='1';
          else
          cVar1S4S78P035P064N052P037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='1' )then
          cVar1S5S78P035P064N052P037(0) <='1';
          else
          cVar1S5S78P035P064N052P037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='1' )then
          cVar1S6S78P035P064N052P037(0) <='1';
          else
          cVar1S6S78P035P064N052P037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='1' )then
          cVar1S7S78P035P064N052P037(0) <='1';
          else
          cVar1S7S78P035P064N052P037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='0' )then
          cVar1S8S78P035P064N052N037(0) <='1';
          else
          cVar1S8S78P035P064N052N037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='0' )then
          cVar1S9S78P035P064N052N037(0) <='1';
          else
          cVar1S9S78P035P064N052N037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND E( 4)='0' AND B( 0)='0' )then
          cVar1S10S78P035P064N052N037(0) <='1';
          else
          cVar1S10S78P035P064N052N037(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='0' AND A( 9)='0' )then
          cVar1S11S78P035N064P012P001(0) <='1';
          else
          cVar1S11S78P035N064P012P001(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='0' AND A( 9)='0' )then
          cVar1S12S78P035N064P012P001(0) <='1';
          else
          cVar1S12S78P035N064P012P001(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='0' AND A( 9)='0' )then
          cVar1S13S78P035N064P012P001(0) <='1';
          else
          cVar1S13S78P035N064P012P001(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='1' AND B( 9)='1' )then
          cVar1S14S78P035N064P012P036(0) <='1';
          else
          cVar1S14S78P035N064P012P036(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='1' AND B( 9)='1' )then
          cVar1S15S78P035N064P012P036(0) <='1';
          else
          cVar1S15S78P035N064P012P036(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND A(13)='1' AND B( 9)='0' )then
          cVar1S16S78P035N064P012N036(0) <='1';
          else
          cVar1S16S78P035N064P012N036(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='0' AND A( 2)='1' )then
          cVar1S17S78N035P016P064P015(0) <='1';
          else
          cVar1S17S78N035P016P064P015(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='0' AND A( 2)='1' )then
          cVar1S18S78N035P016P064P015(0) <='1';
          else
          cVar1S18S78N035P016P064P015(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='0' AND A( 2)='0' )then
          cVar1S19S78N035P016P064N015(0) <='1';
          else
          cVar1S19S78N035P016P064N015(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='0' AND A( 2)='0' )then
          cVar1S20S78N035P016P064N015(0) <='1';
          else
          cVar1S20S78N035P016P064N015(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='0' AND A( 2)='0' )then
          cVar1S21S78N035P016P064N015(0) <='1';
          else
          cVar1S21S78N035P016P064N015(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S22S78N035P016P064P048(0) <='1';
          else
          cVar1S22S78N035P016P064P048(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S23S78N035P016P064P048(0) <='1';
          else
          cVar1S23S78N035P016P064P048(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='0' )then
          cVar1S24S78N035P016P064P048(0) <='1';
          else
          cVar1S24S78N035P016P064P048(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='0' AND E( 1)='1' AND E( 5)='1' )then
          cVar1S25S78N035P016P064P048(0) <='1';
          else
          cVar1S25S78N035P016P064P048(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='1' AND A(17)='0' )then
          cVar1S26S78N035P016P053P004(0) <='1';
          else
          cVar1S26S78N035P016P053P004(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='1' AND A(17)='0' )then
          cVar1S27S78N035P016P053P004(0) <='1';
          else
          cVar1S27S78N035P016P053P004(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='1' AND A(17)='0' )then
          cVar1S28S78N035P016P053P004(0) <='1';
          else
          cVar1S28S78N035P016P053P004(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='0' AND B(13)='0' )then
          cVar1S29S78N035P016N053P028(0) <='1';
          else
          cVar1S29S78N035P016N053P028(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='0' AND B(13)='0' )then
          cVar1S30S78N035P016N053P028(0) <='1';
          else
          cVar1S30S78N035P016N053P028(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='0' AND B(13)='0' )then
          cVar1S31S78N035P016N053P028(0) <='1';
          else
          cVar1S31S78N035P016N053P028(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='0' AND B(13)='0' )then
          cVar1S32S78N035P016N053P028(0) <='1';
          else
          cVar1S32S78N035P016N053P028(0) <='0';
          end if;
        if(B( 1)='0' AND A(11)='1' AND E(12)='0' AND B(13)='1' )then
          cVar1S33S78N035P016N053P028(0) <='1';
          else
          cVar1S33S78N035P016N053P028(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='1' AND E(12)='0' )then
          cVar1S0S79P064P035P052P053nsss(0) <='1';
          else
          cVar1S0S79P064P035P052P053nsss(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='0' AND D(11)='0' )then
          cVar1S1S79P064P035N052P055(0) <='1';
          else
          cVar1S1S79P064P035N052P055(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='0' AND D(11)='0' )then
          cVar1S2S79P064P035N052P055(0) <='1';
          else
          cVar1S2S79P064P035N052P055(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='0' AND D(11)='0' )then
          cVar1S3S79P064P035N052P055(0) <='1';
          else
          cVar1S3S79P064P035N052P055(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='0' AND D(11)='1' )then
          cVar1S4S79P064P035N052P055(0) <='1';
          else
          cVar1S4S79P064P035N052P055(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='1' AND E( 4)='0' AND D(11)='1' )then
          cVar1S5S79P064P035N052P055(0) <='1';
          else
          cVar1S5S79P064P035N052P055(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S6S79P064N035P051P048(0) <='1';
          else
          cVar1S6S79P064N035P051P048(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S7S79P064N035P051P048(0) <='1';
          else
          cVar1S7S79P064N035P051P048(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S8S79P064N035P051P048(0) <='1';
          else
          cVar1S8S79P064N035P051P048(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S9S79P064N035P051P048(0) <='1';
          else
          cVar1S9S79P064N035P051P048(0) <='0';
          end if;
        if(E( 1)='1' AND B( 1)='0' AND D(12)='1' AND E( 8)='0' )then
          cVar1S10S79P064N035P051P069(0) <='1';
          else
          cVar1S10S79P064N035P051P069(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='1' )then
          cVar1S11S79N064P035P016P026(0) <='1';
          else
          cVar1S11S79N064P035P016P026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='1' )then
          cVar1S12S79N064P035P016P026(0) <='1';
          else
          cVar1S12S79N064P035P016P026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='0' )then
          cVar1S13S79N064P035P016N026(0) <='1';
          else
          cVar1S13S79N064P035P016N026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='0' )then
          cVar1S14S79N064P035P016N026(0) <='1';
          else
          cVar1S14S79N064P035P016N026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='0' )then
          cVar1S15S79N064P035P016N026(0) <='1';
          else
          cVar1S15S79N064P035P016N026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='0' AND B(14)='0' )then
          cVar1S16S79N064P035P016N026(0) <='1';
          else
          cVar1S16S79N064P035P016N026(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='1' AND E( 4)='1' )then
          cVar1S17S79N064P035P016P052(0) <='1';
          else
          cVar1S17S79N064P035P016P052(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='1' AND E( 4)='1' )then
          cVar1S18S79N064P035P016P052(0) <='1';
          else
          cVar1S18S79N064P035P016P052(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='1' AND E( 4)='1' )then
          cVar1S19S79N064P035P016P052(0) <='1';
          else
          cVar1S19S79N064P035P016P052(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='1' AND E( 4)='0' )then
          cVar1S20S79N064P035P016N052(0) <='1';
          else
          cVar1S20S79N064P035P016N052(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='0' AND A(11)='1' AND E( 4)='0' )then
          cVar1S21S79N064P035P016N052(0) <='1';
          else
          cVar1S21S79N064P035P016N052(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='0' AND A(11)='1' )then
          cVar1S22S79N064P035P013P016(0) <='1';
          else
          cVar1S22S79N064P035P013P016(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='0' AND A(11)='0' )then
          cVar1S23S79N064P035P013N016(0) <='1';
          else
          cVar1S23S79N064P035P013N016(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='0' AND A(11)='0' )then
          cVar1S24S79N064P035P013N016(0) <='1';
          else
          cVar1S24S79N064P035P013N016(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='0' AND A(11)='0' )then
          cVar1S25S79N064P035P013N016(0) <='1';
          else
          cVar1S25S79N064P035P013N016(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='1' AND B(12)='1' )then
          cVar1S26S79N064P035P013P030(0) <='1';
          else
          cVar1S26S79N064P035P013P030(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='1' AND B(12)='1' )then
          cVar1S27S79N064P035P013P030(0) <='1';
          else
          cVar1S27S79N064P035P013P030(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='1' AND B(12)='0' )then
          cVar1S28S79N064P035P013N030(0) <='1';
          else
          cVar1S28S79N064P035P013N030(0) <='0';
          end if;
        if(E( 1)='0' AND B( 1)='1' AND A( 3)='1' AND B(12)='0' )then
          cVar1S29S79N064P035P013N030(0) <='1';
          else
          cVar1S29S79N064P035P013N030(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='0' )then
          cVar1S0S80P037P034P057P058(0) <='1';
          else
          cVar1S0S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='0' )then
          cVar1S1S80P037P034P057P058(0) <='1';
          else
          cVar1S1S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='0' )then
          cVar1S2S80P037P034P057P058(0) <='1';
          else
          cVar1S2S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='1' )then
          cVar1S3S80P037P034P057P058(0) <='1';
          else
          cVar1S3S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='1' )then
          cVar1S4S80P037P034P057P058(0) <='1';
          else
          cVar1S4S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='0' AND D( 2)='1' )then
          cVar1S5S80P037P034P057P058(0) <='1';
          else
          cVar1S5S80P037P034P057P058(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='1' AND A(12)='1' )then
          cVar1S6S80P037P034P057P014(0) <='1';
          else
          cVar1S6S80P037P034P057P014(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='1' AND A(12)='1' )then
          cVar1S7S80P037P034P057P014(0) <='1';
          else
          cVar1S7S80P037P034P057P014(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='1' AND E(11)='1' AND A(12)='0' )then
          cVar1S8S80P037P034P057N014(0) <='1';
          else
          cVar1S8S80P037P034P057N014(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='1' AND A(13)='0' )then
          cVar1S9S80P037N034P017P012(0) <='1';
          else
          cVar1S9S80P037N034P017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='1' AND A(13)='0' )then
          cVar1S10S80P037N034P017P012(0) <='1';
          else
          cVar1S10S80P037N034P017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='1' AND A(13)='0' )then
          cVar1S11S80P037N034P017P012(0) <='1';
          else
          cVar1S11S80P037N034P017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='1' AND A(13)='1' )then
          cVar1S12S80P037N034P017P012(0) <='1';
          else
          cVar1S12S80P037N034P017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='1' AND A(13)='1' )then
          cVar1S13S80P037N034P017P012(0) <='1';
          else
          cVar1S13S80P037N034P017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='1' )then
          cVar1S14S80P037N034N017P012(0) <='1';
          else
          cVar1S14S80P037N034N017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='1' )then
          cVar1S15S80P037N034N017P012(0) <='1';
          else
          cVar1S15S80P037N034N017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='1' )then
          cVar1S16S80P037N034N017P012(0) <='1';
          else
          cVar1S16S80P037N034N017P012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='0' )then
          cVar1S17S80P037N034N017N012(0) <='1';
          else
          cVar1S17S80P037N034N017N012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='0' )then
          cVar1S18S80P037N034N017N012(0) <='1';
          else
          cVar1S18S80P037N034N017N012(0) <='0';
          end if;
        if(B( 0)='0' AND B(10)='0' AND A( 1)='0' AND A(13)='0' )then
          cVar1S19S80P037N034N017N012(0) <='1';
          else
          cVar1S19S80P037N034N017N012(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='1' AND B( 4)='1' )then
          cVar1S20S80P037P015P052P029nsss(0) <='1';
          else
          cVar1S20S80P037P015P052P029nsss(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='1' AND B( 4)='0' )then
          cVar1S21S80P037P015P052N029(0) <='1';
          else
          cVar1S21S80P037P015P052N029(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='0' AND B( 6)='1' )then
          cVar1S22S80P037P015N052P025(0) <='1';
          else
          cVar1S22S80P037P015N052P025(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='0' AND B( 6)='1' )then
          cVar1S23S80P037P015N052P025(0) <='1';
          else
          cVar1S23S80P037P015N052P025(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='0' AND B( 6)='0' )then
          cVar1S24S80P037P015N052N025(0) <='1';
          else
          cVar1S24S80P037P015N052N025(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='1' AND E( 4)='0' AND B( 6)='0' )then
          cVar1S25S80P037P015N052N025(0) <='1';
          else
          cVar1S25S80P037P015N052N025(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='1' AND D(11)='0' )then
          cVar1S26S80P037N015P018P055(0) <='1';
          else
          cVar1S26S80P037N015P018P055(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='1' AND D(11)='0' )then
          cVar1S27S80P037N015P018P055(0) <='1';
          else
          cVar1S27S80P037N015P018P055(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='1' AND D(11)='0' )then
          cVar1S28S80P037N015P018P055(0) <='1';
          else
          cVar1S28S80P037N015P018P055(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='1' AND D(11)='0' )then
          cVar1S29S80P037N015P018P055(0) <='1';
          else
          cVar1S29S80P037N015P018P055(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='1' AND D(11)='1' )then
          cVar1S30S80P037N015P018P055(0) <='1';
          else
          cVar1S30S80P037N015P018P055(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='0' )then
          cVar1S31S80P037N015N018P034(0) <='1';
          else
          cVar1S31S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='0' )then
          cVar1S32S80P037N015N018P034(0) <='1';
          else
          cVar1S32S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='0' )then
          cVar1S33S80P037N015N018P034(0) <='1';
          else
          cVar1S33S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='0' )then
          cVar1S34S80P037N015N018P034(0) <='1';
          else
          cVar1S34S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='1' )then
          cVar1S35S80P037N015N018P034(0) <='1';
          else
          cVar1S35S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='1' )then
          cVar1S36S80P037N015N018P034(0) <='1';
          else
          cVar1S36S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='1' AND A( 2)='0' AND A(10)='0' AND B(10)='1' )then
          cVar1S37S80P037N015N018P034(0) <='1';
          else
          cVar1S37S80P037N015N018P034(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='0' )then
          cVar1S0S81P037P032P017P056(0) <='1';
          else
          cVar1S0S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='0' )then
          cVar1S1S81P037P032P017P056(0) <='1';
          else
          cVar1S1S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='0' )then
          cVar1S2S81P037P032P017P056(0) <='1';
          else
          cVar1S2S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='1' )then
          cVar1S3S81P037P032P017P056(0) <='1';
          else
          cVar1S3S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='1' )then
          cVar1S4S81P037P032P017P056(0) <='1';
          else
          cVar1S4S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='0' AND E( 3)='1' )then
          cVar1S5S81P037P032P017P056(0) <='1';
          else
          cVar1S5S81P037P032P017P056(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='1' AND B( 9)='1' )then
          cVar1S6S81P037P032P017P036(0) <='1';
          else
          cVar1S6S81P037P032P017P036(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='1' AND B( 9)='1' )then
          cVar1S7S81P037P032P017P036(0) <='1';
          else
          cVar1S7S81P037P032P017P036(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='1' AND B( 9)='0' )then
          cVar1S8S81P037P032P017N036(0) <='1';
          else
          cVar1S8S81P037P032P017N036(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='0' AND A( 1)='1' AND B( 9)='0' )then
          cVar1S9S81P037P032P017N036(0) <='1';
          else
          cVar1S9S81P037P032P017N036(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='0' AND B( 3)='0' )then
          cVar1S10S81P037P032P013P031(0) <='1';
          else
          cVar1S10S81P037P032P013P031(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='0' AND B( 3)='0' )then
          cVar1S11S81P037P032P013P031(0) <='1';
          else
          cVar1S11S81P037P032P013P031(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='0' AND B( 3)='1' )then
          cVar1S12S81P037P032P013P031(0) <='1';
          else
          cVar1S12S81P037P032P013P031(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='0' AND B( 3)='1' )then
          cVar1S13S81P037P032P013P031(0) <='1';
          else
          cVar1S13S81P037P032P013P031(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='1' AND D(10)='1' )then
          cVar1S14S81P037P032P013P059(0) <='1';
          else
          cVar1S14S81P037P032P013P059(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='1' AND D(10)='1' )then
          cVar1S15S81P037P032P013P059(0) <='1';
          else
          cVar1S15S81P037P032P013P059(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='1' AND D(10)='1' )then
          cVar1S16S81P037P032P013P059(0) <='1';
          else
          cVar1S16S81P037P032P013P059(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='1' AND D(10)='0' )then
          cVar1S17S81P037P032P013N059(0) <='1';
          else
          cVar1S17S81P037P032P013N059(0) <='0';
          end if;
        if(B( 0)='0' AND B(11)='1' AND A( 3)='1' AND D(10)='0' )then
          cVar1S18S81P037P032P013N059(0) <='1';
          else
          cVar1S18S81P037P032P013N059(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='1' AND A( 3)='1' )then
          cVar1S19S81P037P052P008P013nsss(0) <='1';
          else
          cVar1S19S81P037P052P008P013nsss(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar1S20S81P037P052P008N013(0) <='1';
          else
          cVar1S20S81P037P052P008N013(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar1S21S81P037P052P008N013(0) <='1';
          else
          cVar1S21S81P037P052P008N013(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar1S22S81P037P052P008N013(0) <='1';
          else
          cVar1S22S81P037P052P008N013(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='1' )then
          cVar1S23S81P037P052N008P068(0) <='1';
          else
          cVar1S23S81P037P052N008P068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='1' )then
          cVar1S24S81P037P052N008P068(0) <='1';
          else
          cVar1S24S81P037P052N008P068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='1' )then
          cVar1S25S81P037P052N008P068(0) <='1';
          else
          cVar1S25S81P037P052N008P068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='0' )then
          cVar1S26S81P037P052N008N068(0) <='1';
          else
          cVar1S26S81P037P052N008N068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='0' )then
          cVar1S27S81P037P052N008N068(0) <='1';
          else
          cVar1S27S81P037P052N008N068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='1' AND A(15)='0' AND E( 0)='0' )then
          cVar1S28S81P037P052N008N068(0) <='1';
          else
          cVar1S28S81P037P052N008N068(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='1' AND E( 6)='1' )then
          cVar1S29S81P037N052P025P044nsss(0) <='1';
          else
          cVar1S29S81P037N052P025P044nsss(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='1' AND E( 6)='0' )then
          cVar1S30S81P037N052P025N044(0) <='1';
          else
          cVar1S30S81P037N052P025N044(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='1' AND E( 6)='0' )then
          cVar1S31S81P037N052P025N044(0) <='1';
          else
          cVar1S31S81P037N052P025N044(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='1' )then
          cVar1S32S81P037N052N025P024(0) <='1';
          else
          cVar1S32S81P037N052N025P024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='1' )then
          cVar1S33S81P037N052N025P024(0) <='1';
          else
          cVar1S33S81P037N052N025P024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='1' )then
          cVar1S34S81P037N052N025P024(0) <='1';
          else
          cVar1S34S81P037N052N025P024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='0' )then
          cVar1S35S81P037N052N025N024(0) <='1';
          else
          cVar1S35S81P037N052N025N024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='0' )then
          cVar1S36S81P037N052N025N024(0) <='1';
          else
          cVar1S36S81P037N052N025N024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='0' )then
          cVar1S37S81P037N052N025N024(0) <='1';
          else
          cVar1S37S81P037N052N025N024(0) <='0';
          end if;
        if(B( 0)='1' AND E( 4)='0' AND B( 6)='0' AND B(15)='0' )then
          cVar1S38S81P037N052N025N024(0) <='1';
          else
          cVar1S38S81P037N052N025N024(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S0S82P037P031P054P034(0) <='1';
          else
          cVar1S0S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S1S82P037P031P054P034(0) <='1';
          else
          cVar1S1S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S2S82P037P031P054P034(0) <='1';
          else
          cVar1S2S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='1' )then
          cVar1S3S82P037P031P054P034(0) <='1';
          else
          cVar1S3S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='1' )then
          cVar1S4S82P037P031P054P034(0) <='1';
          else
          cVar1S4S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='0' AND B(10)='1' )then
          cVar1S5S82P037P031P054P034(0) <='1';
          else
          cVar1S5S82P037P031P054P034(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='1' AND E( 9)='1' )then
          cVar1S6S82P037P031P054P065(0) <='1';
          else
          cVar1S6S82P037P031P054P065(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='1' AND E( 9)='0' )then
          cVar1S7S82P037P031P054N065(0) <='1';
          else
          cVar1S7S82P037P031P054N065(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='1' AND E( 9)='0' )then
          cVar1S8S82P037P031P054N065(0) <='1';
          else
          cVar1S8S82P037P031P054N065(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='0' AND D( 3)='1' AND E( 9)='0' )then
          cVar1S9S82P037P031P054N065(0) <='1';
          else
          cVar1S9S82P037P031P054N065(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='1' AND D( 2)='1' AND A( 6)='0' )then
          cVar1S10S82P037P031P058P007(0) <='1';
          else
          cVar1S10S82P037P031P058P007(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='1' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S11S82P037P031N058P054(0) <='1';
          else
          cVar1S11S82P037P031N058P054(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='1' AND D( 2)='0' AND D( 3)='1' )then
          cVar1S12S82P037P031N058P054(0) <='1';
          else
          cVar1S12S82P037P031N058P054(0) <='0';
          end if;
        if(B( 0)='1' AND B( 3)='1' AND D( 2)='0' AND D( 3)='0' )then
          cVar1S13S82P037P031N058N054(0) <='1';
          else
          cVar1S13S82P037P031N058N054(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='1' AND E( 2)='0' )then
          cVar1S14S82N037P017P044P060(0) <='1';
          else
          cVar1S14S82N037P017P044P060(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S15S82N037P017N044P023(0) <='1';
          else
          cVar1S15S82N037P017N044P023(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S16S82N037P017N044P023(0) <='1';
          else
          cVar1S16S82N037P017N044P023(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S17S82N037P017N044P023(0) <='1';
          else
          cVar1S17S82N037P017N044P023(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='0' AND B( 7)='1' )then
          cVar1S18S82N037P017N044P023(0) <='1';
          else
          cVar1S18S82N037P017N044P023(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='1' AND E( 6)='0' AND B( 7)='1' )then
          cVar1S19S82N037P017N044P023(0) <='1';
          else
          cVar1S19S82N037P017N044P023(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='1' AND A( 5)='1' )then
          cVar1S20S82N037N017P029P009(0) <='1';
          else
          cVar1S20S82N037N017P029P009(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='1' AND A( 5)='1' )then
          cVar1S21S82N037N017P029P009(0) <='1';
          else
          cVar1S21S82N037N017P029P009(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='1' AND A( 5)='0' )then
          cVar1S22S82N037N017P029N009(0) <='1';
          else
          cVar1S22S82N037N017P029N009(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='1' AND A( 5)='0' )then
          cVar1S23S82N037N017P029N009(0) <='1';
          else
          cVar1S23S82N037N017P029N009(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='0' AND D( 8)='1' )then
          cVar1S24S82N037N017N029P067(0) <='1';
          else
          cVar1S24S82N037N017N029P067(0) <='0';
          end if;
        if(B( 0)='0' AND A( 1)='0' AND B( 4)='0' AND D( 8)='0' )then
          cVar1S25S82N037N017N029N067(0) <='1';
          else
          cVar1S25S82N037N017N029N067(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S0S83P017P037P000P047(0) <='1';
          else
          cVar1S0S83P017P037P000P047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S1S83P017P037P000P047(0) <='1';
          else
          cVar1S1S83P017P037P000P047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='1' )then
          cVar1S2S83P017P037P000P047(0) <='1';
          else
          cVar1S2S83P017P037P000P047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S3S83P017P037P000N047(0) <='1';
          else
          cVar1S3S83P017P037P000N047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S4S83P017P037P000N047(0) <='1';
          else
          cVar1S4S83P017P037P000N047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='0' AND D(13)='0' )then
          cVar1S5S83P017P037P000N047(0) <='1';
          else
          cVar1S5S83P017P037P000N047(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='1' AND B( 8)='1' )then
          cVar1S6S83P017P037P000P021nsss(0) <='1';
          else
          cVar1S6S83P017P037P000P021nsss(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='0' AND A(19)='1' AND B( 8)='0' )then
          cVar1S7S83P017P037P000N021(0) <='1';
          else
          cVar1S7S83P017P037P000N021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='1' AND A( 8)='1' )then
          cVar1S8S83P017P037P019P003(0) <='1';
          else
          cVar1S8S83P017P037P019P003(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='1' AND A( 8)='0' )then
          cVar1S9S83P017P037P019N003(0) <='1';
          else
          cVar1S9S83P017P037P019N003(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='1' AND A( 8)='0' )then
          cVar1S10S83P017P037P019N003(0) <='1';
          else
          cVar1S10S83P017P037P019N003(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='1' AND A( 8)='0' )then
          cVar1S11S83P017P037P019N003(0) <='1';
          else
          cVar1S11S83P017P037P019N003(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='0' AND A( 9)='0' )then
          cVar1S12S83P017P037N019P001(0) <='1';
          else
          cVar1S12S83P017P037N019P001(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='0' AND A( 9)='0' )then
          cVar1S13S83P017P037N019P001(0) <='1';
          else
          cVar1S13S83P017P037N019P001(0) <='0';
          end if;
        if(A( 1)='0' AND B( 0)='1' AND A( 0)='0' AND A( 9)='0' )then
          cVar1S14S83P017P037N019P001(0) <='1';
          else
          cVar1S14S83P017P037N019P001(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='1' AND E( 2)='0' AND A(14)='0' )then
          cVar1S15S83P017P044P060P010(0) <='1';
          else
          cVar1S15S83P017P044P060P010(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='1' AND E( 2)='0' AND A(14)='1' )then
          cVar1S16S83P017P044P060P010(0) <='1';
          else
          cVar1S16S83P017P044P060P010(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND E( 4)='1' )then
          cVar1S17S83P017N044P023P052(0) <='1';
          else
          cVar1S17S83P017N044P023P052(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND E( 4)='1' )then
          cVar1S18S83P017N044P023P052(0) <='1';
          else
          cVar1S18S83P017N044P023P052(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND E( 4)='0' )then
          cVar1S19S83P017N044P023N052(0) <='1';
          else
          cVar1S19S83P017N044P023N052(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND E( 4)='0' )then
          cVar1S20S83P017N044P023N052(0) <='1';
          else
          cVar1S20S83P017N044P023N052(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND E( 4)='0' )then
          cVar1S21S83P017N044P023N052(0) <='1';
          else
          cVar1S21S83P017N044P023N052(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='1' AND E( 9)='1' )then
          cVar1S22S83P017N044P023P065nsss(0) <='1';
          else
          cVar1S22S83P017N044P023P065nsss(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='1' AND E( 9)='0' )then
          cVar1S23S83P017N044P023N065(0) <='1';
          else
          cVar1S23S83P017N044P023N065(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='0' AND E( 1)='0' )then
          cVar1S0S84P019P018P057P064(0) <='1';
          else
          cVar1S0S84P019P018P057P064(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='0' AND E( 1)='0' )then
          cVar1S1S84P019P018P057P064(0) <='1';
          else
          cVar1S1S84P019P018P057P064(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='0' AND E( 1)='1' )then
          cVar1S2S84P019P018P057P064(0) <='1';
          else
          cVar1S2S84P019P018P057P064(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='0' AND E( 1)='1' )then
          cVar1S3S84P019P018P057P064(0) <='1';
          else
          cVar1S3S84P019P018P057P064(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='0' AND E( 1)='1' )then
          cVar1S4S84P019P018P057P064(0) <='1';
          else
          cVar1S4S84P019P018P057P064(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='1' AND A( 8)='1' )then
          cVar1S5S84P019P018P057P003(0) <='1';
          else
          cVar1S5S84P019P018P057P003(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='1' AND A( 8)='0' )then
          cVar1S6S84P019P018P057N003(0) <='1';
          else
          cVar1S6S84P019P018P057N003(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='1' AND A( 8)='0' )then
          cVar1S7S84P019P018P057N003(0) <='1';
          else
          cVar1S7S84P019P018P057N003(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND E(11)='1' AND A( 8)='0' )then
          cVar1S8S84P019P018P057N003(0) <='1';
          else
          cVar1S8S84P019P018P057N003(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S9S84P019P018P033P014(0) <='1';
          else
          cVar1S9S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S10S84P019P018P033P014(0) <='1';
          else
          cVar1S10S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S11S84P019P018P033P014(0) <='1';
          else
          cVar1S11S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='1' )then
          cVar1S12S84P019P018P033P014(0) <='1';
          else
          cVar1S12S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='1' )then
          cVar1S13S84P019P018P033P014(0) <='1';
          else
          cVar1S13S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='1' )then
          cVar1S14S84P019P018P033P014(0) <='1';
          else
          cVar1S14S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='0' AND A(12)='1' )then
          cVar1S15S84P019P018P033P014(0) <='1';
          else
          cVar1S15S84P019P018P033P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='1' AND A( 3)='1' )then
          cVar1S16S84P019P018P033P013(0) <='1';
          else
          cVar1S16S84P019P018P033P013(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='1' AND A( 3)='1' )then
          cVar1S17S84P019P018P033P013(0) <='1';
          else
          cVar1S17S84P019P018P033P013(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='1' AND A( 3)='1' )then
          cVar1S18S84P019P018P033P013(0) <='1';
          else
          cVar1S18S84P019P018P033P013(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='1' AND A( 3)='0' )then
          cVar1S19S84P019P018P033N013(0) <='1';
          else
          cVar1S19S84P019P018P033N013(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND B( 2)='1' AND A( 3)='0' )then
          cVar1S20S84P019P018P033N013(0) <='1';
          else
          cVar1S20S84P019P018P033N013(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='1' AND E( 1)='0' )then
          cVar1S21S84N019P047P006P064(0) <='1';
          else
          cVar1S21S84N019P047P006P064(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='1' AND E( 1)='0' )then
          cVar1S22S84N019P047P006P064(0) <='1';
          else
          cVar1S22S84N019P047P006P064(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='0' AND D( 0)='0' )then
          cVar1S23S84N019P047N006P066(0) <='1';
          else
          cVar1S23S84N019P047N006P066(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='0' AND D( 0)='0' )then
          cVar1S24S84N019P047N006P066(0) <='1';
          else
          cVar1S24S84N019P047N006P066(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='0' AND D( 0)='0' )then
          cVar1S25S84N019P047N006P066(0) <='1';
          else
          cVar1S25S84N019P047N006P066(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='0' AND D( 0)='1' )then
          cVar1S26S84N019P047N006P066(0) <='1';
          else
          cVar1S26S84N019P047N006P066(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='1' AND A(16)='0' AND D( 0)='1' )then
          cVar1S27S84N019P047N006P066(0) <='1';
          else
          cVar1S27S84N019P047N006P066(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='1' AND E( 6)='0' )then
          cVar1S28S84N019N047P043P044(0) <='1';
          else
          cVar1S28S84N019N047P043P044(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='1' AND E( 6)='0' )then
          cVar1S29S84N019N047P043P044(0) <='1';
          else
          cVar1S29S84N019N047P043P044(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='1' AND E( 6)='0' )then
          cVar1S30S84N019N047P043P044(0) <='1';
          else
          cVar1S30S84N019N047P043P044(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='1' AND E( 6)='1' )then
          cVar1S31S84N019N047P043P044(0) <='1';
          else
          cVar1S31S84N019N047P043P044(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='0' )then
          cVar1S32S84N019N047N043P024(0) <='1';
          else
          cVar1S32S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='0' )then
          cVar1S33S84N019N047N043P024(0) <='1';
          else
          cVar1S33S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='0' )then
          cVar1S34S84N019N047N043P024(0) <='1';
          else
          cVar1S34S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='1' )then
          cVar1S35S84N019N047N043P024(0) <='1';
          else
          cVar1S35S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='1' )then
          cVar1S36S84N019N047N043P024(0) <='1';
          else
          cVar1S36S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(13)='0' AND D(14)='0' AND B(15)='1' )then
          cVar1S37S84N019N047N043P024(0) <='1';
          else
          cVar1S37S84N019N047N043P024(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='0' )then
          cVar1S0S85P019P051P067P007(0) <='1';
          else
          cVar1S0S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='0' )then
          cVar1S1S85P019P051P067P007(0) <='1';
          else
          cVar1S1S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='0' )then
          cVar1S2S85P019P051P067P007(0) <='1';
          else
          cVar1S2S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='1' )then
          cVar1S3S85P019P051P067P007(0) <='1';
          else
          cVar1S3S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='1' )then
          cVar1S4S85P019P051P067P007(0) <='1';
          else
          cVar1S4S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='1' )then
          cVar1S5S85P019P051P067P007(0) <='1';
          else
          cVar1S5S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='1' AND A( 6)='1' )then
          cVar1S6S85P019P051P067P007(0) <='1';
          else
          cVar1S6S85P019P051P067P007(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='0' )then
          cVar1S7S85P019P051N067P001(0) <='1';
          else
          cVar1S7S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='0' )then
          cVar1S8S85P019P051N067P001(0) <='1';
          else
          cVar1S8S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='0' )then
          cVar1S9S85P019P051N067P001(0) <='1';
          else
          cVar1S9S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='0' )then
          cVar1S10S85P019P051N067P001(0) <='1';
          else
          cVar1S10S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='1' )then
          cVar1S11S85P019P051N067P001(0) <='1';
          else
          cVar1S11S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='1' )then
          cVar1S12S85P019P051N067P001(0) <='1';
          else
          cVar1S12S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='0' AND D( 8)='0' AND A( 9)='1' )then
          cVar1S13S85P019P051N067P001(0) <='1';
          else
          cVar1S13S85P019P051N067P001(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='1' AND B( 5)='1' )then
          cVar1S14S85P019P051P008P027nsss(0) <='1';
          else
          cVar1S14S85P019P051P008P027nsss(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='1' AND B( 5)='0' )then
          cVar1S15S85P019P051P008N027(0) <='1';
          else
          cVar1S15S85P019P051P008N027(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='1' AND B( 5)='0' )then
          cVar1S16S85P019P051P008N027(0) <='1';
          else
          cVar1S16S85P019P051P008N027(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='0' AND E(11)='0' )then
          cVar1S17S85P019P051N008P057(0) <='1';
          else
          cVar1S17S85P019P051N008P057(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='0' AND E(11)='0' )then
          cVar1S18S85P019P051N008P057(0) <='1';
          else
          cVar1S18S85P019P051N008P057(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='0' AND E(11)='0' )then
          cVar1S19S85P019P051N008P057(0) <='1';
          else
          cVar1S19S85P019P051N008P057(0) <='0';
          end if;
        if(A( 0)='0' AND D(12)='1' AND A(15)='0' AND E(11)='1' )then
          cVar1S20S85P019P051N008P057(0) <='1';
          else
          cVar1S20S85P019P051N008P057(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='0' )then
          cVar1S21S85P019P018P014P033(0) <='1';
          else
          cVar1S21S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='0' )then
          cVar1S22S85P019P018P014P033(0) <='1';
          else
          cVar1S22S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='0' )then
          cVar1S23S85P019P018P014P033(0) <='1';
          else
          cVar1S23S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='1' )then
          cVar1S24S85P019P018P014P033(0) <='1';
          else
          cVar1S24S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='1' )then
          cVar1S25S85P019P018P014P033(0) <='1';
          else
          cVar1S25S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='0' AND B( 2)='1' )then
          cVar1S26S85P019P018P014P033(0) <='1';
          else
          cVar1S26S85P019P018P014P033(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='1' AND B( 7)='1' )then
          cVar1S27S85P019P018P014P023(0) <='1';
          else
          cVar1S27S85P019P018P014P023(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='1' AND B( 7)='0' )then
          cVar1S28S85P019P018P014N023(0) <='1';
          else
          cVar1S28S85P019P018P014N023(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='1' AND B( 7)='0' )then
          cVar1S29S85P019P018P014N023(0) <='1';
          else
          cVar1S29S85P019P018P014N023(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='1' AND B( 7)='0' )then
          cVar1S30S85P019P018P014N023(0) <='1';
          else
          cVar1S30S85P019P018P014N023(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND A(12)='1' AND B( 7)='0' )then
          cVar1S31S85P019P018P014N023(0) <='1';
          else
          cVar1S31S85P019P018P014N023(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='1' AND A(13)='1' )then
          cVar1S32S85P019N018P033P012(0) <='1';
          else
          cVar1S32S85P019N018P033P012(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='1' AND A(13)='1' )then
          cVar1S33S85P019N018P033P012(0) <='1';
          else
          cVar1S33S85P019N018P033P012(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='1' AND A(13)='0' )then
          cVar1S34S85P019N018P033N012(0) <='1';
          else
          cVar1S34S85P019N018P033N012(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='1' AND A(13)='0' )then
          cVar1S35S85P019N018P033N012(0) <='1';
          else
          cVar1S35S85P019N018P033N012(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='1' )then
          cVar1S36S85P019N018N033P010(0) <='1';
          else
          cVar1S36S85P019N018N033P010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='1' )then
          cVar1S37S85P019N018N033P010(0) <='1';
          else
          cVar1S37S85P019N018N033P010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='1' )then
          cVar1S38S85P019N018N033P010(0) <='1';
          else
          cVar1S38S85P019N018N033P010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='0' )then
          cVar1S39S85P019N018N033N010(0) <='1';
          else
          cVar1S39S85P019N018N033N010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='0' )then
          cVar1S40S85P019N018N033N010(0) <='1';
          else
          cVar1S40S85P019N018N033N010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 2)='0' AND A(14)='0' )then
          cVar1S41S85P019N018N033N010(0) <='1';
          else
          cVar1S41S85P019N018N033N010(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='1' )then
          cVar1S0S86P019P018P036P014(0) <='1';
          else
          cVar1S0S86P019P018P036P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='1' )then
          cVar1S1S86P019P018P036P014(0) <='1';
          else
          cVar1S1S86P019P018P036P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='1' )then
          cVar1S2S86P019P018P036P014(0) <='1';
          else
          cVar1S2S86P019P018P036P014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='0' )then
          cVar1S3S86P019P018P036N014(0) <='1';
          else
          cVar1S3S86P019P018P036N014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='0' )then
          cVar1S4S86P019P018P036N014(0) <='1';
          else
          cVar1S4S86P019P018P036N014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='1' AND A(12)='0' )then
          cVar1S5S86P019P018P036N014(0) <='1';
          else
          cVar1S5S86P019P018P036N014(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='0' )then
          cVar1S6S86P019P018N036P069(0) <='1';
          else
          cVar1S6S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='0' )then
          cVar1S7S86P019P018N036P069(0) <='1';
          else
          cVar1S7S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='0' )then
          cVar1S8S86P019P018N036P069(0) <='1';
          else
          cVar1S8S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='0' )then
          cVar1S9S86P019P018N036P069(0) <='1';
          else
          cVar1S9S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='1' )then
          cVar1S10S86P019P018N036P069(0) <='1';
          else
          cVar1S10S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='0' AND B( 9)='0' AND E( 8)='1' )then
          cVar1S11S86P019P018N036P069(0) <='1';
          else
          cVar1S11S86P019P018N036P069(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='1' AND B(12)='1' )then
          cVar1S12S86P019P018P055P030(0) <='1';
          else
          cVar1S12S86P019P018P055P030(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='1' AND B(12)='1' )then
          cVar1S13S86P019P018P055P030(0) <='1';
          else
          cVar1S13S86P019P018P055P030(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='1' AND B(12)='0' )then
          cVar1S14S86P019P018P055N030(0) <='1';
          else
          cVar1S14S86P019P018P055N030(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='1' AND B(12)='0' )then
          cVar1S15S86P019P018P055N030(0) <='1';
          else
          cVar1S15S86P019P018P055N030(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='1' AND B(12)='0' )then
          cVar1S16S86P019P018P055N030(0) <='1';
          else
          cVar1S16S86P019P018P055N030(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='0' AND D( 5)='0' )then
          cVar1S17S86P019P018N055P046(0) <='1';
          else
          cVar1S17S86P019P018N055P046(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='0' AND D( 5)='0' )then
          cVar1S18S86P019P018N055P046(0) <='1';
          else
          cVar1S18S86P019P018N055P046(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='0' AND D( 5)='0' )then
          cVar1S19S86P019P018N055P046(0) <='1';
          else
          cVar1S19S86P019P018N055P046(0) <='0';
          end if;
        if(A( 0)='1' AND A(10)='1' AND D(11)='0' AND D( 5)='1' )then
          cVar1S20S86P019P018N055P046(0) <='1';
          else
          cVar1S20S86P019P018N055P046(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='0' AND B( 3)='0' )then
          cVar1S21S86N019P067P002P031(0) <='1';
          else
          cVar1S21S86N019P067P002P031(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='0' AND B( 3)='0' )then
          cVar1S22S86N019P067P002P031(0) <='1';
          else
          cVar1S22S86N019P067P002P031(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='0' AND B( 3)='0' )then
          cVar1S23S86N019P067P002P031(0) <='1';
          else
          cVar1S23S86N019P067P002P031(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='0' AND B( 3)='1' )then
          cVar1S24S86N019P067P002P031(0) <='1';
          else
          cVar1S24S86N019P067P002P031(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='0' AND B( 3)='1' )then
          cVar1S25S86N019P067P002P031(0) <='1';
          else
          cVar1S25S86N019P067P002P031(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='1' AND E( 1)='1' )then
          cVar1S26S86N019P067P002P064nsss(0) <='1';
          else
          cVar1S26S86N019P067P002P064nsss(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='1' AND A(18)='1' AND E( 1)='0' )then
          cVar1S27S86N019P067P002N064(0) <='1';
          else
          cVar1S27S86N019P067P002N064(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='1' AND A( 4)='1' )then
          cVar1S28S86N019N067P017P011(0) <='1';
          else
          cVar1S28S86N019N067P017P011(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='1' AND A( 4)='1' )then
          cVar1S29S86N019N067P017P011(0) <='1';
          else
          cVar1S29S86N019N067P017P011(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='1' AND A( 4)='0' )then
          cVar1S30S86N019N067P017N011(0) <='1';
          else
          cVar1S30S86N019N067P017N011(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='1' AND A( 4)='0' )then
          cVar1S31S86N019N067P017N011(0) <='1';
          else
          cVar1S31S86N019N067P017N011(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='1' AND A( 4)='0' )then
          cVar1S32S86N019N067P017N011(0) <='1';
          else
          cVar1S32S86N019N067P017N011(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S33S86N019N067N017P069(0) <='1';
          else
          cVar1S33S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S34S86N019N067N017P069(0) <='1';
          else
          cVar1S34S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S35S86N019N067N017P069(0) <='1';
          else
          cVar1S35S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='0' )then
          cVar1S36S86N019N067N017P069(0) <='1';
          else
          cVar1S36S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S37S86N019N067N017P069(0) <='1';
          else
          cVar1S37S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S38S86N019N067N017P069(0) <='1';
          else
          cVar1S38S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S39S86N019N067N017P069(0) <='1';
          else
          cVar1S39S86N019N067N017P069(0) <='0';
          end if;
        if(A( 0)='0' AND D( 8)='0' AND A( 1)='0' AND E( 8)='1' )then
          cVar1S40S86N019N067N017P069(0) <='1';
          else
          cVar1S40S86N019N067N017P069(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='1' )then
          cVar1S0S87P017P002P038P066(0) <='1';
          else
          cVar1S0S87P017P002P038P066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='1' )then
          cVar1S1S87P017P002P038P066(0) <='1';
          else
          cVar1S1S87P017P002P038P066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='1' )then
          cVar1S2S87P017P002P038P066(0) <='1';
          else
          cVar1S2S87P017P002P038P066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='1' )then
          cVar1S3S87P017P002P038P066(0) <='1';
          else
          cVar1S3S87P017P002P038P066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='0' )then
          cVar1S4S87P017P002P038N066(0) <='1';
          else
          cVar1S4S87P017P002P038N066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='0' )then
          cVar1S5S87P017P002P038N066(0) <='1';
          else
          cVar1S5S87P017P002P038N066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='0' AND D( 0)='0' )then
          cVar1S6S87P017P002P038N066(0) <='1';
          else
          cVar1S6S87P017P002P038N066(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='1' AND A(17)='1' )then
          cVar1S7S87P017P002P038P004nsss(0) <='1';
          else
          cVar1S7S87P017P002P038P004nsss(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='0' AND D( 7)='1' AND A(17)='0' )then
          cVar1S8S87P017P002P038N004(0) <='1';
          else
          cVar1S8S87P017P002P038N004(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='1' )then
          cVar1S9S87P017P002P040nsss(0) <='1';
          else
          cVar1S9S87P017P002P040nsss(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='0' AND A( 3)='1' )then
          cVar1S10S87P017P002N040P013(0) <='1';
          else
          cVar1S10S87P017P002N040P013(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='0' AND A( 3)='1' )then
          cVar1S11S87P017P002N040P013(0) <='1';
          else
          cVar1S11S87P017P002N040P013(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='0' AND A( 3)='0' )then
          cVar1S12S87P017P002N040N013(0) <='1';
          else
          cVar1S12S87P017P002N040N013(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='0' AND A( 3)='0' )then
          cVar1S13S87P017P002N040N013(0) <='1';
          else
          cVar1S13S87P017P002N040N013(0) <='0';
          end if;
        if(A( 1)='1' AND A(18)='1' AND E( 7)='0' AND A( 3)='0' )then
          cVar1S14S87P017P002N040N013(0) <='1';
          else
          cVar1S14S87P017P002N040N013(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='1' )then
          cVar1S15S87N017P019P052P003(0) <='1';
          else
          cVar1S15S87N017P019P052P003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='1' )then
          cVar1S16S87N017P019P052P003(0) <='1';
          else
          cVar1S16S87N017P019P052P003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='1' )then
          cVar1S17S87N017P019P052P003(0) <='1';
          else
          cVar1S17S87N017P019P052P003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='0' )then
          cVar1S18S87N017P019P052N003(0) <='1';
          else
          cVar1S18S87N017P019P052N003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='0' )then
          cVar1S19S87N017P019P052N003(0) <='1';
          else
          cVar1S19S87N017P019P052N003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='0' AND A( 8)='0' )then
          cVar1S20S87N017P019P052N003(0) <='1';
          else
          cVar1S20S87N017P019P052N003(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='1' AND A( 5)='1' )then
          cVar1S21S87N017P019P052P009(0) <='1';
          else
          cVar1S21S87N017P019P052P009(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='1' AND A( 5)='1' )then
          cVar1S22S87N017P019P052P009(0) <='1';
          else
          cVar1S22S87N017P019P052P009(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S23S87N017P019P052N009(0) <='1';
          else
          cVar1S23S87N017P019P052N009(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S24S87N017P019P052N009(0) <='1';
          else
          cVar1S24S87N017P019P052N009(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S25S87N017P019P052N009(0) <='1';
          else
          cVar1S25S87N017P019P052N009(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S26S87N017N019P069P067(0) <='1';
          else
          cVar1S26S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S27S87N017N019P069P067(0) <='1';
          else
          cVar1S27S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S28S87N017N019P069P067(0) <='1';
          else
          cVar1S28S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S29S87N017N019P069P067(0) <='1';
          else
          cVar1S29S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S30S87N017N019P069P067(0) <='1';
          else
          cVar1S30S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S31S87N017N019P069P067(0) <='1';
          else
          cVar1S31S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S32S87N017N019P069P067(0) <='1';
          else
          cVar1S32S87N017N019P069P067(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='1' )then
          cVar1S33S87N017N019P069P064(0) <='1';
          else
          cVar1S33S87N017N019P069P064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='1' )then
          cVar1S34S87N017N019P069P064(0) <='1';
          else
          cVar1S34S87N017N019P069P064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='1' )then
          cVar1S35S87N017N019P069P064(0) <='1';
          else
          cVar1S35S87N017N019P069P064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='1' )then
          cVar1S36S87N017N019P069P064(0) <='1';
          else
          cVar1S36S87N017N019P069P064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='0' )then
          cVar1S37S87N017N019P069N064(0) <='1';
          else
          cVar1S37S87N017N019P069N064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='0' )then
          cVar1S38S87N017N019P069N064(0) <='1';
          else
          cVar1S38S87N017N019P069N064(0) <='0';
          end if;
        if(A( 1)='0' AND A( 0)='0' AND E( 8)='1' AND E( 1)='0' )then
          cVar1S39S87N017N019P069N064(0) <='1';
          else
          cVar1S39S87N017N019P069N064(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='0' )then
          cVar1S0S88P014P016P018P012(0) <='1';
          else
          cVar1S0S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='0' )then
          cVar1S1S88P014P016P018P012(0) <='1';
          else
          cVar1S1S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='0' )then
          cVar1S2S88P014P016P018P012(0) <='1';
          else
          cVar1S2S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='1' )then
          cVar1S3S88P014P016P018P012(0) <='1';
          else
          cVar1S3S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='1' )then
          cVar1S4S88P014P016P018P012(0) <='1';
          else
          cVar1S4S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='0' AND A(13)='1' )then
          cVar1S5S88P014P016P018P012(0) <='1';
          else
          cVar1S5S88P014P016P018P012(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='1' )then
          cVar1S6S88P014P016P018P033(0) <='1';
          else
          cVar1S6S88P014P016P018P033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='1' )then
          cVar1S7S88P014P016P018P033(0) <='1';
          else
          cVar1S7S88P014P016P018P033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='1' )then
          cVar1S8S88P014P016P018P033(0) <='1';
          else
          cVar1S8S88P014P016P018P033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='0' )then
          cVar1S9S88P014P016P018N033(0) <='1';
          else
          cVar1S9S88P014P016P018N033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='0' )then
          cVar1S10S88P014P016P018N033(0) <='1';
          else
          cVar1S10S88P014P016P018N033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='0' )then
          cVar1S11S88P014P016P018N033(0) <='1';
          else
          cVar1S11S88P014P016P018N033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='1' AND A(10)='1' AND B( 2)='0' )then
          cVar1S12S88P014P016P018N033(0) <='1';
          else
          cVar1S12S88P014P016P018N033(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar1S13S88P014N016P021P040(0) <='1';
          else
          cVar1S13S88P014N016P021P040(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar1S14S88P014N016P021P040(0) <='1';
          else
          cVar1S14S88P014N016P021P040(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar1S15S88P014N016P021P040(0) <='1';
          else
          cVar1S15S88P014N016P021P040(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='1' AND E( 7)='0' )then
          cVar1S16S88P014N016P021N040(0) <='1';
          else
          cVar1S16S88P014N016P021N040(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='1' AND E( 7)='0' )then
          cVar1S17S88P014N016P021N040(0) <='1';
          else
          cVar1S17S88P014N016P021N040(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='0' AND D( 3)='1' )then
          cVar1S18S88P014N016N021P054(0) <='1';
          else
          cVar1S18S88P014N016N021P054(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='0' AND D( 3)='1' )then
          cVar1S19S88P014N016N021P054(0) <='1';
          else
          cVar1S19S88P014N016N021P054(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='0' AND D( 3)='1' )then
          cVar1S20S88P014N016N021P054(0) <='1';
          else
          cVar1S20S88P014N016N021P054(0) <='0';
          end if;
        if(A(12)='0' AND A(11)='0' AND B( 8)='0' AND D( 3)='0' )then
          cVar1S21S88P014N016N021N054(0) <='1';
          else
          cVar1S21S88P014N016N021N054(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='1' AND A( 0)='1' )then
          cVar1S22S88P014P021P003P019(0) <='1';
          else
          cVar1S22S88P014P021P003P019(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='1' AND A( 0)='0' )then
          cVar1S23S88P014P021P003N019(0) <='1';
          else
          cVar1S23S88P014P021P003N019(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='1' )then
          cVar1S24S88P014P021N003P023(0) <='1';
          else
          cVar1S24S88P014P021N003P023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='1' )then
          cVar1S25S88P014P021N003P023(0) <='1';
          else
          cVar1S25S88P014P021N003P023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='1' )then
          cVar1S26S88P014P021N003P023(0) <='1';
          else
          cVar1S26S88P014P021N003P023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='0' )then
          cVar1S27S88P014P021N003N023(0) <='1';
          else
          cVar1S27S88P014P021N003N023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='0' )then
          cVar1S28S88P014P021N003N023(0) <='1';
          else
          cVar1S28S88P014P021N003N023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A( 8)='0' AND B( 7)='0' )then
          cVar1S29S88P014P021N003N023(0) <='1';
          else
          cVar1S29S88P014P021N003N023(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='1' )then
          cVar1S30S88P014P021P026P037(0) <='1';
          else
          cVar1S30S88P014P021P026P037(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='1' )then
          cVar1S31S88P014P021P026P037(0) <='1';
          else
          cVar1S31S88P014P021P026P037(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='0' )then
          cVar1S32S88P014P021P026N037(0) <='1';
          else
          cVar1S32S88P014P021P026N037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='1' )then
          cVar1S0S89P014P017P015P037(0) <='1';
          else
          cVar1S0S89P014P017P015P037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='1' )then
          cVar1S1S89P014P017P015P037(0) <='1';
          else
          cVar1S1S89P014P017P015P037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='1' )then
          cVar1S2S89P014P017P015P037(0) <='1';
          else
          cVar1S2S89P014P017P015P037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='0' )then
          cVar1S3S89P014P017P015N037(0) <='1';
          else
          cVar1S3S89P014P017P015N037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='0' )then
          cVar1S4S89P014P017P015N037(0) <='1';
          else
          cVar1S4S89P014P017P015N037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='0' AND B( 0)='0' )then
          cVar1S5S89P014P017P015N037(0) <='1';
          else
          cVar1S5S89P014P017P015N037(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='1' AND B(12)='1' )then
          cVar1S6S89P014P017P015P030(0) <='1';
          else
          cVar1S6S89P014P017P015P030(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='1' AND B(12)='1' )then
          cVar1S7S89P014P017P015P030(0) <='1';
          else
          cVar1S7S89P014P017P015P030(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='1' AND B(12)='1' )then
          cVar1S8S89P014P017P015P030(0) <='1';
          else
          cVar1S8S89P014P017P015P030(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='1' AND B(12)='0' )then
          cVar1S9S89P014P017P015N030(0) <='1';
          else
          cVar1S9S89P014P017P015N030(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='1' AND A( 2)='1' AND B(12)='0' )then
          cVar1S10S89P014P017P015N030(0) <='1';
          else
          cVar1S10S89P014P017P015N030(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='1' )then
          cVar1S11S89P014N017P044P015(0) <='1';
          else
          cVar1S11S89P014N017P044P015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='1' )then
          cVar1S12S89P014N017P044P015(0) <='1';
          else
          cVar1S12S89P014N017P044P015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='1' )then
          cVar1S13S89P014N017P044P015(0) <='1';
          else
          cVar1S13S89P014N017P044P015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='0' )then
          cVar1S14S89P014N017P044N015(0) <='1';
          else
          cVar1S14S89P014N017P044N015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='0' )then
          cVar1S15S89P014N017P044N015(0) <='1';
          else
          cVar1S15S89P014N017P044N015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='1' AND A( 2)='0' )then
          cVar1S16S89P014N017P044N015(0) <='1';
          else
          cVar1S16S89P014N017P044N015(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='0' AND B( 5)='1' )then
          cVar1S17S89P014N017N044P027(0) <='1';
          else
          cVar1S17S89P014N017N044P027(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='0' AND B( 5)='1' )then
          cVar1S18S89P014N017N044P027(0) <='1';
          else
          cVar1S18S89P014N017N044P027(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='0' AND B( 5)='0' )then
          cVar1S19S89P014N017N044N027(0) <='1';
          else
          cVar1S19S89P014N017N044N027(0) <='0';
          end if;
        if(A(12)='0' AND A( 1)='0' AND E( 6)='0' AND B( 5)='0' )then
          cVar1S20S89P014N017N044N027(0) <='1';
          else
          cVar1S20S89P014N017N044N027(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='0' AND E( 7)='0' )then
          cVar1S21S89P014P021P012P040(0) <='1';
          else
          cVar1S21S89P014P021P012P040(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='0' AND E( 7)='0' )then
          cVar1S22S89P014P021P012P040(0) <='1';
          else
          cVar1S22S89P014P021P012P040(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='0' AND E( 7)='0' )then
          cVar1S23S89P014P021P012P040(0) <='1';
          else
          cVar1S23S89P014P021P012P040(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='0' AND E( 7)='0' )then
          cVar1S24S89P014P021P012P040(0) <='1';
          else
          cVar1S24S89P014P021P012P040(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='0' AND E( 7)='1' )then
          cVar1S25S89P014P021P012P040(0) <='1';
          else
          cVar1S25S89P014P021P012P040(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='1' AND D(15)='0' )then
          cVar1S26S89P014P021P012P039(0) <='1';
          else
          cVar1S26S89P014P021P012P039(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='1' AND D(15)='0' )then
          cVar1S27S89P014P021P012P039(0) <='1';
          else
          cVar1S27S89P014P021P012P039(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='1' AND D(15)='0' )then
          cVar1S28S89P014P021P012P039(0) <='1';
          else
          cVar1S28S89P014P021P012P039(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='0' AND A(13)='1' AND D(15)='0' )then
          cVar1S29S89P014P021P012P039(0) <='1';
          else
          cVar1S29S89P014P021P012P039(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='1' )then
          cVar1S30S89P014P021P026P037(0) <='1';
          else
          cVar1S30S89P014P021P026P037(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='1' )then
          cVar1S31S89P014P021P026P037(0) <='1';
          else
          cVar1S31S89P014P021P026P037(0) <='0';
          end if;
        if(A(12)='1' AND B( 8)='1' AND B(14)='0' AND B( 0)='0' )then
          cVar1S32S89P014P021P026N037(0) <='1';
          else
          cVar1S32S89P014P021P026N037(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='1' )then
          cVar1S0S90P017P014P019P042(0) <='1';
          else
          cVar1S0S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='1' )then
          cVar1S1S90P017P014P019P042(0) <='1';
          else
          cVar1S1S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='1' )then
          cVar1S2S90P017P014P019P042(0) <='1';
          else
          cVar1S2S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='0' )then
          cVar1S3S90P017P014P019N042(0) <='1';
          else
          cVar1S3S90P017P014P019N042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='0' )then
          cVar1S4S90P017P014P019N042(0) <='1';
          else
          cVar1S4S90P017P014P019N042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='0' AND D( 6)='0' )then
          cVar1S5S90P017P014P019N042(0) <='1';
          else
          cVar1S5S90P017P014P019N042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='1' AND D( 6)='0' )then
          cVar1S6S90P017P014P019P042(0) <='1';
          else
          cVar1S6S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='1' AND D( 6)='0' )then
          cVar1S7S90P017P014P019P042(0) <='1';
          else
          cVar1S7S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='0' AND A( 0)='1' AND D( 6)='1' )then
          cVar1S8S90P017P014P019P042(0) <='1';
          else
          cVar1S8S90P017P014P019P042(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S9S90P017P014P047P024(0) <='1';
          else
          cVar1S9S90P017P014P047P024(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S10S90P017P014P047P024(0) <='1';
          else
          cVar1S10S90P017P014P047P024(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='0' AND B(15)='1' )then
          cVar1S11S90P017P014P047P024(0) <='1';
          else
          cVar1S11S90P017P014P047P024(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='0' AND B(15)='1' )then
          cVar1S12S90P017P014P047P024(0) <='1';
          else
          cVar1S12S90P017P014P047P024(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='0' AND B(15)='1' )then
          cVar1S13S90P017P014P047P024(0) <='1';
          else
          cVar1S13S90P017P014P047P024(0) <='0';
          end if;
        if(A( 1)='1' AND A(12)='1' AND D(13)='1' AND B(15)='1' )then
          cVar1S14S90P017P014P047P024nsss(0) <='1';
          else
          cVar1S14S90P017P014P047P024nsss(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='1' AND B( 6)='1' )then
          cVar1S15S90N017P068P004P025(0) <='1';
          else
          cVar1S15S90N017P068P004P025(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='1' AND B( 6)='0' )then
          cVar1S16S90N017P068P004N025(0) <='1';
          else
          cVar1S16S90N017P068P004N025(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='1' AND B( 6)='0' )then
          cVar1S17S90N017P068P004N025(0) <='1';
          else
          cVar1S17S90N017P068P004N025(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='1' AND B( 6)='0' )then
          cVar1S18S90N017P068P004N025(0) <='1';
          else
          cVar1S18S90N017P068P004N025(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='0' AND B(13)='1' )then
          cVar1S19S90N017P068N004P028(0) <='1';
          else
          cVar1S19S90N017P068N004P028(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='0' AND B(13)='0' )then
          cVar1S20S90N017P068N004N028(0) <='1';
          else
          cVar1S20S90N017P068N004N028(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(17)='0' AND B(13)='0' )then
          cVar1S21S90N017P068N004N028(0) <='1';
          else
          cVar1S21S90N017P068N004N028(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S22S90N017P068P064P062(0) <='1';
          else
          cVar1S22S90N017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S23S90N017P068P064P062(0) <='1';
          else
          cVar1S23S90N017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S24S90N017P068P064P062(0) <='1';
          else
          cVar1S24S90N017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S25S90N017P068P064P062(0) <='1';
          else
          cVar1S25S90N017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S26S90N017P068P064P019(0) <='1';
          else
          cVar1S26S90N017P068P064P019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S27S90N017P068P064P019(0) <='1';
          else
          cVar1S27S90N017P068P064P019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S28S90N017P068P064N019(0) <='1';
          else
          cVar1S28S90N017P068P064N019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S29S90N017P068P064N019(0) <='1';
          else
          cVar1S29S90N017P068P064N019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='1' )then
          cVar1S0S91P017P068P010P004(0) <='1';
          else
          cVar1S0S91P017P068P010P004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='1' )then
          cVar1S1S91P017P068P010P004(0) <='1';
          else
          cVar1S1S91P017P068P010P004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='1' )then
          cVar1S2S91P017P068P010P004(0) <='1';
          else
          cVar1S2S91P017P068P010P004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='0' )then
          cVar1S3S91P017P068P010N004(0) <='1';
          else
          cVar1S3S91P017P068P010N004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='0' )then
          cVar1S4S91P017P068P010N004(0) <='1';
          else
          cVar1S4S91P017P068P010N004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='0' AND A(17)='0' )then
          cVar1S5S91P017P068P010N004(0) <='1';
          else
          cVar1S5S91P017P068P010N004(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='1' AND B( 8)='0' )then
          cVar1S6S91P017P068P010P021(0) <='1';
          else
          cVar1S6S91P017P068P010P021(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='1' AND B( 8)='1' )then
          cVar1S7S91P017P068P010P021(0) <='1';
          else
          cVar1S7S91P017P068P010P021(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='0' AND A(14)='1' AND B( 8)='1' )then
          cVar1S8S91P017P068P010P021(0) <='1';
          else
          cVar1S8S91P017P068P010P021(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S9S91P017P068P064P062(0) <='1';
          else
          cVar1S9S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S10S91P017P068P064P062(0) <='1';
          else
          cVar1S10S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='0' )then
          cVar1S11S91P017P068P064P062(0) <='1';
          else
          cVar1S11S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S12S91P017P068P064P062(0) <='1';
          else
          cVar1S12S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S13S91P017P068P064P062(0) <='1';
          else
          cVar1S13S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S14S91P017P068P064P062(0) <='1';
          else
          cVar1S14S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='0' AND D( 1)='1' )then
          cVar1S15S91P017P068P064P062(0) <='1';
          else
          cVar1S15S91P017P068P064P062(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S16S91P017P068P064P019(0) <='1';
          else
          cVar1S16S91P017P068P064P019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S17S91P017P068P064P019(0) <='1';
          else
          cVar1S17S91P017P068P064P019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S18S91P017P068P064N019(0) <='1';
          else
          cVar1S18S91P017P068P064N019(0) <='0';
          end if;
        if(A( 1)='0' AND E( 0)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S19S91P017P068P064N019(0) <='1';
          else
          cVar1S19S91P017P068P064N019(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='1' AND E( 2)='0' AND A(14)='0' )then
          cVar1S20S91P017P044P060P010(0) <='1';
          else
          cVar1S20S91P017P044P060P010(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='1' AND E( 2)='0' AND A(14)='1' )then
          cVar1S21S91P017P044P060P010(0) <='1';
          else
          cVar1S21S91P017P044P060P010(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='0' )then
          cVar1S22S91P017N044P023P042(0) <='1';
          else
          cVar1S22S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='0' )then
          cVar1S23S91P017N044P023P042(0) <='1';
          else
          cVar1S23S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='0' )then
          cVar1S24S91P017N044P023P042(0) <='1';
          else
          cVar1S24S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='0' )then
          cVar1S25S91P017N044P023P042(0) <='1';
          else
          cVar1S25S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='1' )then
          cVar1S26S91P017N044P023P042(0) <='1';
          else
          cVar1S26S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='0' AND D( 6)='1' )then
          cVar1S27S91P017N044P023P042(0) <='1';
          else
          cVar1S27S91P017N044P023P042(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='1' AND E( 9)='1' )then
          cVar1S28S91P017N044P023P065nsss(0) <='1';
          else
          cVar1S28S91P017N044P023P065nsss(0) <='0';
          end if;
        if(A( 1)='1' AND E( 6)='0' AND B( 7)='1' AND E( 9)='0' )then
          cVar1S29S91P017N044P023N065(0) <='1';
          else
          cVar1S29S91P017N044P023N065(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='0' )then
          cVar1S0S92P017P059P061P013(0) <='1';
          else
          cVar1S0S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='0' )then
          cVar1S1S92P017P059P061P013(0) <='1';
          else
          cVar1S1S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='0' )then
          cVar1S2S92P017P059P061P013(0) <='1';
          else
          cVar1S2S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='0' )then
          cVar1S3S92P017P059P061P013(0) <='1';
          else
          cVar1S3S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='1' )then
          cVar1S4S92P017P059P061P013(0) <='1';
          else
          cVar1S4S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='1' )then
          cVar1S5S92P017P059P061P013(0) <='1';
          else
          cVar1S5S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='1' )then
          cVar1S6S92P017P059P061P013(0) <='1';
          else
          cVar1S6S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='0' AND A( 3)='1' )then
          cVar1S7S92P017P059P061P013(0) <='1';
          else
          cVar1S7S92P017P059P061P013(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='1' AND D( 0)='1' )then
          cVar1S8S92P017P059P061P066(0) <='1';
          else
          cVar1S8S92P017P059P061P066(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='1' AND D( 0)='1' )then
          cVar1S9S92P017P059P061P066(0) <='1';
          else
          cVar1S9S92P017P059P061P066(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='0' AND E(10)='1' AND D( 0)='0' )then
          cVar1S10S92P017P059P061N066(0) <='1';
          else
          cVar1S10S92P017P059P061N066(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='1' AND A(13)='0' )then
          cVar1S11S92P017P059P030P012(0) <='1';
          else
          cVar1S11S92P017P059P030P012(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='1' AND A(13)='0' )then
          cVar1S12S92P017P059P030P012(0) <='1';
          else
          cVar1S12S92P017P059P030P012(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='1' AND A(13)='1' )then
          cVar1S13S92P017P059P030P012(0) <='1';
          else
          cVar1S13S92P017P059P030P012(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='0' AND D(11)='0' )then
          cVar1S14S92P017P059N030P055(0) <='1';
          else
          cVar1S14S92P017P059N030P055(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='0' AND D(11)='0' )then
          cVar1S15S92P017P059N030P055(0) <='1';
          else
          cVar1S15S92P017P059N030P055(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='0' AND D(11)='0' )then
          cVar1S16S92P017P059N030P055(0) <='1';
          else
          cVar1S16S92P017P059N030P055(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='0' AND D(11)='0' )then
          cVar1S17S92P017P059N030P055(0) <='1';
          else
          cVar1S17S92P017P059N030P055(0) <='0';
          end if;
        if(A( 1)='1' AND D(10)='1' AND B(12)='0' AND D(11)='1' )then
          cVar1S18S92P017P059N030P055(0) <='1';
          else
          cVar1S18S92P017P059N030P055(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='1' AND E( 5)='1' )then
          cVar1S19S92N017P006P027P048nsss(0) <='1';
          else
          cVar1S19S92N017P006P027P048nsss(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='1' AND E( 5)='0' )then
          cVar1S20S92N017P006P027N048(0) <='1';
          else
          cVar1S20S92N017P006P027N048(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='1' AND E( 5)='0' )then
          cVar1S21S92N017P006P027N048(0) <='1';
          else
          cVar1S21S92N017P006P027N048(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='0' AND A( 2)='1' )then
          cVar1S22S92N017P006N027P015(0) <='1';
          else
          cVar1S22S92N017P006N027P015(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='0' AND A( 2)='1' )then
          cVar1S23S92N017P006N027P015(0) <='1';
          else
          cVar1S23S92N017P006N027P015(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='0' AND A( 2)='0' )then
          cVar1S24S92N017P006N027N015(0) <='1';
          else
          cVar1S24S92N017P006N027N015(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='1' AND B( 5)='0' AND A( 2)='0' )then
          cVar1S25S92N017P006N027N015(0) <='1';
          else
          cVar1S25S92N017P006N027N015(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='1' AND B(13)='0' )then
          cVar1S26S92N017N006P030P028(0) <='1';
          else
          cVar1S26S92N017N006P030P028(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='1' AND B(13)='0' )then
          cVar1S27S92N017N006P030P028(0) <='1';
          else
          cVar1S27S92N017N006P030P028(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='1' AND B(13)='0' )then
          cVar1S28S92N017N006P030P028(0) <='1';
          else
          cVar1S28S92N017N006P030P028(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='1' AND B(13)='1' )then
          cVar1S29S92N017N006P030P028(0) <='1';
          else
          cVar1S29S92N017N006P030P028(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='1' AND B(13)='1' )then
          cVar1S30S92N017N006P030P028(0) <='1';
          else
          cVar1S30S92N017N006P030P028(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='0' AND A(12)='1' )then
          cVar1S31S92N017N006N030P014(0) <='1';
          else
          cVar1S31S92N017N006N030P014(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='0' AND A(12)='1' )then
          cVar1S32S92N017N006N030P014(0) <='1';
          else
          cVar1S32S92N017N006N030P014(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='0' AND A(12)='1' )then
          cVar1S33S92N017N006N030P014(0) <='1';
          else
          cVar1S33S92N017N006N030P014(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='0' AND A(12)='0' )then
          cVar1S34S92N017N006N030N014(0) <='1';
          else
          cVar1S34S92N017N006N030N014(0) <='0';
          end if;
        if(A( 1)='0' AND A(16)='0' AND B(12)='0' AND A(12)='0' )then
          cVar1S35S92N017N006N030N014(0) <='1';
          else
          cVar1S35S92N017N006N030N014(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='0' )then
          cVar1S0S93P017P030P014P010(0) <='1';
          else
          cVar1S0S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='0' )then
          cVar1S1S93P017P030P014P010(0) <='1';
          else
          cVar1S1S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='0' )then
          cVar1S2S93P017P030P014P010(0) <='1';
          else
          cVar1S2S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='0' )then
          cVar1S3S93P017P030P014P010(0) <='1';
          else
          cVar1S3S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='1' )then
          cVar1S4S93P017P030P014P010(0) <='1';
          else
          cVar1S4S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='1' )then
          cVar1S5S93P017P030P014P010(0) <='1';
          else
          cVar1S5S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='0' AND A(14)='1' )then
          cVar1S6S93P017P030P014P010(0) <='1';
          else
          cVar1S6S93P017P030P014P010(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='1' AND B( 8)='0' )then
          cVar1S7S93P017P030P014P021(0) <='1';
          else
          cVar1S7S93P017P030P014P021(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='1' AND B( 8)='0' )then
          cVar1S8S93P017P030P014P021(0) <='1';
          else
          cVar1S8S93P017P030P014P021(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='1' AND B( 8)='0' )then
          cVar1S9S93P017P030P014P021(0) <='1';
          else
          cVar1S9S93P017P030P014P021(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='1' AND B( 8)='0' )then
          cVar1S10S93P017P030P014P021(0) <='1';
          else
          cVar1S10S93P017P030P014P021(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='0' AND A(12)='1' AND B( 8)='1' )then
          cVar1S11S93P017P030P014P021(0) <='1';
          else
          cVar1S11S93P017P030P014P021(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='1' AND A( 3)='1' )then
          cVar1S12S93P017P030P061P013nsss(0) <='1';
          else
          cVar1S12S93P017P030P061P013nsss(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='1' AND A( 3)='0' )then
          cVar1S13S93P017P030P061N013(0) <='1';
          else
          cVar1S13S93P017P030P061N013(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='1' AND A( 3)='0' )then
          cVar1S14S93P017P030P061N013(0) <='1';
          else
          cVar1S14S93P017P030P061N013(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='0' AND B(11)='0' )then
          cVar1S15S93P017P030N061P032(0) <='1';
          else
          cVar1S15S93P017P030N061P032(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='0' AND B(11)='0' )then
          cVar1S16S93P017P030N061P032(0) <='1';
          else
          cVar1S16S93P017P030N061P032(0) <='0';
          end if;
        if(A( 1)='0' AND B(12)='1' AND E(10)='0' AND B(11)='1' )then
          cVar1S17S93P017P030N061P032(0) <='1';
          else
          cVar1S17S93P017P030N061P032(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='0' )then
          cVar1S18S93P017P013P003P008(0) <='1';
          else
          cVar1S18S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='0' )then
          cVar1S19S93P017P013P003P008(0) <='1';
          else
          cVar1S19S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='0' )then
          cVar1S20S93P017P013P003P008(0) <='1';
          else
          cVar1S20S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='0' )then
          cVar1S21S93P017P013P003P008(0) <='1';
          else
          cVar1S21S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='1' )then
          cVar1S22S93P017P013P003P008(0) <='1';
          else
          cVar1S22S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='0' AND A(15)='1' )then
          cVar1S23S93P017P013P003P008(0) <='1';
          else
          cVar1S23S93P017P013P003P008(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='1' AND E(12)='0' )then
          cVar1S24S93P017P013P003P053(0) <='1';
          else
          cVar1S24S93P017P013P003P053(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='1' AND A( 8)='1' AND E(12)='0' )then
          cVar1S25S93P017P013P003P053(0) <='1';
          else
          cVar1S25S93P017P013P003P053(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='1' AND E( 0)='1' )then
          cVar1S26S93P017N013P003P068(0) <='1';
          else
          cVar1S26S93P017N013P003P068(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='1' AND E( 0)='1' )then
          cVar1S27S93P017N013P003P068(0) <='1';
          else
          cVar1S27S93P017N013P003P068(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='1' AND E( 0)='1' )then
          cVar1S28S93P017N013P003P068(0) <='1';
          else
          cVar1S28S93P017N013P003P068(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='1' AND E( 0)='0' )then
          cVar1S29S93P017N013P003N068(0) <='1';
          else
          cVar1S29S93P017N013P003N068(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='1' AND E( 0)='0' )then
          cVar1S30S93P017N013P003N068(0) <='1';
          else
          cVar1S30S93P017N013P003N068(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='0' AND A(18)='0' )then
          cVar1S31S93P017N013N003P002(0) <='1';
          else
          cVar1S31S93P017N013N003P002(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='0' AND A(18)='0' )then
          cVar1S32S93P017N013N003P002(0) <='1';
          else
          cVar1S32S93P017N013N003P002(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='0' AND A(18)='1' )then
          cVar1S33S93P017N013N003P002(0) <='1';
          else
          cVar1S33S93P017N013N003P002(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='0' AND A(18)='1' )then
          cVar1S34S93P017N013N003P002(0) <='1';
          else
          cVar1S34S93P017N013N003P002(0) <='0';
          end if;
        if(A( 1)='1' AND A( 3)='0' AND A( 8)='0' AND A(18)='1' )then
          cVar1S35S93P017N013N003P002(0) <='1';
          else
          cVar1S35S93P017N013N003P002(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='1' AND A( 6)='0' )then
          cVar1S0S94P013P032P033P007(0) <='1';
          else
          cVar1S0S94P013P032P033P007(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='1' AND A( 6)='0' )then
          cVar1S1S94P013P032P033P007(0) <='1';
          else
          cVar1S1S94P013P032P033P007(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='1' AND A( 6)='1' )then
          cVar1S2S94P013P032P033P007(0) <='1';
          else
          cVar1S2S94P013P032P033P007(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='1' AND A( 6)='1' )then
          cVar1S3S94P013P032P033P007(0) <='1';
          else
          cVar1S3S94P013P032P033P007(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='0' AND B( 3)='1' )then
          cVar1S4S94P013P032N033P031(0) <='1';
          else
          cVar1S4S94P013P032N033P031(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='0' AND B( 3)='1' )then
          cVar1S5S94P013P032N033P031(0) <='1';
          else
          cVar1S5S94P013P032N033P031(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='0' AND B( 3)='0' )then
          cVar1S6S94P013P032N033N031(0) <='1';
          else
          cVar1S6S94P013P032N033N031(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='0' AND B( 3)='0' )then
          cVar1S7S94P013P032N033N031(0) <='1';
          else
          cVar1S7S94P013P032N033N031(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND B( 2)='0' AND B( 3)='0' )then
          cVar1S8S94P013P032N033N031(0) <='1';
          else
          cVar1S8S94P013P032N033N031(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='1' )then
          cVar1S9S94P013P032P061P067(0) <='1';
          else
          cVar1S9S94P013P032P061P067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='1' )then
          cVar1S10S94P013P032P061P067(0) <='1';
          else
          cVar1S10S94P013P032P061P067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S11S94P013P032P061N067(0) <='1';
          else
          cVar1S11S94P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S12S94P013P032P061N067(0) <='1';
          else
          cVar1S12S94P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S13S94P013P032P061N067(0) <='1';
          else
          cVar1S13S94P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='1' )then
          cVar1S14S94P013P032N061P063(0) <='1';
          else
          cVar1S14S94P013P032N061P063(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='0' )then
          cVar1S15S94P013P032N061N063(0) <='1';
          else
          cVar1S15S94P013P032N061N063(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='0' )then
          cVar1S16S94P013P032N061N063(0) <='1';
          else
          cVar1S16S94P013P032N061N063(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='1' )then
          cVar1S17S94N013P017P068P018(0) <='1';
          else
          cVar1S17S94N013P017P068P018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='1' )then
          cVar1S18S94N013P017P068P018(0) <='1';
          else
          cVar1S18S94N013P017P068P018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='1' )then
          cVar1S19S94N013P017P068P018(0) <='1';
          else
          cVar1S19S94N013P017P068P018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S20S94N013P017P068N018(0) <='1';
          else
          cVar1S20S94N013P017P068N018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S21S94N013P017P068N018(0) <='1';
          else
          cVar1S21S94N013P017P068N018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar1S22S94N013P017P068N018(0) <='1';
          else
          cVar1S22S94N013P017P068N018(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='1' AND A( 8)='1' )then
          cVar1S23S94N013P017P068P003(0) <='1';
          else
          cVar1S23S94N013P017P068P003(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='1' AND A( 8)='1' )then
          cVar1S24S94N013P017P068P003(0) <='1';
          else
          cVar1S24S94N013P017P068P003(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='1' AND A( 8)='1' )then
          cVar1S25S94N013P017P068P003(0) <='1';
          else
          cVar1S25S94N013P017P068P003(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='1' AND E( 0)='1' AND A( 8)='0' )then
          cVar1S26S94N013P017P068N003(0) <='1';
          else
          cVar1S26S94N013P017P068N003(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='0' )then
          cVar1S27S94N013N017P015P036(0) <='1';
          else
          cVar1S27S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='0' )then
          cVar1S28S94N013N017P015P036(0) <='1';
          else
          cVar1S28S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='0' )then
          cVar1S29S94N013N017P015P036(0) <='1';
          else
          cVar1S29S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='1' )then
          cVar1S30S94N013N017P015P036(0) <='1';
          else
          cVar1S30S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='1' )then
          cVar1S31S94N013N017P015P036(0) <='1';
          else
          cVar1S31S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='1' AND B( 9)='1' )then
          cVar1S32S94N013N017P015P036(0) <='1';
          else
          cVar1S32S94N013N017P015P036(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='0' AND A( 0)='1' )then
          cVar1S33S94N013N017N015P019(0) <='1';
          else
          cVar1S33S94N013N017N015P019(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='0' AND A( 0)='1' )then
          cVar1S34S94N013N017N015P019(0) <='1';
          else
          cVar1S34S94N013N017N015P019(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='0' AND A( 0)='1' )then
          cVar1S35S94N013N017N015P019(0) <='1';
          else
          cVar1S35S94N013N017N015P019(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='0' AND A( 0)='0' )then
          cVar1S36S94N013N017N015N019(0) <='1';
          else
          cVar1S36S94N013N017N015N019(0) <='0';
          end if;
        if(A( 3)='0' AND A( 1)='0' AND A( 2)='0' AND A( 0)='0' )then
          cVar1S37S94N013N017N015N019(0) <='1';
          else
          cVar1S37S94N013N017N015N019(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='0' )then
          cVar1S0S95P013P032P011P003(0) <='1';
          else
          cVar1S0S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='0' )then
          cVar1S1S95P013P032P011P003(0) <='1';
          else
          cVar1S1S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='0' )then
          cVar1S2S95P013P032P011P003(0) <='1';
          else
          cVar1S2S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='0' )then
          cVar1S3S95P013P032P011P003(0) <='1';
          else
          cVar1S3S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='1' )then
          cVar1S4S95P013P032P011P003(0) <='1';
          else
          cVar1S4S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='0' AND A( 8)='1' )then
          cVar1S5S95P013P032P011P003(0) <='1';
          else
          cVar1S5S95P013P032P011P003(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='1' )then
          cVar1S6S95P013P032P011P036(0) <='1';
          else
          cVar1S6S95P013P032P011P036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='1' )then
          cVar1S7S95P013P032P011P036(0) <='1';
          else
          cVar1S7S95P013P032P011P036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='1' )then
          cVar1S8S95P013P032P011P036(0) <='1';
          else
          cVar1S8S95P013P032P011P036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='0' )then
          cVar1S9S95P013P032P011N036(0) <='1';
          else
          cVar1S9S95P013P032P011N036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='0' )then
          cVar1S10S95P013P032P011N036(0) <='1';
          else
          cVar1S10S95P013P032P011N036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='0' )then
          cVar1S11S95P013P032P011N036(0) <='1';
          else
          cVar1S11S95P013P032P011N036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='0' AND A( 4)='1' AND B( 9)='0' )then
          cVar1S12S95P013P032P011N036(0) <='1';
          else
          cVar1S12S95P013P032P011N036(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='1' )then
          cVar1S13S95P013P032P061P067nsss(0) <='1';
          else
          cVar1S13S95P013P032P061P067nsss(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S14S95P013P032P061N067(0) <='1';
          else
          cVar1S14S95P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S15S95P013P032P061N067(0) <='1';
          else
          cVar1S15S95P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S16S95P013P032P061N067(0) <='1';
          else
          cVar1S16S95P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='1' AND D( 8)='0' )then
          cVar1S17S95P013P032P061N067(0) <='1';
          else
          cVar1S17S95P013P032P061N067(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='1' )then
          cVar1S18S95P013P032N061P063(0) <='1';
          else
          cVar1S18S95P013P032N061P063(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='0' )then
          cVar1S19S95P013P032N061N063(0) <='1';
          else
          cVar1S19S95P013P032N061N063(0) <='0';
          end if;
        if(A( 3)='1' AND B(11)='1' AND E(10)='0' AND D( 9)='0' )then
          cVar1S20S95P013P032N061N063(0) <='1';
          else
          cVar1S20S95P013P032N061N063(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='1' AND A(17)='1' )then
          cVar1S21S95N013P019P041P004(0) <='1';
          else
          cVar1S21S95N013P019P041P004(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='1' AND A(17)='1' )then
          cVar1S22S95N013P019P041P004(0) <='1';
          else
          cVar1S22S95N013P019P041P004(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='1' AND A(17)='0' )then
          cVar1S23S95N013P019P041N004(0) <='1';
          else
          cVar1S23S95N013P019P041N004(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='1' AND A(17)='0' )then
          cVar1S24S95N013P019P041N004(0) <='1';
          else
          cVar1S24S95N013P019P041N004(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='1' AND A(17)='0' )then
          cVar1S25S95N013P019P041N004(0) <='1';
          else
          cVar1S25S95N013P019P041N004(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='0' AND B(17)='0' )then
          cVar1S26S95N013P019N041P020(0) <='1';
          else
          cVar1S26S95N013P019N041P020(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='0' AND B(17)='0' )then
          cVar1S27S95N013P019N041P020(0) <='1';
          else
          cVar1S27S95N013P019N041P020(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='0' AND B(17)='1' )then
          cVar1S28S95N013P019N041P020(0) <='1';
          else
          cVar1S28S95N013P019N041P020(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='0' AND E(15)='0' AND B(17)='1' )then
          cVar1S29S95N013P019N041P020(0) <='1';
          else
          cVar1S29S95N013P019N041P020(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='1' AND D( 0)='0' )then
          cVar1S30S95N013P019P017P066(0) <='1';
          else
          cVar1S30S95N013P019P017P066(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='1' AND D( 0)='0' )then
          cVar1S31S95N013P019P017P066(0) <='1';
          else
          cVar1S31S95N013P019P017P066(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='1' AND D( 0)='0' )then
          cVar1S32S95N013P019P017P066(0) <='1';
          else
          cVar1S32S95N013P019P017P066(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='1' AND D( 0)='0' )then
          cVar1S33S95N013P019P017P066(0) <='1';
          else
          cVar1S33S95N013P019P017P066(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='1' AND D( 0)='1' )then
          cVar1S34S95N013P019P017P066(0) <='1';
          else
          cVar1S34S95N013P019P017P066(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='1' )then
          cVar1S35S95N013P019N017P048(0) <='1';
          else
          cVar1S35S95N013P019N017P048(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='1' )then
          cVar1S36S95N013P019N017P048(0) <='1';
          else
          cVar1S36S95N013P019N017P048(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='1' )then
          cVar1S37S95N013P019N017P048(0) <='1';
          else
          cVar1S37S95N013P019N017P048(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='0' )then
          cVar1S38S95N013P019N017N048(0) <='1';
          else
          cVar1S38S95N013P019N017N048(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='0' )then
          cVar1S39S95N013P019N017N048(0) <='1';
          else
          cVar1S39S95N013P019N017N048(0) <='0';
          end if;
        if(A( 3)='0' AND A( 0)='1' AND A( 1)='0' AND E( 5)='0' )then
          cVar1S40S95N013P019N017N048(0) <='1';
          else
          cVar1S40S95N013P019N017N048(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S0S96P019P012P058P011(0) <='1';
          else
          cVar1S0S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S1S96P019P012P058P011(0) <='1';
          else
          cVar1S1S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S2S96P019P012P058P011(0) <='1';
          else
          cVar1S2S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S3S96P019P012P058P011(0) <='1';
          else
          cVar1S3S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S4S96P019P012P058P011(0) <='1';
          else
          cVar1S4S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S5S96P019P012P058P011(0) <='1';
          else
          cVar1S5S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S6S96P019P012P058P011(0) <='1';
          else
          cVar1S6S96P019P012P058P011(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='0' )then
          cVar1S7S96P019P012P058P068(0) <='1';
          else
          cVar1S7S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='0' )then
          cVar1S8S96P019P012P058P068(0) <='1';
          else
          cVar1S8S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='0' )then
          cVar1S9S96P019P012P058P068(0) <='1';
          else
          cVar1S9S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='0' )then
          cVar1S10S96P019P012P058P068(0) <='1';
          else
          cVar1S10S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='1' )then
          cVar1S11S96P019P012P058P068(0) <='1';
          else
          cVar1S11S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='0' AND D( 2)='1' AND E( 0)='1' )then
          cVar1S12S96P019P012P058P068(0) <='1';
          else
          cVar1S12S96P019P012P058P068(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='1' )then
          cVar1S13S96P019P012P043P056(0) <='1';
          else
          cVar1S13S96P019P012P043P056(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='1' )then
          cVar1S14S96P019P012P043P056(0) <='1';
          else
          cVar1S14S96P019P012P043P056(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='1' )then
          cVar1S15S96P019P012P043P056(0) <='1';
          else
          cVar1S15S96P019P012P043P056(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='0' )then
          cVar1S16S96P019P012P043N056(0) <='1';
          else
          cVar1S16S96P019P012P043N056(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='0' )then
          cVar1S17S96P019P012P043N056(0) <='1';
          else
          cVar1S17S96P019P012P043N056(0) <='0';
          end if;
        if(A( 0)='0' AND A(13)='1' AND D(14)='0' AND E( 3)='0' )then
          cVar1S18S96P019P012P043N056(0) <='1';
          else
          cVar1S18S96P019P012P043N056(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='1' AND A( 2)='0' )then
          cVar1S19S96P019P003P057P015nsss(0) <='1';
          else
          cVar1S19S96P019P003P057P015nsss(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='1' AND A( 2)='1' )then
          cVar1S20S96P019P003P057P015(0) <='1';
          else
          cVar1S20S96P019P003P057P015(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='0' AND E( 0)='1' )then
          cVar1S21S96P019P003N057P068(0) <='1';
          else
          cVar1S21S96P019P003N057P068(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='0' AND E( 0)='1' )then
          cVar1S22S96P019P003N057P068(0) <='1';
          else
          cVar1S22S96P019P003N057P068(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='0' AND E( 0)='0' )then
          cVar1S23S96P019P003N057N068(0) <='1';
          else
          cVar1S23S96P019P003N057N068(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='0' AND E( 0)='0' )then
          cVar1S24S96P019P003N057N068(0) <='1';
          else
          cVar1S24S96P019P003N057N068(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='1' AND E(11)='0' AND E( 0)='0' )then
          cVar1S25S96P019P003N057N068(0) <='1';
          else
          cVar1S25S96P019P003N057N068(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='1' )then
          cVar1S26S96P019N003P057P025(0) <='1';
          else
          cVar1S26S96P019N003P057P025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='1' )then
          cVar1S27S96P019N003P057P025(0) <='1';
          else
          cVar1S27S96P019N003P057P025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='0' )then
          cVar1S28S96P019N003P057N025(0) <='1';
          else
          cVar1S28S96P019N003P057N025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='0' )then
          cVar1S29S96P019N003P057N025(0) <='1';
          else
          cVar1S29S96P019N003P057N025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='0' )then
          cVar1S30S96P019N003P057N025(0) <='1';
          else
          cVar1S30S96P019N003P057N025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='0' AND B( 6)='0' )then
          cVar1S31S96P019N003P057N025(0) <='1';
          else
          cVar1S31S96P019N003P057N025(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='1' AND D( 0)='0' )then
          cVar1S32S96P019N003P057P066(0) <='1';
          else
          cVar1S32S96P019N003P057P066(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='1' AND D( 0)='0' )then
          cVar1S33S96P019N003P057P066(0) <='1';
          else
          cVar1S33S96P019N003P057P066(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='1' AND D( 0)='0' )then
          cVar1S34S96P019N003P057P066(0) <='1';
          else
          cVar1S34S96P019N003P057P066(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='1' AND D( 0)='1' )then
          cVar1S35S96P019N003P057P066(0) <='1';
          else
          cVar1S35S96P019N003P057P066(0) <='0';
          end if;
        if(A( 0)='1' AND A( 8)='0' AND E(11)='1' AND D( 0)='1' )then
          cVar1S36S96P019N003P057P066(0) <='1';
          else
          cVar1S36S96P019N003P057P066(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='1' AND A( 6)='1' )then
          cVar1S0S97P019P057P069P007(0) <='1';
          else
          cVar1S0S97P019P057P069P007(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='1' AND A( 6)='1' )then
          cVar1S1S97P019P057P069P007(0) <='1';
          else
          cVar1S1S97P019P057P069P007(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='1' AND A( 6)='0' )then
          cVar1S2S97P019P057P069N007(0) <='1';
          else
          cVar1S2S97P019P057P069N007(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='1' AND A( 6)='0' )then
          cVar1S3S97P019P057P069N007(0) <='1';
          else
          cVar1S3S97P019P057P069N007(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='1' AND A( 6)='0' )then
          cVar1S4S97P019P057P069N007(0) <='1';
          else
          cVar1S4S97P019P057P069N007(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='0' AND D( 7)='0' )then
          cVar1S5S97P019P057N069P038(0) <='1';
          else
          cVar1S5S97P019P057N069P038(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='0' AND D( 7)='0' )then
          cVar1S6S97P019P057N069P038(0) <='1';
          else
          cVar1S6S97P019P057N069P038(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='0' AND D( 7)='0' )then
          cVar1S7S97P019P057N069P038(0) <='1';
          else
          cVar1S7S97P019P057N069P038(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='0' AND E( 8)='0' AND D( 7)='1' )then
          cVar1S8S97P019P057N069P038(0) <='1';
          else
          cVar1S8S97P019P057N069P038(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='1' AND A( 2)='0' )then
          cVar1S9S97P019P057P003P015nsss(0) <='1';
          else
          cVar1S9S97P019P057P003P015nsss(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='1' AND A( 2)='1' )then
          cVar1S10S97P019P057P003P015(0) <='1';
          else
          cVar1S10S97P019P057P003P015(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='0' AND A( 4)='1' )then
          cVar1S11S97P019P057N003P011(0) <='1';
          else
          cVar1S11S97P019P057N003P011(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='0' AND A( 4)='1' )then
          cVar1S12S97P019P057N003P011(0) <='1';
          else
          cVar1S12S97P019P057N003P011(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='0' AND A( 4)='0' )then
          cVar1S13S97P019P057N003N011(0) <='1';
          else
          cVar1S13S97P019P057N003N011(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='0' AND A( 4)='0' )then
          cVar1S14S97P019P057N003N011(0) <='1';
          else
          cVar1S14S97P019P057N003N011(0) <='0';
          end if;
        if(A( 0)='1' AND E(11)='1' AND A( 8)='0' AND A( 4)='0' )then
          cVar1S15S97P019P057N003N011(0) <='1';
          else
          cVar1S15S97P019P057N003N011(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND D(11)='0' )then
          cVar1S16S97N019P060P021P055(0) <='1';
          else
          cVar1S16S97N019P060P021P055(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND D(11)='0' )then
          cVar1S17S97N019P060P021P055(0) <='1';
          else
          cVar1S17S97N019P060P021P055(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND D(11)='0' )then
          cVar1S18S97N019P060P021P055(0) <='1';
          else
          cVar1S18S97N019P060P021P055(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND D(11)='1' )then
          cVar1S19S97N019P060P021P055(0) <='1';
          else
          cVar1S19S97N019P060P021P055(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND D(11)='1' )then
          cVar1S20S97N019P060P021P055(0) <='1';
          else
          cVar1S20S97N019P060P021P055(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='1' AND B( 2)='1' )then
          cVar1S21S97N019P060P021P033nsss(0) <='1';
          else
          cVar1S21S97N019P060P021P033nsss(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='0' AND B( 9)='1' )then
          cVar1S22S97N019N060P068P036(0) <='1';
          else
          cVar1S22S97N019N060P068P036(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='0' AND B( 9)='1' )then
          cVar1S23S97N019N060P068P036(0) <='1';
          else
          cVar1S23S97N019N060P068P036(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='0' AND B( 9)='0' )then
          cVar1S24S97N019N060P068N036(0) <='1';
          else
          cVar1S24S97N019N060P068N036(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='0' AND B( 9)='0' )then
          cVar1S25S97N019N060P068N036(0) <='1';
          else
          cVar1S25S97N019N060P068N036(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='0' AND B( 9)='0' )then
          cVar1S26S97N019N060P068N036(0) <='1';
          else
          cVar1S26S97N019N060P068N036(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='1' AND B( 7)='0' )then
          cVar1S27S97N019N060P068P023(0) <='1';
          else
          cVar1S27S97N019N060P068P023(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='1' AND B( 7)='0' )then
          cVar1S28S97N019N060P068P023(0) <='1';
          else
          cVar1S28S97N019N060P068P023(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='1' AND B( 7)='0' )then
          cVar1S29S97N019N060P068P023(0) <='1';
          else
          cVar1S29S97N019N060P068P023(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='1' AND B( 7)='0' )then
          cVar1S30S97N019N060P068P023(0) <='1';
          else
          cVar1S30S97N019N060P068P023(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND E( 0)='1' AND B( 7)='1' )then
          cVar1S31S97N019N060P068P023(0) <='1';
          else
          cVar1S31S97N019N060P068P023(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S0S98P019P060P033P003(0) <='1';
          else
          cVar1S0S98P019P060P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S1S98P019P060P033P003(0) <='1';
          else
          cVar1S1S98P019P060P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S2S98P019P060P033P003(0) <='1';
          else
          cVar1S2S98P019P060P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='1' AND A( 8)='0' )then
          cVar1S3S98P019P060P033P003(0) <='1';
          else
          cVar1S3S98P019P060P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='1' AND A( 8)='1' )then
          cVar1S4S98P019P060P033P003(0) <='1';
          else
          cVar1S4S98P019P060P033P003(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='0' AND D( 2)='0' )then
          cVar1S5S98P019P060N033P058(0) <='1';
          else
          cVar1S5S98P019P060N033P058(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='0' AND D( 2)='0' )then
          cVar1S6S98P019P060N033P058(0) <='1';
          else
          cVar1S6S98P019P060N033P058(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='0' AND D( 2)='1' )then
          cVar1S7S98P019P060N033P058(0) <='1';
          else
          cVar1S7S98P019P060N033P058(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='0' AND B( 2)='0' AND D( 2)='1' )then
          cVar1S8S98P019P060N033P058(0) <='1';
          else
          cVar1S8S98P019P060N033P058(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND A(14)='1' )then
          cVar1S9S98P019P060P021P010(0) <='1';
          else
          cVar1S9S98P019P060P021P010(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND A(14)='1' )then
          cVar1S10S98P019P060P021P010(0) <='1';
          else
          cVar1S10S98P019P060P021P010(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND A(14)='1' )then
          cVar1S11S98P019P060P021P010(0) <='1';
          else
          cVar1S11S98P019P060P021P010(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S12S98P019P060P021N010(0) <='1';
          else
          cVar1S12S98P019P060P021N010(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='0' AND A(14)='0' )then
          cVar1S13S98P019P060P021N010(0) <='1';
          else
          cVar1S13S98P019P060P021N010(0) <='0';
          end if;
        if(A( 0)='0' AND E( 2)='1' AND B( 8)='1' AND B( 2)='1' )then
          cVar1S14S98P019P060P021P033nsss(0) <='1';
          else
          cVar1S14S98P019P060P021P033nsss(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='1' AND A( 1)='0' )then
          cVar1S15S98P019P069P013P017(0) <='1';
          else
          cVar1S15S98P019P069P013P017(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='1' AND A( 1)='0' )then
          cVar1S16S98P019P069P013P017(0) <='1';
          else
          cVar1S16S98P019P069P013P017(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='1' AND A( 1)='1' )then
          cVar1S17S98P019P069P013P017(0) <='1';
          else
          cVar1S17S98P019P069P013P017(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='1' AND A( 1)='1' )then
          cVar1S18S98P019P069P013P017(0) <='1';
          else
          cVar1S18S98P019P069P013P017(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='0' AND B(16)='1' )then
          cVar1S19S98P019P069N013P022nsss(0) <='1';
          else
          cVar1S19S98P019P069N013P022nsss(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='0' AND B(16)='0' )then
          cVar1S20S98P019P069N013N022(0) <='1';
          else
          cVar1S20S98P019P069N013N022(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='0' AND B(16)='0' )then
          cVar1S21S98P019P069N013N022(0) <='1';
          else
          cVar1S21S98P019P069N013N022(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A( 3)='0' AND B(16)='0' )then
          cVar1S22S98P019P069N013N022(0) <='1';
          else
          cVar1S22S98P019P069N013N022(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='1' AND D( 9)='1' )then
          cVar1S23S98P019N069P058P063(0) <='1';
          else
          cVar1S23S98P019N069P058P063(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='1' AND D( 9)='1' )then
          cVar1S24S98P019N069P058P063(0) <='1';
          else
          cVar1S24S98P019N069P058P063(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='1' AND D( 9)='0' )then
          cVar1S25S98P019N069P058N063(0) <='1';
          else
          cVar1S25S98P019N069P058N063(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='1' AND D( 9)='0' )then
          cVar1S26S98P019N069P058N063(0) <='1';
          else
          cVar1S26S98P019N069P058N063(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='0' AND E( 2)='0' )then
          cVar1S27S98P019N069N058P060(0) <='1';
          else
          cVar1S27S98P019N069N058P060(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='0' AND E( 2)='0' )then
          cVar1S28S98P019N069N058P060(0) <='1';
          else
          cVar1S28S98P019N069N058P060(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='0' AND E( 2)='0' )then
          cVar1S29S98P019N069N058P060(0) <='1';
          else
          cVar1S29S98P019N069N058P060(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND D( 2)='0' AND E( 2)='1' )then
          cVar1S30S98P019N069N058P060(0) <='1';
          else
          cVar1S30S98P019N069N058P060(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='1' AND B( 5)='1' )then
          cVar1S0S99P019P069P006P027nsss(0) <='1';
          else
          cVar1S0S99P019P069P006P027nsss(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='1' AND B( 5)='0' )then
          cVar1S1S99P019P069P006N027(0) <='1';
          else
          cVar1S1S99P019P069P006N027(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='1' AND B( 5)='0' )then
          cVar1S2S99P019P069P006N027(0) <='1';
          else
          cVar1S2S99P019P069P006N027(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='1' AND B( 5)='0' )then
          cVar1S3S99P019P069P006N027(0) <='1';
          else
          cVar1S3S99P019P069P006N027(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='0' AND D(13)='0' )then
          cVar1S4S99P019P069N006P047(0) <='1';
          else
          cVar1S4S99P019P069N006P047(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='0' AND D(13)='0' )then
          cVar1S5S99P019P069N006P047(0) <='1';
          else
          cVar1S5S99P019P069N006P047(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='0' AND D(13)='0' )then
          cVar1S6S99P019P069N006P047(0) <='1';
          else
          cVar1S6S99P019P069N006P047(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='1' AND A(16)='0' AND D(13)='1' )then
          cVar1S7S99P019P069N006P047(0) <='1';
          else
          cVar1S7S99P019P069N006P047(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='1' )then
          cVar1S8S99P019N069P060P016(0) <='1';
          else
          cVar1S8S99P019N069P060P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='1' )then
          cVar1S9S99P019N069P060P016(0) <='1';
          else
          cVar1S9S99P019N069P060P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='1' )then
          cVar1S10S99P019N069P060P016(0) <='1';
          else
          cVar1S10S99P019N069P060P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='1' )then
          cVar1S11S99P019N069P060P016(0) <='1';
          else
          cVar1S11S99P019N069P060P016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='0' )then
          cVar1S12S99P019N069P060N016(0) <='1';
          else
          cVar1S12S99P019N069P060N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='0' )then
          cVar1S13S99P019N069P060N016(0) <='1';
          else
          cVar1S13S99P019N069P060N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='0' )then
          cVar1S14S99P019N069P060N016(0) <='1';
          else
          cVar1S14S99P019N069P060N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='0' AND A(11)='0' )then
          cVar1S15S99P019N069P060N016(0) <='1';
          else
          cVar1S15S99P019N069P060N016(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='1' AND D( 2)='1' )then
          cVar1S16S99P019N069P060P058(0) <='1';
          else
          cVar1S16S99P019N069P060P058(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='1' AND D( 2)='0' )then
          cVar1S17S99P019N069P060N058(0) <='1';
          else
          cVar1S17S99P019N069P060N058(0) <='0';
          end if;
        if(A( 0)='1' AND E( 8)='0' AND E( 2)='1' AND D( 2)='0' )then
          cVar1S18S99P019N069P060N058(0) <='1';
          else
          cVar1S18S99P019N069P060N058(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='0' AND A( 8)='0' )then
          cVar1S19S99N019P033P030P003(0) <='1';
          else
          cVar1S19S99N019P033P030P003(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='0' AND A( 8)='0' )then
          cVar1S20S99N019P033P030P003(0) <='1';
          else
          cVar1S20S99N019P033P030P003(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='0' AND A( 8)='0' )then
          cVar1S21S99N019P033P030P003(0) <='1';
          else
          cVar1S21S99N019P033P030P003(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='0' AND A( 8)='1' )then
          cVar1S22S99N019P033P030P003(0) <='1';
          else
          cVar1S22S99N019P033P030P003(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='1' AND A(13)='0' )then
          cVar1S23S99N019P033P030P012(0) <='1';
          else
          cVar1S23S99N019P033P030P012(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='1' AND A(13)='0' )then
          cVar1S24S99N019P033P030P012(0) <='1';
          else
          cVar1S24S99N019P033P030P012(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='1' AND A(13)='0' )then
          cVar1S25S99N019P033P030P012(0) <='1';
          else
          cVar1S25S99N019P033P030P012(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='1' AND B(12)='1' AND A(13)='1' )then
          cVar1S26S99N019P033P030P012(0) <='1';
          else
          cVar1S26S99N019P033P030P012(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='1' )then
          cVar1S27S99N019N033P036P027(0) <='1';
          else
          cVar1S27S99N019N033P036P027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='1' )then
          cVar1S28S99N019N033P036P027(0) <='1';
          else
          cVar1S28S99N019N033P036P027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='1' )then
          cVar1S29S99N019N033P036P027(0) <='1';
          else
          cVar1S29S99N019N033P036P027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='0' )then
          cVar1S30S99N019N033P036N027(0) <='1';
          else
          cVar1S30S99N019N033P036N027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='0' )then
          cVar1S31S99N019N033P036N027(0) <='1';
          else
          cVar1S31S99N019N033P036N027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='0' AND B( 5)='0' )then
          cVar1S32S99N019N033P036N027(0) <='1';
          else
          cVar1S32S99N019N033P036N027(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='1' AND B( 8)='0' )then
          cVar1S33S99N019N033P036P021(0) <='1';
          else
          cVar1S33S99N019N033P036P021(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='1' AND B( 8)='0' )then
          cVar1S34S99N019N033P036P021(0) <='1';
          else
          cVar1S34S99N019N033P036P021(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='1' AND B( 8)='1' )then
          cVar1S35S99N019N033P036P021(0) <='1';
          else
          cVar1S35S99N019N033P036P021(0) <='0';
          end if;
        if(A( 0)='0' AND B( 2)='0' AND B( 9)='1' AND B( 8)='1' )then
          cVar1S36S99N019N033P036P021(0) <='1';
          else
          cVar1S36S99N019N033P036P021(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='1' )then
          cVar1S0S100P036P012P019P014(0) <='1';
          else
          cVar1S0S100P036P012P019P014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='1' )then
          cVar1S1S100P036P012P019P014(0) <='1';
          else
          cVar1S1S100P036P012P019P014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='1' )then
          cVar1S2S100P036P012P019P014(0) <='1';
          else
          cVar1S2S100P036P012P019P014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='0' )then
          cVar1S3S100P036P012P019N014(0) <='1';
          else
          cVar1S3S100P036P012P019N014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='0' )then
          cVar1S4S100P036P012P019N014(0) <='1';
          else
          cVar1S4S100P036P012P019N014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='0' )then
          cVar1S5S100P036P012P019N014(0) <='1';
          else
          cVar1S5S100P036P012P019N014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='0' AND A(12)='0' )then
          cVar1S6S100P036P012P019N014(0) <='1';
          else
          cVar1S6S100P036P012P019N014(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='1' )then
          cVar1S7S100P036P012P019P016(0) <='1';
          else
          cVar1S7S100P036P012P019P016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='1' )then
          cVar1S8S100P036P012P019P016(0) <='1';
          else
          cVar1S8S100P036P012P019P016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='1' )then
          cVar1S9S100P036P012P019P016(0) <='1';
          else
          cVar1S9S100P036P012P019P016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='1' )then
          cVar1S10S100P036P012P019P016(0) <='1';
          else
          cVar1S10S100P036P012P019P016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='0' )then
          cVar1S11S100P036P012P019N016(0) <='1';
          else
          cVar1S11S100P036P012P019N016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='0' )then
          cVar1S12S100P036P012P019N016(0) <='1';
          else
          cVar1S12S100P036P012P019N016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='0' AND A( 0)='1' AND A(11)='0' )then
          cVar1S13S100P036P012P019N016(0) <='1';
          else
          cVar1S13S100P036P012P019N016(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='1' )then
          cVar1S14S100P036P012P018P066(0) <='1';
          else
          cVar1S14S100P036P012P018P066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='1' )then
          cVar1S15S100P036P012P018P066(0) <='1';
          else
          cVar1S15S100P036P012P018P066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='1' )then
          cVar1S16S100P036P012P018P066(0) <='1';
          else
          cVar1S16S100P036P012P018P066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='1' )then
          cVar1S17S100P036P012P018P066(0) <='1';
          else
          cVar1S17S100P036P012P018P066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='0' )then
          cVar1S18S100P036P012P018N066(0) <='1';
          else
          cVar1S18S100P036P012P018N066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='0' )then
          cVar1S19S100P036P012P018N066(0) <='1';
          else
          cVar1S19S100P036P012P018N066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='1' AND D( 0)='0' )then
          cVar1S20S100P036P012P018N066(0) <='1';
          else
          cVar1S20S100P036P012P018N066(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='0' AND D(14)='0' )then
          cVar1S21S100P036P012N018P043(0) <='1';
          else
          cVar1S21S100P036P012N018P043(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='0' AND D(14)='0' )then
          cVar1S22S100P036P012N018P043(0) <='1';
          else
          cVar1S22S100P036P012N018P043(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='0' AND D(14)='0' )then
          cVar1S23S100P036P012N018P043(0) <='1';
          else
          cVar1S23S100P036P012N018P043(0) <='0';
          end if;
        if(B( 9)='0' AND A(13)='1' AND A(10)='0' AND D(14)='1' )then
          cVar1S24S100P036P012N018P043(0) <='1';
          else
          cVar1S24S100P036P012N018P043(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S25S100P036P006P053P033(0) <='1';
          else
          cVar1S25S100P036P006P053P033(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S26S100P036P006P053P033(0) <='1';
          else
          cVar1S26S100P036P006P053P033(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S27S100P036P006P053P033(0) <='1';
          else
          cVar1S27S100P036P006P053P033(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='1' AND E(12)='0' AND B( 2)='1' )then
          cVar1S28S100P036P006P053P033(0) <='1';
          else
          cVar1S28S100P036P006P053P033(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='1' AND B(14)='1' )then
          cVar1S29S100P036N006P008P026(0) <='1';
          else
          cVar1S29S100P036N006P008P026(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='1' AND B(14)='0' )then
          cVar1S30S100P036N006P008N026(0) <='1';
          else
          cVar1S30S100P036N006P008N026(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='1' AND B(14)='0' )then
          cVar1S31S100P036N006P008N026(0) <='1';
          else
          cVar1S31S100P036N006P008N026(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='1' AND B(14)='0' )then
          cVar1S32S100P036N006P008N026(0) <='1';
          else
          cVar1S32S100P036N006P008N026(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='0' AND D(13)='0' )then
          cVar1S33S100P036N006N008P047(0) <='1';
          else
          cVar1S33S100P036N006N008P047(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='0' AND D(13)='0' )then
          cVar1S34S100P036N006N008P047(0) <='1';
          else
          cVar1S34S100P036N006N008P047(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='0' AND D(13)='0' )then
          cVar1S35S100P036N006N008P047(0) <='1';
          else
          cVar1S35S100P036N006N008P047(0) <='0';
          end if;
        if(B( 9)='1' AND A(16)='0' AND A(15)='0' AND D(13)='1' )then
          cVar1S36S100P036N006N008P047(0) <='1';
          else
          cVar1S36S100P036N006N008P047(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S0S101P036P005P023P029(0) <='1';
          else
          cVar1S0S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S1S101P036P005P023P029(0) <='1';
          else
          cVar1S1S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S2S101P036P005P023P029(0) <='1';
          else
          cVar1S2S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S3S101P036P005P023P029(0) <='1';
          else
          cVar1S3S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='1' )then
          cVar1S4S101P036P005P023P029(0) <='1';
          else
          cVar1S4S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='0' AND B( 4)='1' )then
          cVar1S5S101P036P005P023P029(0) <='1';
          else
          cVar1S5S101P036P005P023P029(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='1' AND A(17)='1' )then
          cVar1S6S101P036P005P023P004nsss(0) <='1';
          else
          cVar1S6S101P036P005P023P004nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND B( 7)='1' AND A(17)='0' )then
          cVar1S7S101P036P005P023N004(0) <='1';
          else
          cVar1S7S101P036P005P023N004(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND E( 8)='1' AND A( 3)='0' )then
          cVar1S8S101P036P005P069P013(0) <='1';
          else
          cVar1S8S101P036P005P069P013(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND E( 8)='1' AND A( 3)='0' )then
          cVar1S9S101P036P005P069P013(0) <='1';
          else
          cVar1S9S101P036P005P069P013(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND E( 8)='0' AND B(11)='1' )then
          cVar1S10S101P036P005N069P032nsss(0) <='1';
          else
          cVar1S10S101P036P005N069P032nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND E( 8)='0' AND B(11)='0' )then
          cVar1S11S101P036P005N069N032(0) <='1';
          else
          cVar1S11S101P036P005N069N032(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='1' )then
          cVar1S12S101N036P014P061P069(0) <='1';
          else
          cVar1S12S101N036P014P061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='1' )then
          cVar1S13S101N036P014P061P069(0) <='1';
          else
          cVar1S13S101N036P014P061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='1' )then
          cVar1S14S101N036P014P061P069(0) <='1';
          else
          cVar1S14S101N036P014P061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S15S101N036P014P061N069(0) <='1';
          else
          cVar1S15S101N036P014P061N069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S16S101N036P014P061N069(0) <='1';
          else
          cVar1S16S101N036P014P061N069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='1' AND E( 8)='0' )then
          cVar1S17S101N036P014P061N069(0) <='1';
          else
          cVar1S17S101N036P014P061N069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='0' AND E( 8)='0' )then
          cVar1S18S101N036P014N061P069(0) <='1';
          else
          cVar1S18S101N036P014N061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='0' AND E( 8)='0' )then
          cVar1S19S101N036P014N061P069(0) <='1';
          else
          cVar1S19S101N036P014N061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='0' AND E( 8)='0' )then
          cVar1S20S101N036P014N061P069(0) <='1';
          else
          cVar1S20S101N036P014N061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='0' AND E( 8)='1' )then
          cVar1S21S101N036P014N061P069(0) <='1';
          else
          cVar1S21S101N036P014N061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='1' AND E(10)='0' AND E( 8)='1' )then
          cVar1S22S101N036P014N061P069(0) <='1';
          else
          cVar1S22S101N036P014N061P069(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='1' AND B( 7)='0' )then
          cVar1S23S101N036N014P012P023(0) <='1';
          else
          cVar1S23S101N036N014P012P023(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='1' AND B( 7)='0' )then
          cVar1S24S101N036N014P012P023(0) <='1';
          else
          cVar1S24S101N036N014P012P023(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='1' AND B( 7)='0' )then
          cVar1S25S101N036N014P012P023(0) <='1';
          else
          cVar1S25S101N036N014P012P023(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='1' AND B( 7)='0' )then
          cVar1S26S101N036N014P012P023(0) <='1';
          else
          cVar1S26S101N036N014P012P023(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='1' AND B( 7)='1' )then
          cVar1S27S101N036N014P012P023(0) <='1';
          else
          cVar1S27S101N036N014P012P023(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='0' AND A( 2)='0' )then
          cVar1S28S101N036N014N012P015(0) <='1';
          else
          cVar1S28S101N036N014N012P015(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='0' AND A( 2)='0' )then
          cVar1S29S101N036N014N012P015(0) <='1';
          else
          cVar1S29S101N036N014N012P015(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='0' AND A( 2)='0' )then
          cVar1S30S101N036N014N012P015(0) <='1';
          else
          cVar1S30S101N036N014N012P015(0) <='0';
          end if;
        if(B( 9)='0' AND A(12)='0' AND A(13)='0' AND A( 2)='1' )then
          cVar1S31S101N036N014N012P015(0) <='1';
          else
          cVar1S31S101N036N014N012P015(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='1' AND B( 3)='0' )then
          cVar1S0S102P036P016P030P031(0) <='1';
          else
          cVar1S0S102P036P016P030P031(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='1' AND B( 3)='0' )then
          cVar1S1S102P036P016P030P031(0) <='1';
          else
          cVar1S1S102P036P016P030P031(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='1' AND B( 3)='0' )then
          cVar1S2S102P036P016P030P031(0) <='1';
          else
          cVar1S2S102P036P016P030P031(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='1' AND B( 3)='1' )then
          cVar1S3S102P036P016P030P031(0) <='1';
          else
          cVar1S3S102P036P016P030P031(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='1' )then
          cVar1S4S102P036P016N030P028(0) <='1';
          else
          cVar1S4S102P036P016N030P028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='1' )then
          cVar1S5S102P036P016N030P028(0) <='1';
          else
          cVar1S5S102P036P016N030P028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='1' )then
          cVar1S6S102P036P016N030P028(0) <='1';
          else
          cVar1S6S102P036P016N030P028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='1' )then
          cVar1S7S102P036P016N030P028(0) <='1';
          else
          cVar1S7S102P036P016N030P028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='0' )then
          cVar1S8S102P036P016N030N028(0) <='1';
          else
          cVar1S8S102P036P016N030N028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='0' )then
          cVar1S9S102P036P016N030N028(0) <='1';
          else
          cVar1S9S102P036P016N030N028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='0' AND B(12)='0' AND B(13)='0' )then
          cVar1S10S102P036P016N030N028(0) <='1';
          else
          cVar1S10S102P036P016N030N028(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='1' AND D(15)='0' )then
          cVar1S11S102P036P016P014P039(0) <='1';
          else
          cVar1S11S102P036P016P014P039(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='1' AND D(15)='0' )then
          cVar1S12S102P036P016P014P039(0) <='1';
          else
          cVar1S12S102P036P016P014P039(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='1' AND D(15)='0' )then
          cVar1S13S102P036P016P014P039(0) <='1';
          else
          cVar1S13S102P036P016P014P039(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='1' AND D(15)='0' )then
          cVar1S14S102P036P016P014P039(0) <='1';
          else
          cVar1S14S102P036P016P014P039(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='1' )then
          cVar1S15S102P036P016N014P037(0) <='1';
          else
          cVar1S15S102P036P016N014P037(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='1' )then
          cVar1S16S102P036P016N014P037(0) <='1';
          else
          cVar1S16S102P036P016N014P037(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='1' )then
          cVar1S17S102P036P016N014P037(0) <='1';
          else
          cVar1S17S102P036P016N014P037(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='0' )then
          cVar1S18S102P036P016N014N037(0) <='1';
          else
          cVar1S18S102P036P016N014N037(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='0' )then
          cVar1S19S102P036P016N014N037(0) <='1';
          else
          cVar1S19S102P036P016N014N037(0) <='0';
          end if;
        if(B( 9)='0' AND A(11)='1' AND A(12)='0' AND B( 0)='0' )then
          cVar1S20S102P036P016N014N037(0) <='1';
          else
          cVar1S20S102P036P016N014N037(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='1' AND E( 8)='1' AND A( 5)='0' )then
          cVar1S21S102P036P000P069P009nsss(0) <='1';
          else
          cVar1S21S102P036P000P069P009nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='1' AND E( 8)='0' AND A( 3)='0' )then
          cVar1S22S102P036P000N069P013(0) <='1';
          else
          cVar1S22S102P036P000N069P013(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='1' AND E( 8)='0' AND A( 3)='0' )then
          cVar1S23S102P036P000N069P013(0) <='1';
          else
          cVar1S23S102P036P000N069P013(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='1' AND B( 0)='0' )then
          cVar1S24S102P036N000P030P037(0) <='1';
          else
          cVar1S24S102P036N000P030P037(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='1' AND B( 0)='1' )then
          cVar1S25S102P036N000P030P037(0) <='1';
          else
          cVar1S25S102P036N000P030P037(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='1' AND B( 0)='1' )then
          cVar1S26S102P036N000P030P037(0) <='1';
          else
          cVar1S26S102P036N000P030P037(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S27S102P036N000N030P057(0) <='1';
          else
          cVar1S27S102P036N000N030P057(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S28S102P036N000N030P057(0) <='1';
          else
          cVar1S28S102P036N000N030P057(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S29S102P036N000N030P057(0) <='1';
          else
          cVar1S29S102P036N000N030P057(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='0' AND E(11)='1' )then
          cVar1S30S102P036N000N030P057(0) <='1';
          else
          cVar1S30S102P036N000N030P057(0) <='0';
          end if;
        if(B( 9)='1' AND A(19)='0' AND B(12)='0' AND E(11)='1' )then
          cVar1S31S102P036N000N030P057(0) <='1';
          else
          cVar1S31S102P036N000N030P057(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='0' AND D(14)='1' )then
          cVar1S0S103P036P001P023P043(0) <='1';
          else
          cVar1S0S103P036P001P023P043(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='0' AND D(14)='1' )then
          cVar1S1S103P036P001P023P043(0) <='1';
          else
          cVar1S1S103P036P001P023P043(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='0' AND D(14)='0' )then
          cVar1S2S103P036P001P023N043(0) <='1';
          else
          cVar1S2S103P036P001P023N043(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='0' AND D(14)='0' )then
          cVar1S3S103P036P001P023N043(0) <='1';
          else
          cVar1S3S103P036P001P023N043(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='0' AND D(14)='0' )then
          cVar1S4S103P036P001P023N043(0) <='1';
          else
          cVar1S4S103P036P001P023N043(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='0' AND B( 7)='1' AND D( 6)='1' )then
          cVar1S5S103P036P001P023P042(0) <='1';
          else
          cVar1S5S103P036P001P023P042(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='1' AND B(10)='1' AND B( 0)='0' )then
          cVar1S6S103P036P001P034P037nsss(0) <='1';
          else
          cVar1S6S103P036P001P034P037nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='1' AND B(10)='0' AND B( 2)='1' )then
          cVar1S7S103P036P001N034P033nsss(0) <='1';
          else
          cVar1S7S103P036P001N034P033nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A( 9)='1' AND B(10)='0' AND B( 2)='0' )then
          cVar1S8S103P036P001N034N033(0) <='1';
          else
          cVar1S8S103P036P001N034N033(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='0' )then
          cVar1S9S103N036P011P040P010(0) <='1';
          else
          cVar1S9S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='0' )then
          cVar1S10S103N036P011P040P010(0) <='1';
          else
          cVar1S10S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='0' )then
          cVar1S11S103N036P011P040P010(0) <='1';
          else
          cVar1S11S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='0' )then
          cVar1S12S103N036P011P040P010(0) <='1';
          else
          cVar1S12S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='1' )then
          cVar1S13S103N036P011P040P010(0) <='1';
          else
          cVar1S13S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='0' AND A(14)='1' )then
          cVar1S14S103N036P011P040P010(0) <='1';
          else
          cVar1S14S103N036P011P040P010(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='1' AND D( 7)='1' )then
          cVar1S15S103N036P011P040P038nsss(0) <='1';
          else
          cVar1S15S103N036P011P040P038nsss(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='1' AND E( 7)='1' AND D( 7)='0' )then
          cVar1S16S103N036P011P040N038(0) <='1';
          else
          cVar1S16S103N036P011P040N038(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='0' )then
          cVar1S17S103N036N011P016P055(0) <='1';
          else
          cVar1S17S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='0' )then
          cVar1S18S103N036N011P016P055(0) <='1';
          else
          cVar1S18S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='0' )then
          cVar1S19S103N036N011P016P055(0) <='1';
          else
          cVar1S19S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='0' )then
          cVar1S20S103N036N011P016P055(0) <='1';
          else
          cVar1S20S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='1' )then
          cVar1S21S103N036N011P016P055(0) <='1';
          else
          cVar1S21S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='1' AND D(11)='1' )then
          cVar1S22S103N036N011P016P055(0) <='1';
          else
          cVar1S22S103N036N011P016P055(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='1' )then
          cVar1S23S103N036N011N016P013(0) <='1';
          else
          cVar1S23S103N036N011N016P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='1' )then
          cVar1S24S103N036N011N016P013(0) <='1';
          else
          cVar1S24S103N036N011N016P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='1' )then
          cVar1S25S103N036N011N016P013(0) <='1';
          else
          cVar1S25S103N036N011N016P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='1' )then
          cVar1S26S103N036N011N016P013(0) <='1';
          else
          cVar1S26S103N036N011N016P013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='0' )then
          cVar1S27S103N036N011N016N013(0) <='1';
          else
          cVar1S27S103N036N011N016N013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='0' )then
          cVar1S28S103N036N011N016N013(0) <='1';
          else
          cVar1S28S103N036N011N016N013(0) <='0';
          end if;
        if(B( 9)='0' AND A( 4)='0' AND A(11)='0' AND A( 3)='0' )then
          cVar1S29S103N036N011N016N013(0) <='1';
          else
          cVar1S29S103N036N011N016N013(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='1' AND E( 5)='0' )then
          cVar1S0S104P036P051P026P048(0) <='1';
          else
          cVar1S0S104P036P051P026P048(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='1' AND E( 5)='0' )then
          cVar1S1S104P036P051P026P048(0) <='1';
          else
          cVar1S1S104P036P051P026P048(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='0' AND B(13)='1' )then
          cVar1S2S104P036P051N026P028(0) <='1';
          else
          cVar1S2S104P036P051N026P028(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='0' AND B(13)='1' )then
          cVar1S3S104P036P051N026P028(0) <='1';
          else
          cVar1S3S104P036P051N026P028(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='0' AND B(13)='1' )then
          cVar1S4S104P036P051N026P028(0) <='1';
          else
          cVar1S4S104P036P051N026P028(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='1' AND B(14)='0' AND B(13)='0' )then
          cVar1S5S104P036P051N026N028(0) <='1';
          else
          cVar1S5S104P036P051N026N028(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='0' )then
          cVar1S6S104P036N051P053P009(0) <='1';
          else
          cVar1S6S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='0' )then
          cVar1S7S104P036N051P053P009(0) <='1';
          else
          cVar1S7S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='0' )then
          cVar1S8S104P036N051P053P009(0) <='1';
          else
          cVar1S8S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='0' )then
          cVar1S9S104P036N051P053P009(0) <='1';
          else
          cVar1S9S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='1' )then
          cVar1S10S104P036N051P053P009(0) <='1';
          else
          cVar1S10S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='0' AND A( 5)='1' )then
          cVar1S11S104P036N051P053P009(0) <='1';
          else
          cVar1S11S104P036N051P053P009(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='1' AND B(14)='0' )then
          cVar1S12S104P036N051P053P026(0) <='1';
          else
          cVar1S12S104P036N051P053P026(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='1' AND B(14)='0' )then
          cVar1S13S104P036N051P053P026(0) <='1';
          else
          cVar1S13S104P036N051P053P026(0) <='0';
          end if;
        if(B( 9)='0' AND D(12)='0' AND E(12)='1' AND B(14)='0' )then
          cVar1S14S104P036N051P053P026(0) <='1';
          else
          cVar1S14S104P036N051P053P026(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='1' )then
          cVar1S15S104P036P043P022nsss(0) <='1';
          else
          cVar1S15S104P036P043P022nsss(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND B(15)='1' )then
          cVar1S16S104P036P043N022P024nsss(0) <='1';
          else
          cVar1S16S104P036P043N022P024nsss(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND B(15)='0' )then
          cVar1S17S104P036P043N022N024(0) <='1';
          else
          cVar1S17S104P036P043N022N024(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='1' AND B(16)='0' AND B(15)='0' )then
          cVar1S18S104P036P043N022N024(0) <='1';
          else
          cVar1S18S104P036P043N022N024(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND D( 7)='0' )then
          cVar1S19S104P036N043P045P038(0) <='1';
          else
          cVar1S19S104P036N043P045P038(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND D( 7)='0' )then
          cVar1S20S104P036N043P045P038(0) <='1';
          else
          cVar1S20S104P036N043P045P038(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='0' AND D( 7)='1' )then
          cVar1S21S104P036N043P045P038(0) <='1';
          else
          cVar1S21S104P036N043P045P038(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='1' AND A(11)='1' )then
          cVar1S22S104P036N043P045P016(0) <='1';
          else
          cVar1S22S104P036N043P045P016(0) <='0';
          end if;
        if(B( 9)='1' AND D(14)='0' AND E(14)='1' AND A(11)='0' )then
          cVar1S23S104P036N043P045N016(0) <='1';
          else
          cVar1S23S104P036N043P045N016(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='0' AND B(12)='1' )then
          cVar1S0S105P013P061P016P030(0) <='1';
          else
          cVar1S0S105P013P061P016P030(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='0' AND B(12)='0' )then
          cVar1S1S105P013P061P016N030(0) <='1';
          else
          cVar1S1S105P013P061P016N030(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='0' AND B(12)='0' )then
          cVar1S2S105P013P061P016N030(0) <='1';
          else
          cVar1S2S105P013P061P016N030(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='1' AND B( 2)='1' )then
          cVar1S3S105P013P061P016P033(0) <='1';
          else
          cVar1S3S105P013P061P016P033(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='1' AND B( 2)='0' )then
          cVar1S4S105P013P061P016N033(0) <='1';
          else
          cVar1S4S105P013P061P016N033(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='1' AND B( 2)='0' )then
          cVar1S5S105P013P061P016N033(0) <='1';
          else
          cVar1S5S105P013P061P016N033(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='1' AND A(11)='1' AND B( 2)='0' )then
          cVar1S6S105P013P061P016N033(0) <='1';
          else
          cVar1S6S105P013P061P016N033(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S7S105P013N061P032P051(0) <='1';
          else
          cVar1S7S105P013N061P032P051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S8S105P013N061P032P051(0) <='1';
          else
          cVar1S8S105P013N061P032P051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S9S105P013N061P032P051(0) <='1';
          else
          cVar1S9S105P013N061P032P051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S10S105P013N061P032P051(0) <='1';
          else
          cVar1S10S105P013N061P032P051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S11S105P013N061P032N051(0) <='1';
          else
          cVar1S11S105P013N061P032N051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S12S105P013N061P032N051(0) <='1';
          else
          cVar1S12S105P013N061P032N051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S13S105P013N061P032N051(0) <='1';
          else
          cVar1S13S105P013N061P032N051(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='1' AND D( 9)='1' )then
          cVar1S14S105P013N061P032P063(0) <='1';
          else
          cVar1S14S105P013N061P032P063(0) <='0';
          end if;
        if(A( 3)='1' AND E(10)='0' AND B(11)='1' AND D( 9)='0' )then
          cVar1S15S105P013N061P032N063(0) <='1';
          else
          cVar1S15S105P013N061P032N063(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='0' )then
          cVar1S16S105N013P036P002P011(0) <='1';
          else
          cVar1S16S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='0' )then
          cVar1S17S105N013P036P002P011(0) <='1';
          else
          cVar1S17S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='1' )then
          cVar1S18S105N013P036P002P011(0) <='1';
          else
          cVar1S18S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='1' )then
          cVar1S19S105N013P036P002P011(0) <='1';
          else
          cVar1S19S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='1' )then
          cVar1S20S105N013P036P002P011(0) <='1';
          else
          cVar1S20S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='0' AND A( 4)='1' )then
          cVar1S21S105N013P036P002P011(0) <='1';
          else
          cVar1S21S105N013P036P002P011(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='1' AND A(18)='1' AND E( 0)='0' )then
          cVar1S22S105N013P036P002P068(0) <='1';
          else
          cVar1S22S105N013P036P002P068(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='1' AND D(11)='1' )then
          cVar1S23S105N013N036P028P055(0) <='1';
          else
          cVar1S23S105N013N036P028P055(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='1' AND D(11)='1' )then
          cVar1S24S105N013N036P028P055(0) <='1';
          else
          cVar1S24S105N013N036P028P055(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='1' AND D(11)='0' )then
          cVar1S25S105N013N036P028N055(0) <='1';
          else
          cVar1S25S105N013N036P028N055(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='1' AND D(11)='0' )then
          cVar1S26S105N013N036P028N055(0) <='1';
          else
          cVar1S26S105N013N036P028N055(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='0' AND B(14)='1' )then
          cVar1S27S105N013N036N028P026(0) <='1';
          else
          cVar1S27S105N013N036N028P026(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='0' AND B(14)='0' )then
          cVar1S28S105N013N036N028N026(0) <='1';
          else
          cVar1S28S105N013N036N028N026(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='0' AND B(14)='0' )then
          cVar1S29S105N013N036N028N026(0) <='1';
          else
          cVar1S29S105N013N036N028N026(0) <='0';
          end if;
        if(A( 3)='0' AND B( 9)='0' AND B(13)='0' AND B(14)='0' )then
          cVar1S30S105N013N036N028N026(0) <='1';
          else
          cVar1S30S105N013N036N028N026(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S0S106P036P064P002P048(0) <='1';
          else
          cVar1S0S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S1S106P036P064P002P048(0) <='1';
          else
          cVar1S1S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S2S106P036P064P002P048(0) <='1';
          else
          cVar1S2S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S3S106P036P064P002P048(0) <='1';
          else
          cVar1S3S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='1' )then
          cVar1S4S106P036P064P002P048(0) <='1';
          else
          cVar1S4S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='0' AND E( 5)='1' )then
          cVar1S5S106P036P064P002P048(0) <='1';
          else
          cVar1S5S106P036P064P002P048(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='1' AND A(13)='0' )then
          cVar1S6S106P036P064P002P012(0) <='1';
          else
          cVar1S6S106P036P064P002P012(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A(18)='1' AND A(13)='0' )then
          cVar1S7S106P036P064P002P012(0) <='1';
          else
          cVar1S7S106P036P064P002P012(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='1' )then
          cVar1S8S106P036N064P062P015(0) <='1';
          else
          cVar1S8S106P036N064P062P015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='1' )then
          cVar1S9S106P036N064P062P015(0) <='1';
          else
          cVar1S9S106P036N064P062P015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='0' )then
          cVar1S10S106P036N064P062N015(0) <='1';
          else
          cVar1S10S106P036N064P062N015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='0' )then
          cVar1S11S106P036N064P062N015(0) <='1';
          else
          cVar1S11S106P036N064P062N015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='0' )then
          cVar1S12S106P036N064P062N015(0) <='1';
          else
          cVar1S12S106P036N064P062N015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='0' AND A( 2)='0' )then
          cVar1S13S106P036N064P062N015(0) <='1';
          else
          cVar1S13S106P036N064P062N015(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='1' AND D( 6)='0' )then
          cVar1S14S106P036N064P062P042(0) <='1';
          else
          cVar1S14S106P036N064P062P042(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='1' AND D( 6)='0' )then
          cVar1S15S106P036N064P062P042(0) <='1';
          else
          cVar1S15S106P036N064P062P042(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='1' AND D( 6)='0' )then
          cVar1S16S106P036N064P062P042(0) <='1';
          else
          cVar1S16S106P036N064P062P042(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D( 1)='1' AND D( 6)='0' )then
          cVar1S17S106P036N064P062P042(0) <='1';
          else
          cVar1S17S106P036N064P062P042(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='1' AND A(15)='0' )then
          cVar1S18S106P036P005P013P008(0) <='1';
          else
          cVar1S18S106P036P005P013P008(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='1' AND A(15)='0' )then
          cVar1S19S106P036P005P013P008(0) <='1';
          else
          cVar1S19S106P036P005P013P008(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='1' AND A(15)='0' )then
          cVar1S20S106P036P005P013P008(0) <='1';
          else
          cVar1S20S106P036P005P013P008(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='1' AND A(15)='0' )then
          cVar1S21S106P036P005P013P008(0) <='1';
          else
          cVar1S21S106P036P005P013P008(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='1' AND A(15)='1' )then
          cVar1S22S106P036P005P013P008(0) <='1';
          else
          cVar1S22S106P036P005P013P008(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='0' AND E(10)='0' )then
          cVar1S23S106P036P005N013P061(0) <='1';
          else
          cVar1S23S106P036P005N013P061(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='0' AND E(10)='0' )then
          cVar1S24S106P036P005N013P061(0) <='1';
          else
          cVar1S24S106P036P005N013P061(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='0' AND E(10)='1' )then
          cVar1S25S106P036P005N013P061(0) <='1';
          else
          cVar1S25S106P036P005N013P061(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='0' AND E(10)='1' )then
          cVar1S26S106P036P005N013P061(0) <='1';
          else
          cVar1S26S106P036P005N013P061(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 3)='0' AND E(10)='1' )then
          cVar1S27S106P036P005N013P061(0) <='1';
          else
          cVar1S27S106P036P005N013P061(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND B(17)='1' )then
          cVar1S28S106P036P005P031P020nsss(0) <='1';
          else
          cVar1S28S106P036P005P031P020nsss(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND B(17)='0' )then
          cVar1S29S106P036P005P031N020(0) <='1';
          else
          cVar1S29S106P036P005P031N020(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND B(17)='0' )then
          cVar1S30S106P036P005P031N020(0) <='1';
          else
          cVar1S30S106P036P005P031N020(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND B(17)='0' )then
          cVar1S31S106P036P005P031N020(0) <='1';
          else
          cVar1S31S106P036P005P031N020(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S0S107P036P005P019P047(0) <='1';
          else
          cVar1S0S107P036P005P019P047(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S1S107P036P005P019P047(0) <='1';
          else
          cVar1S1S107P036P005P019P047(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='1' AND D(13)='0' )then
          cVar1S2S107P036P005P019P047(0) <='1';
          else
          cVar1S2S107P036P005P019P047(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='1' AND D(13)='1' )then
          cVar1S3S107P036P005P019P047(0) <='1';
          else
          cVar1S3S107P036P005P019P047(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='0' )then
          cVar1S4S107P036P005N019P048(0) <='1';
          else
          cVar1S4S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='0' )then
          cVar1S5S107P036P005N019P048(0) <='1';
          else
          cVar1S5S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='0' )then
          cVar1S6S107P036P005N019P048(0) <='1';
          else
          cVar1S6S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='0' )then
          cVar1S7S107P036P005N019P048(0) <='1';
          else
          cVar1S7S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='1' )then
          cVar1S8S107P036P005N019P048(0) <='1';
          else
          cVar1S8S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='0' AND A( 0)='0' AND E( 5)='1' )then
          cVar1S9S107P036P005N019P048(0) <='1';
          else
          cVar1S9S107P036P005N019P048(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND E( 8)='1' )then
          cVar1S10S107P036P005P031P069(0) <='1';
          else
          cVar1S10S107P036P005P031P069(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND E( 8)='1' )then
          cVar1S11S107P036P005P031P069(0) <='1';
          else
          cVar1S11S107P036P005P031P069(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND E( 8)='0' )then
          cVar1S12S107P036P005P031N069(0) <='1';
          else
          cVar1S12S107P036P005P031N069(0) <='0';
          end if;
        if(B( 9)='1' AND A( 7)='1' AND B( 3)='0' AND E( 8)='0' )then
          cVar1S13S107P036P005P031N069(0) <='1';
          else
          cVar1S13S107P036P005P031N069(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='1' AND D(10)='1' )then
          cVar1S14S107N036P064P019P059(0) <='1';
          else
          cVar1S14S107N036P064P019P059(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='1' AND D(10)='1' )then
          cVar1S15S107N036P064P019P059(0) <='1';
          else
          cVar1S15S107N036P064P019P059(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='1' AND D(10)='0' )then
          cVar1S16S107N036P064P019N059(0) <='1';
          else
          cVar1S16S107N036P064P019N059(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='1' AND D(10)='0' )then
          cVar1S17S107N036P064P019N059(0) <='1';
          else
          cVar1S17S107N036P064P019N059(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='1' AND D(10)='0' )then
          cVar1S18S107N036P064P019N059(0) <='1';
          else
          cVar1S18S107N036P064P019N059(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='0' )then
          cVar1S19S107N036P064N019P056(0) <='1';
          else
          cVar1S19S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='0' )then
          cVar1S20S107N036P064N019P056(0) <='1';
          else
          cVar1S20S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='1' )then
          cVar1S21S107N036P064N019P056(0) <='1';
          else
          cVar1S21S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='1' )then
          cVar1S22S107N036P064N019P056(0) <='1';
          else
          cVar1S22S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='1' )then
          cVar1S23S107N036P064N019P056(0) <='1';
          else
          cVar1S23S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='1' AND A( 0)='0' AND E( 3)='1' )then
          cVar1S24S107N036P064N019P056(0) <='1';
          else
          cVar1S24S107N036P064N019P056(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='1' AND E(11)='0' )then
          cVar1S25S107N036N064P051P057(0) <='1';
          else
          cVar1S25S107N036N064P051P057(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='1' AND E(11)='0' )then
          cVar1S26S107N036N064P051P057(0) <='1';
          else
          cVar1S26S107N036N064P051P057(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='1' AND E(11)='0' )then
          cVar1S27S107N036N064P051P057(0) <='1';
          else
          cVar1S27S107N036N064P051P057(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='1' AND E(11)='1' )then
          cVar1S28S107N036N064P051P057(0) <='1';
          else
          cVar1S28S107N036N064P051P057(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='1' AND E(11)='1' )then
          cVar1S29S107N036N064P051P057(0) <='1';
          else
          cVar1S29S107N036N064P051P057(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='0' AND E(12)='0' )then
          cVar1S30S107N036N064N051P053(0) <='1';
          else
          cVar1S30S107N036N064N051P053(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='0' AND E(12)='0' )then
          cVar1S31S107N036N064N051P053(0) <='1';
          else
          cVar1S31S107N036N064N051P053(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='0' AND E(12)='0' )then
          cVar1S32S107N036N064N051P053(0) <='1';
          else
          cVar1S32S107N036N064N051P053(0) <='0';
          end if;
        if(B( 9)='0' AND E( 1)='0' AND D(12)='0' AND E(12)='1' )then
          cVar1S33S107N036N064N051P053(0) <='1';
          else
          cVar1S33S107N036N064N051P053(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='0' )then
          cVar1S0S108P064P012P031P054(0) <='1';
          else
          cVar1S0S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='0' )then
          cVar1S1S108P064P012P031P054(0) <='1';
          else
          cVar1S1S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='0' )then
          cVar1S2S108P064P012P031P054(0) <='1';
          else
          cVar1S2S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='1' )then
          cVar1S3S108P064P012P031P054(0) <='1';
          else
          cVar1S3S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='1' )then
          cVar1S4S108P064P012P031P054(0) <='1';
          else
          cVar1S4S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='1' )then
          cVar1S5S108P064P012P031P054(0) <='1';
          else
          cVar1S5S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='0' AND D( 3)='1' )then
          cVar1S6S108P064P012P031P054(0) <='1';
          else
          cVar1S6S108P064P012P031P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='1' AND A( 7)='0' )then
          cVar1S7S108P064P012P031P005(0) <='1';
          else
          cVar1S7S108P064P012P031P005(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='1' AND A( 7)='0' )then
          cVar1S8S108P064P012P031P005(0) <='1';
          else
          cVar1S8S108P064P012P031P005(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='1' AND A( 7)='0' )then
          cVar1S9S108P064P012P031P005(0) <='1';
          else
          cVar1S9S108P064P012P031P005(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='0' AND B( 3)='1' AND A( 7)='1' )then
          cVar1S10S108P064P012P031P005(0) <='1';
          else
          cVar1S10S108P064P012P031P005(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='1' AND B(11)='0' )then
          cVar1S11S108P064P012P030P032(0) <='1';
          else
          cVar1S11S108P064P012P030P032(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='1' AND B(11)='0' )then
          cVar1S12S108P064P012P030P032(0) <='1';
          else
          cVar1S12S108P064P012P030P032(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='1' AND B(11)='0' )then
          cVar1S13S108P064P012P030P032(0) <='1';
          else
          cVar1S13S108P064P012P030P032(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='1' AND B(11)='1' )then
          cVar1S14S108P064P012P030P032(0) <='1';
          else
          cVar1S14S108P064P012P030P032(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='1' AND B(11)='1' )then
          cVar1S15S108P064P012P030P032(0) <='1';
          else
          cVar1S15S108P064P012P030P032(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='0' AND D( 3)='1' )then
          cVar1S16S108P064P012N030P054(0) <='1';
          else
          cVar1S16S108P064P012N030P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='0' AND D( 3)='1' )then
          cVar1S17S108P064P012N030P054(0) <='1';
          else
          cVar1S17S108P064P012N030P054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='0' AND D( 3)='0' )then
          cVar1S18S108P064P012N030N054(0) <='1';
          else
          cVar1S18S108P064P012N030N054(0) <='0';
          end if;
        if(E( 1)='0' AND A(13)='1' AND B(12)='0' AND D( 3)='0' )then
          cVar1S19S108P064P012N030N054(0) <='1';
          else
          cVar1S19S108P064P012N030N054(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='1' )then
          cVar1S20S108P064P068P062P066(0) <='1';
          else
          cVar1S20S108P064P068P062P066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='1' )then
          cVar1S21S108P064P068P062P066(0) <='1';
          else
          cVar1S21S108P064P068P062P066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='1' )then
          cVar1S22S108P064P068P062P066(0) <='1';
          else
          cVar1S22S108P064P068P062P066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='0' )then
          cVar1S23S108P064P068P062N066(0) <='1';
          else
          cVar1S23S108P064P068P062N066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='0' )then
          cVar1S24S108P064P068P062N066(0) <='1';
          else
          cVar1S24S108P064P068P062N066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='0' AND D( 0)='0' )then
          cVar1S25S108P064P068P062N066(0) <='1';
          else
          cVar1S25S108P064P068P062N066(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='1' AND E(14)='1' )then
          cVar1S26S108P064P068P062P045(0) <='1';
          else
          cVar1S26S108P064P068P062P045(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='1' AND E(14)='1' )then
          cVar1S27S108P064P068P062P045(0) <='1';
          else
          cVar1S27S108P064P068P062P045(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='1' AND E(14)='0' )then
          cVar1S28S108P064P068P062N045(0) <='1';
          else
          cVar1S28S108P064P068P062N045(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D( 1)='1' AND E(14)='0' )then
          cVar1S29S108P064P068P062N045(0) <='1';
          else
          cVar1S29S108P064P068P062N045(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='1' AND B( 1)='1' )then
          cVar1S30S108P064P068P012P035(0) <='1';
          else
          cVar1S30S108P064P068P012P035(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='1' AND B( 1)='1' )then
          cVar1S31S108P064P068P012P035(0) <='1';
          else
          cVar1S31S108P064P068P012P035(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='1' AND B( 1)='1' )then
          cVar1S32S108P064P068P012P035(0) <='1';
          else
          cVar1S32S108P064P068P012P035(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='1' AND B( 1)='0' )then
          cVar1S33S108P064P068P012N035(0) <='1';
          else
          cVar1S33S108P064P068P012N035(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='1' AND B( 1)='0' )then
          cVar1S34S108P064P068P012N035(0) <='1';
          else
          cVar1S34S108P064P068P012N035(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='0' AND A( 0)='1' )then
          cVar1S35S108P064P068N012P019(0) <='1';
          else
          cVar1S35S108P064P068N012P019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='0' AND A( 0)='1' )then
          cVar1S36S108P064P068N012P019(0) <='1';
          else
          cVar1S36S108P064P068N012P019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='0' AND A( 0)='0' )then
          cVar1S37S108P064P068N012N019(0) <='1';
          else
          cVar1S37S108P064P068N012N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='0' AND A( 0)='0' )then
          cVar1S38S108P064P068N012N019(0) <='1';
          else
          cVar1S38S108P064P068N012N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND A(13)='0' AND A( 0)='0' )then
          cVar1S39S108P064P068N012N019(0) <='1';
          else
          cVar1S39S108P064P068N012N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='0' AND E( 3)='0' )then
          cVar1S0S109P064P068P055P056(0) <='1';
          else
          cVar1S0S109P064P068P055P056(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='0' AND E( 3)='0' )then
          cVar1S1S109P064P068P055P056(0) <='1';
          else
          cVar1S1S109P064P068P055P056(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='0' AND E( 3)='0' )then
          cVar1S2S109P064P068P055P056(0) <='1';
          else
          cVar1S2S109P064P068P055P056(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='0' AND E( 3)='0' )then
          cVar1S3S109P064P068P055P056(0) <='1';
          else
          cVar1S3S109P064P068P055P056(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='0' AND E( 3)='1' )then
          cVar1S4S109P064P068P055P056(0) <='1';
          else
          cVar1S4S109P064P068P055P056(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='1' AND E( 2)='0' )then
          cVar1S5S109P064P068P055P060(0) <='1';
          else
          cVar1S5S109P064P068P055P060(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='1' AND E( 2)='0' )then
          cVar1S6S109P064P068P055P060(0) <='1';
          else
          cVar1S6S109P064P068P055P060(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='0' AND D(11)='1' AND E( 2)='0' )then
          cVar1S7S109P064P068P055P060(0) <='1';
          else
          cVar1S7S109P064P068P055P060(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND D(12)='0' AND A( 0)='1' )then
          cVar1S8S109P064P068P051P019(0) <='1';
          else
          cVar1S8S109P064P068P051P019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND D(12)='0' AND A( 0)='0' )then
          cVar1S9S109P064P068P051N019(0) <='1';
          else
          cVar1S9S109P064P068P051N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND D(12)='0' AND A( 0)='0' )then
          cVar1S10S109P064P068P051N019(0) <='1';
          else
          cVar1S10S109P064P068P051N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND D(12)='0' AND A( 0)='0' )then
          cVar1S11S109P064P068P051N019(0) <='1';
          else
          cVar1S11S109P064P068P051N019(0) <='0';
          end if;
        if(E( 1)='1' AND E( 0)='1' AND D(12)='1' AND A( 1)='1' )then
          cVar1S12S109P064P068P051P017nsss(0) <='1';
          else
          cVar1S12S109P064P068P051P017nsss(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='1' )then
          cVar1S13S109N064P054P040P015(0) <='1';
          else
          cVar1S13S109N064P054P040P015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='1' )then
          cVar1S14S109N064P054P040P015(0) <='1';
          else
          cVar1S14S109N064P054P040P015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='1' )then
          cVar1S15S109N064P054P040P015(0) <='1';
          else
          cVar1S15S109N064P054P040P015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='1' )then
          cVar1S16S109N064P054P040P015(0) <='1';
          else
          cVar1S16S109N064P054P040P015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='0' )then
          cVar1S17S109N064P054P040N015(0) <='1';
          else
          cVar1S17S109N064P054P040N015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='0' )then
          cVar1S18S109N064P054P040N015(0) <='1';
          else
          cVar1S18S109N064P054P040N015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='1' AND E( 7)='0' AND A( 2)='0' )then
          cVar1S19S109N064P054P040N015(0) <='1';
          else
          cVar1S19S109N064P054P040N015(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='1' )then
          cVar1S20S109N064N054P022P043(0) <='1';
          else
          cVar1S20S109N064N054P022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='1' )then
          cVar1S21S109N064N054P022P043(0) <='1';
          else
          cVar1S21S109N064N054P022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='1' )then
          cVar1S22S109N064N054P022P043(0) <='1';
          else
          cVar1S22S109N064N054P022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='0' )then
          cVar1S23S109N064N054P022N043(0) <='1';
          else
          cVar1S23S109N064N054P022N043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='0' )then
          cVar1S24S109N064N054P022N043(0) <='1';
          else
          cVar1S24S109N064N054P022N043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='1' AND D(14)='0' )then
          cVar1S25S109N064N054P022N043(0) <='1';
          else
          cVar1S25S109N064N054P022N043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='0' AND D(14)='0' )then
          cVar1S26S109N064N054N022P043(0) <='1';
          else
          cVar1S26S109N064N054N022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='0' AND D(14)='0' )then
          cVar1S27S109N064N054N022P043(0) <='1';
          else
          cVar1S27S109N064N054N022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='0' AND D(14)='0' )then
          cVar1S28S109N064N054N022P043(0) <='1';
          else
          cVar1S28S109N064N054N022P043(0) <='0';
          end if;
        if(E( 1)='0' AND D( 3)='0' AND B(16)='0' AND D(14)='1' )then
          cVar1S29S109N064N054N022P043(0) <='1';
          else
          cVar1S29S109N064N054N022P043(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='0' AND B( 5)='0' )then
          cVar1S0S110P064P056P052P027(0) <='1';
          else
          cVar1S0S110P064P056P052P027(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='0' AND B( 5)='0' )then
          cVar1S1S110P064P056P052P027(0) <='1';
          else
          cVar1S1S110P064P056P052P027(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='0' AND B( 5)='1' )then
          cVar1S2S110P064P056P052P027(0) <='1';
          else
          cVar1S2S110P064P056P052P027(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='1' AND A( 5)='1' )then
          cVar1S3S110P064P056P052P009nsss(0) <='1';
          else
          cVar1S3S110P064P056P052P009nsss(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S4S110P064P056P052N009(0) <='1';
          else
          cVar1S4S110P064P056P052N009(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='1' AND E( 4)='1' AND A( 5)='0' )then
          cVar1S5S110P064P056P052N009(0) <='1';
          else
          cVar1S5S110P064P056P052N009(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='0' )then
          cVar1S6S110P064N056P026P049(0) <='1';
          else
          cVar1S6S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='0' )then
          cVar1S7S110P064N056P026P049(0) <='1';
          else
          cVar1S7S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='0' )then
          cVar1S8S110P064N056P026P049(0) <='1';
          else
          cVar1S8S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='0' )then
          cVar1S9S110P064N056P026P049(0) <='1';
          else
          cVar1S9S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='1' )then
          cVar1S10S110P064N056P026P049(0) <='1';
          else
          cVar1S10S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='1' )then
          cVar1S11S110P064N056P026P049(0) <='1';
          else
          cVar1S11S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='0' AND E(13)='1' )then
          cVar1S12S110P064N056P026P049(0) <='1';
          else
          cVar1S12S110P064N056P026P049(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='1' )then
          cVar1S13S110P064N056P026P050(0) <='1';
          else
          cVar1S13S110P064N056P026P050(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='1' )then
          cVar1S14S110P064N056P026P050(0) <='1';
          else
          cVar1S14S110P064N056P026P050(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='1' )then
          cVar1S15S110P064N056P026P050(0) <='1';
          else
          cVar1S15S110P064N056P026P050(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='0' )then
          cVar1S16S110P064N056P026N050(0) <='1';
          else
          cVar1S16S110P064N056P026N050(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='0' )then
          cVar1S17S110P064N056P026N050(0) <='1';
          else
          cVar1S17S110P064N056P026N050(0) <='0';
          end if;
        if(E( 1)='0' AND E( 3)='0' AND B(14)='1' AND D( 4)='0' )then
          cVar1S18S110P064N056P026N050(0) <='1';
          else
          cVar1S18S110P064N056P026N050(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='1' AND D(13)='0' AND B(14)='0' )then
          cVar1S19S110P064P013P047P026(0) <='1';
          else
          cVar1S19S110P064P013P047P026(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='1' AND D(13)='0' AND B(14)='0' )then
          cVar1S20S110P064P013P047P026(0) <='1';
          else
          cVar1S20S110P064P013P047P026(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='1' AND D(13)='0' AND B(14)='0' )then
          cVar1S21S110P064P013P047P026(0) <='1';
          else
          cVar1S21S110P064P013P047P026(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='1' AND D(13)='0' AND B(14)='0' )then
          cVar1S22S110P064P013P047P026(0) <='1';
          else
          cVar1S22S110P064P013P047P026(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='1' AND D(13)='0' AND B(14)='1' )then
          cVar1S23S110P064P013P047P026(0) <='1';
          else
          cVar1S23S110P064P013P047P026(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='0' AND B( 2)='0' AND B(16)='0' )then
          cVar1S24S110P064N013P033P022(0) <='1';
          else
          cVar1S24S110P064N013P033P022(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='0' AND B( 2)='0' AND B(16)='1' )then
          cVar1S25S110P064N013P033P022(0) <='1';
          else
          cVar1S25S110P064N013P033P022(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='0' AND B( 2)='1' AND D( 4)='0' )then
          cVar1S26S110P064N013P033P050(0) <='1';
          else
          cVar1S26S110P064N013P033P050(0) <='0';
          end if;
        if(E( 1)='1' AND A( 3)='0' AND B( 2)='1' AND D( 4)='0' )then
          cVar1S27S110P064N013P033P050(0) <='1';
          else
          cVar1S27S110P064N013P033P050(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='0' AND A(10)='0' )then
          cVar1S0S111P064P033P041P018(0) <='1';
          else
          cVar1S0S111P064P033P041P018(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='0' AND A(10)='0' )then
          cVar1S1S111P064P033P041P018(0) <='1';
          else
          cVar1S1S111P064P033P041P018(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='0' AND A(10)='0' )then
          cVar1S2S111P064P033P041P018(0) <='1';
          else
          cVar1S2S111P064P033P041P018(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='0' AND A(10)='1' )then
          cVar1S3S111P064P033P041P018(0) <='1';
          else
          cVar1S3S111P064P033P041P018(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='0' AND A(10)='1' )then
          cVar1S4S111P064P033P041P018(0) <='1';
          else
          cVar1S4S111P064P033P041P018(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='0' AND E(15)='1' AND A( 8)='1' )then
          cVar1S5S111P064P033P041P003nsss(0) <='1';
          else
          cVar1S5S111P064P033P041P003nsss(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='1' AND E( 5)='0' AND D( 4)='0' )then
          cVar1S6S111P064P033P048P050(0) <='1';
          else
          cVar1S6S111P064P033P048P050(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='1' AND E( 5)='0' AND D( 4)='0' )then
          cVar1S7S111P064P033P048P050(0) <='1';
          else
          cVar1S7S111P064P033P048P050(0) <='0';
          end if;
        if(E( 1)='1' AND B( 2)='1' AND E( 5)='0' AND D( 4)='0' )then
          cVar1S8S111P064P033P048P050(0) <='1';
          else
          cVar1S8S111P064P033P048P050(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S9S111N064P016P047P024(0) <='1';
          else
          cVar1S9S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S10S111N064P016P047P024(0) <='1';
          else
          cVar1S10S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S11S111N064P016P047P024(0) <='1';
          else
          cVar1S11S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='0' )then
          cVar1S12S111N064P016P047P024(0) <='1';
          else
          cVar1S12S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='1' )then
          cVar1S13S111N064P016P047P024(0) <='1';
          else
          cVar1S13S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='0' AND B(15)='1' )then
          cVar1S14S111N064P016P047P024(0) <='1';
          else
          cVar1S14S111N064P016P047P024(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='1' AND B(10)='1' )then
          cVar1S15S111N064P016P047P034(0) <='1';
          else
          cVar1S15S111N064P016P047P034(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='1' AND B(10)='0' )then
          cVar1S16S111N064P016P047N034(0) <='1';
          else
          cVar1S16S111N064P016P047N034(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='1' AND D(13)='1' AND B(10)='0' )then
          cVar1S17S111N064P016P047N034(0) <='1';
          else
          cVar1S17S111N064P016P047N034(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='1' )then
          cVar1S18S111N064N016P018P015(0) <='1';
          else
          cVar1S18S111N064N016P018P015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='1' )then
          cVar1S19S111N064N016P018P015(0) <='1';
          else
          cVar1S19S111N064N016P018P015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='1' )then
          cVar1S20S111N064N016P018P015(0) <='1';
          else
          cVar1S20S111N064N016P018P015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='1' )then
          cVar1S21S111N064N016P018P015(0) <='1';
          else
          cVar1S21S111N064N016P018P015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='0' )then
          cVar1S22S111N064N016P018N015(0) <='1';
          else
          cVar1S22S111N064N016P018N015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='0' )then
          cVar1S23S111N064N016P018N015(0) <='1';
          else
          cVar1S23S111N064N016P018N015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='1' AND A( 2)='0' )then
          cVar1S24S111N064N016P018N015(0) <='1';
          else
          cVar1S24S111N064N016P018N015(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='0' AND D(10)='1' )then
          cVar1S25S111N064N016N018P059(0) <='1';
          else
          cVar1S25S111N064N016N018P059(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='0' AND D(10)='0' )then
          cVar1S26S111N064N016N018N059(0) <='1';
          else
          cVar1S26S111N064N016N018N059(0) <='0';
          end if;
        if(E( 1)='0' AND A(11)='0' AND A(10)='0' AND D(10)='0' )then
          cVar1S27S111N064N016N018N059(0) <='1';
          else
          cVar1S27S111N064N016N018N059(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='0' )then
          cVar1S0S112P018P016P027P066(0) <='1';
          else
          cVar1S0S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='0' )then
          cVar1S1S112P018P016P027P066(0) <='1';
          else
          cVar1S1S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='0' )then
          cVar1S2S112P018P016P027P066(0) <='1';
          else
          cVar1S2S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='0' )then
          cVar1S3S112P018P016P027P066(0) <='1';
          else
          cVar1S3S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='1' )then
          cVar1S4S112P018P016P027P066(0) <='1';
          else
          cVar1S4S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='1' )then
          cVar1S5S112P018P016P027P066(0) <='1';
          else
          cVar1S5S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='1' )then
          cVar1S6S112P018P016P027P066(0) <='1';
          else
          cVar1S6S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='0' AND D( 0)='1' )then
          cVar1S7S112P018P016P027P066(0) <='1';
          else
          cVar1S7S112P018P016P027P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='1' )then
          cVar1S8S112P018P016P027P009(0) <='1';
          else
          cVar1S8S112P018P016P027P009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='1' )then
          cVar1S9S112P018P016P027P009(0) <='1';
          else
          cVar1S9S112P018P016P027P009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='1' )then
          cVar1S10S112P018P016P027P009(0) <='1';
          else
          cVar1S10S112P018P016P027P009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='0' )then
          cVar1S11S112P018P016P027N009(0) <='1';
          else
          cVar1S11S112P018P016P027N009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='0' )then
          cVar1S12S112P018P016P027N009(0) <='1';
          else
          cVar1S12S112P018P016P027N009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B( 5)='1' AND A( 5)='0' )then
          cVar1S13S112P018P016P027N009(0) <='1';
          else
          cVar1S13S112P018P016P027N009(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='1' AND E( 9)='0' )then
          cVar1S14S112P018P016P059P065(0) <='1';
          else
          cVar1S14S112P018P016P059P065(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='1' AND E( 9)='0' )then
          cVar1S15S112P018P016P059P065(0) <='1';
          else
          cVar1S15S112P018P016P059P065(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='1' AND E( 9)='1' )then
          cVar1S16S112P018P016P059P065(0) <='1';
          else
          cVar1S16S112P018P016P059P065(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='0' AND D( 0)='0' )then
          cVar1S17S112P018P016N059P066(0) <='1';
          else
          cVar1S17S112P018P016N059P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='0' AND D( 0)='0' )then
          cVar1S18S112P018P016N059P066(0) <='1';
          else
          cVar1S18S112P018P016N059P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='0' AND D( 0)='0' )then
          cVar1S19S112P018P016N059P066(0) <='1';
          else
          cVar1S19S112P018P016N059P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='0' AND D( 0)='1' )then
          cVar1S20S112P018P016N059P066(0) <='1';
          else
          cVar1S20S112P018P016N059P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND D(10)='0' AND D( 0)='1' )then
          cVar1S21S112P018P016N059P066(0) <='1';
          else
          cVar1S21S112P018P016N059P066(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='1' AND E( 7)='0' AND E( 9)='0' )then
          cVar1S22S112N018P054P040P065(0) <='1';
          else
          cVar1S22S112N018P054P040P065(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='1' AND E( 7)='0' AND E( 9)='0' )then
          cVar1S23S112N018P054P040P065(0) <='1';
          else
          cVar1S23S112N018P054P040P065(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='1' AND E( 7)='0' AND E( 9)='0' )then
          cVar1S24S112N018P054P040P065(0) <='1';
          else
          cVar1S24S112N018P054P040P065(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='1' AND E( 7)='0' AND E( 9)='1' )then
          cVar1S25S112N018P054P040P065(0) <='1';
          else
          cVar1S25S112N018P054P040P065(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='1' AND E( 7)='0' AND E( 9)='1' )then
          cVar1S26S112N018P054P040P065(0) <='1';
          else
          cVar1S26S112N018P054P040P065(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='1' )then
          cVar1S27S112N018N054P014P055(0) <='1';
          else
          cVar1S27S112N018N054P014P055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='1' )then
          cVar1S28S112N018N054P014P055(0) <='1';
          else
          cVar1S28S112N018N054P014P055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='0' )then
          cVar1S29S112N018N054P014N055(0) <='1';
          else
          cVar1S29S112N018N054P014N055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='0' )then
          cVar1S30S112N018N054P014N055(0) <='1';
          else
          cVar1S30S112N018N054P014N055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='0' )then
          cVar1S31S112N018N054P014N055(0) <='1';
          else
          cVar1S31S112N018N054P014N055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='0' AND D(11)='0' )then
          cVar1S32S112N018N054P014N055(0) <='1';
          else
          cVar1S32S112N018N054P014N055(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='1' AND B( 3)='0' )then
          cVar1S33S112N018N054P014P031(0) <='1';
          else
          cVar1S33S112N018N054P014P031(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='1' AND B( 3)='0' )then
          cVar1S34S112N018N054P014P031(0) <='1';
          else
          cVar1S34S112N018N054P014P031(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='1' AND B( 3)='0' )then
          cVar1S35S112N018N054P014P031(0) <='1';
          else
          cVar1S35S112N018N054P014P031(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='1' AND B( 3)='0' )then
          cVar1S36S112N018N054P014P031(0) <='1';
          else
          cVar1S36S112N018N054P014P031(0) <='0';
          end if;
        if(A(10)='0' AND D( 3)='0' AND A(12)='1' AND B( 3)='1' )then
          cVar1S37S112N018N054P014P031(0) <='1';
          else
          cVar1S37S112N018N054P014P031(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='0' )then
          cVar1S0S113P014P018P056P011(0) <='1';
          else
          cVar1S0S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='0' )then
          cVar1S1S113P014P018P056P011(0) <='1';
          else
          cVar1S1S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='0' )then
          cVar1S2S113P014P018P056P011(0) <='1';
          else
          cVar1S2S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='0' )then
          cVar1S3S113P014P018P056P011(0) <='1';
          else
          cVar1S3S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='1' )then
          cVar1S4S113P014P018P056P011(0) <='1';
          else
          cVar1S4S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='1' )then
          cVar1S5S113P014P018P056P011(0) <='1';
          else
          cVar1S5S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='1' )then
          cVar1S6S113P014P018P056P011(0) <='1';
          else
          cVar1S6S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='0' AND A( 4)='1' )then
          cVar1S7S113P014P018P056P011(0) <='1';
          else
          cVar1S7S113P014P018P056P011(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='1' AND A( 1)='1' )then
          cVar1S8S113P014P018P056P017(0) <='1';
          else
          cVar1S8S113P014P018P056P017(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='1' AND A( 1)='1' )then
          cVar1S9S113P014P018P056P017(0) <='1';
          else
          cVar1S9S113P014P018P056P017(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='1' AND A( 1)='0' )then
          cVar1S10S113P014P018P056N017(0) <='1';
          else
          cVar1S10S113P014P018P056N017(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='1' AND A( 1)='0' )then
          cVar1S11S113P014P018P056N017(0) <='1';
          else
          cVar1S11S113P014P018P056N017(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='0' AND E( 3)='1' AND A( 1)='0' )then
          cVar1S12S113P014P018P056N017(0) <='1';
          else
          cVar1S12S113P014P018P056N017(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='0' )then
          cVar1S13S113P014P018P067P050(0) <='1';
          else
          cVar1S13S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='0' )then
          cVar1S14S113P014P018P067P050(0) <='1';
          else
          cVar1S14S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='0' )then
          cVar1S15S113P014P018P067P050(0) <='1';
          else
          cVar1S15S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='0' )then
          cVar1S16S113P014P018P067P050(0) <='1';
          else
          cVar1S16S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='1' )then
          cVar1S17S113P014P018P067P050(0) <='1';
          else
          cVar1S17S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='1' )then
          cVar1S18S113P014P018P067P050(0) <='1';
          else
          cVar1S18S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='1' AND D( 4)='1' )then
          cVar1S19S113P014P018P067P050(0) <='1';
          else
          cVar1S19S113P014P018P067P050(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='1' )then
          cVar1S20S113P014P018N067P012(0) <='1';
          else
          cVar1S20S113P014P018N067P012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='1' )then
          cVar1S21S113P014P018N067P012(0) <='1';
          else
          cVar1S21S113P014P018N067P012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='1' )then
          cVar1S22S113P014P018N067P012(0) <='1';
          else
          cVar1S22S113P014P018N067P012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='1' )then
          cVar1S23S113P014P018N067P012(0) <='1';
          else
          cVar1S23S113P014P018N067P012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='0' )then
          cVar1S24S113P014P018N067N012(0) <='1';
          else
          cVar1S24S113P014P018N067N012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='0' )then
          cVar1S25S113P014P018N067N012(0) <='1';
          else
          cVar1S25S113P014P018N067N012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='0' )then
          cVar1S26S113P014P018N067N012(0) <='1';
          else
          cVar1S26S113P014P018N067N012(0) <='0';
          end if;
        if(A(12)='0' AND A(10)='1' AND D( 8)='0' AND A(13)='0' )then
          cVar1S27S113P014P018N067N012(0) <='1';
          else
          cVar1S27S113P014P018N067N012(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='0' AND B( 7)='1' )then
          cVar1S28S113P014P018P022P023(0) <='1';
          else
          cVar1S28S113P014P018P022P023(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='0' AND B( 7)='0' )then
          cVar1S29S113P014P018P022N023(0) <='1';
          else
          cVar1S29S113P014P018P022N023(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='0' AND B( 7)='0' )then
          cVar1S30S113P014P018P022N023(0) <='1';
          else
          cVar1S30S113P014P018P022N023(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='0' AND B( 7)='0' )then
          cVar1S31S113P014P018P022N023(0) <='1';
          else
          cVar1S31S113P014P018P022N023(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='0' AND B( 7)='0' )then
          cVar1S32S113P014P018P022N023(0) <='1';
          else
          cVar1S32S113P014P018P022N023(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='1' AND B( 0)='1' )then
          cVar1S33S113P014P018P022P037nsss(0) <='1';
          else
          cVar1S33S113P014P018P022P037nsss(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='1' AND B(16)='1' AND B( 0)='0' )then
          cVar1S34S113P014P018P022N037(0) <='1';
          else
          cVar1S34S113P014P018P022N037(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='1' )then
          cVar1S35S113P014N018P036P035(0) <='1';
          else
          cVar1S35S113P014N018P036P035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='1' )then
          cVar1S36S113P014N018P036P035(0) <='1';
          else
          cVar1S36S113P014N018P036P035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='1' )then
          cVar1S37S113P014N018P036P035(0) <='1';
          else
          cVar1S37S113P014N018P036P035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='1' )then
          cVar1S38S113P014N018P036P035(0) <='1';
          else
          cVar1S38S113P014N018P036P035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='0' )then
          cVar1S39S113P014N018P036N035(0) <='1';
          else
          cVar1S39S113P014N018P036N035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='0' )then
          cVar1S40S113P014N018P036N035(0) <='1';
          else
          cVar1S40S113P014N018P036N035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='0' )then
          cVar1S41S113P014N018P036N035(0) <='1';
          else
          cVar1S41S113P014N018P036N035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='0' AND B( 1)='0' )then
          cVar1S42S113P014N018P036N035(0) <='1';
          else
          cVar1S42S113P014N018P036N035(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='1' AND E(12)='0' )then
          cVar1S43S113P014N018P036P053(0) <='1';
          else
          cVar1S43S113P014N018P036P053(0) <='0';
          end if;
        if(A(12)='1' AND A(10)='0' AND B( 9)='1' AND E(12)='0' )then
          cVar1S44S113P014N018P036P053(0) <='1';
          else
          cVar1S44S113P014N018P036P053(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='0' AND B(11)='1' )then
          cVar1S0S114P018P064P007P032(0) <='1';
          else
          cVar1S0S114P018P064P007P032(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='0' AND B(11)='0' )then
          cVar1S1S114P018P064P007N032(0) <='1';
          else
          cVar1S1S114P018P064P007N032(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='0' AND B(11)='0' )then
          cVar1S2S114P018P064P007N032(0) <='1';
          else
          cVar1S2S114P018P064P007N032(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='0' AND B(11)='0' )then
          cVar1S3S114P018P064P007N032(0) <='1';
          else
          cVar1S3S114P018P064P007N032(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='0' AND B(11)='0' )then
          cVar1S4S114P018P064P007N032(0) <='1';
          else
          cVar1S4S114P018P064P007N032(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='1' AND D(10)='0' )then
          cVar1S5S114P018P064P007P059(0) <='1';
          else
          cVar1S5S114P018P064P007P059(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='1' AND D(10)='0' )then
          cVar1S6S114P018P064P007P059(0) <='1';
          else
          cVar1S6S114P018P064P007P059(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='1' AND A( 6)='1' AND D(10)='0' )then
          cVar1S7S114P018P064P007P059(0) <='1';
          else
          cVar1S7S114P018P064P007P059(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='1' )then
          cVar1S8S114P018N064P050P034(0) <='1';
          else
          cVar1S8S114P018N064P050P034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='1' )then
          cVar1S9S114P018N064P050P034(0) <='1';
          else
          cVar1S9S114P018N064P050P034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='0' )then
          cVar1S10S114P018N064P050N034(0) <='1';
          else
          cVar1S10S114P018N064P050N034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='0' )then
          cVar1S11S114P018N064P050N034(0) <='1';
          else
          cVar1S11S114P018N064P050N034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='0' )then
          cVar1S12S114P018N064P050N034(0) <='1';
          else
          cVar1S12S114P018N064P050N034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='0' AND B(10)='0' )then
          cVar1S13S114P018N064P050N034(0) <='1';
          else
          cVar1S13S114P018N064P050N034(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='1' AND A(15)='1' )then
          cVar1S14S114P018N064P050P008(0) <='1';
          else
          cVar1S14S114P018N064P050P008(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='1' AND A(15)='1' )then
          cVar1S15S114P018N064P050P008(0) <='1';
          else
          cVar1S15S114P018N064P050P008(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S16S114P018N064P050N008(0) <='1';
          else
          cVar1S16S114P018N064P050N008(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S17S114P018N064P050N008(0) <='1';
          else
          cVar1S17S114P018N064P050N008(0) <='0';
          end if;
        if(A(10)='1' AND E( 1)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S18S114P018N064P050N008(0) <='1';
          else
          cVar1S18S114P018N064P050N008(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='0' )then
          cVar1S19S114N018P014P035P015(0) <='1';
          else
          cVar1S19S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='0' )then
          cVar1S20S114N018P014P035P015(0) <='1';
          else
          cVar1S20S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='0' )then
          cVar1S21S114N018P014P035P015(0) <='1';
          else
          cVar1S21S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='1' )then
          cVar1S22S114N018P014P035P015(0) <='1';
          else
          cVar1S22S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='1' )then
          cVar1S23S114N018P014P035P015(0) <='1';
          else
          cVar1S23S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='1' )then
          cVar1S24S114N018P014P035P015(0) <='1';
          else
          cVar1S24S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='0' AND A( 2)='1' )then
          cVar1S25S114N018P014P035P015(0) <='1';
          else
          cVar1S25S114N018P014P035P015(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='1' AND B(15)='0' )then
          cVar1S26S114N018P014P035P024(0) <='1';
          else
          cVar1S26S114N018P014P035P024(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='1' AND B(15)='0' )then
          cVar1S27S114N018P014P035P024(0) <='1';
          else
          cVar1S27S114N018P014P035P024(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND B( 1)='1' AND B(15)='0' )then
          cVar1S28S114N018P014P035P024(0) <='1';
          else
          cVar1S28S114N018P014P035P024(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='1' )then
          cVar1S29S114N018N014P010P030(0) <='1';
          else
          cVar1S29S114N018N014P010P030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='1' )then
          cVar1S30S114N018N014P010P030(0) <='1';
          else
          cVar1S30S114N018N014P010P030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='1' )then
          cVar1S31S114N018N014P010P030(0) <='1';
          else
          cVar1S31S114N018N014P010P030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='0' )then
          cVar1S32S114N018N014P010N030(0) <='1';
          else
          cVar1S32S114N018N014P010N030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='0' )then
          cVar1S33S114N018N014P010N030(0) <='1';
          else
          cVar1S33S114N018N014P010N030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='1' AND B(12)='0' )then
          cVar1S34S114N018N014P010N030(0) <='1';
          else
          cVar1S34S114N018N014P010N030(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='0' AND A( 4)='1' )then
          cVar1S35S114N018N014N010P011(0) <='1';
          else
          cVar1S35S114N018N014N010P011(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='0' AND A( 4)='1' )then
          cVar1S36S114N018N014N010P011(0) <='1';
          else
          cVar1S36S114N018N014N010P011(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='0' AND A( 4)='0' )then
          cVar1S37S114N018N014N010N011(0) <='1';
          else
          cVar1S37S114N018N014N010N011(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(14)='0' AND A( 4)='0' )then
          cVar1S38S114N018N014N010N011(0) <='1';
          else
          cVar1S38S114N018N014N010N011(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='0' )then
          cVar1S0S115P018P014P069P065(0) <='1';
          else
          cVar1S0S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='0' )then
          cVar1S1S115P018P014P069P065(0) <='1';
          else
          cVar1S1S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='0' )then
          cVar1S2S115P018P014P069P065(0) <='1';
          else
          cVar1S2S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='0' )then
          cVar1S3S115P018P014P069P065(0) <='1';
          else
          cVar1S3S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='1' )then
          cVar1S4S115P018P014P069P065(0) <='1';
          else
          cVar1S4S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='1' )then
          cVar1S5S115P018P014P069P065(0) <='1';
          else
          cVar1S5S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='1' AND E( 9)='1' )then
          cVar1S6S115P018P014P069P065(0) <='1';
          else
          cVar1S6S115P018P014P069P065(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S7S115P018P014N069P067(0) <='1';
          else
          cVar1S7S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S8S115P018P014N069P067(0) <='1';
          else
          cVar1S8S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S9S115P018P014N069P067(0) <='1';
          else
          cVar1S9S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='0' )then
          cVar1S10S115P018P014N069P067(0) <='1';
          else
          cVar1S10S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S11S115P018P014N069P067(0) <='1';
          else
          cVar1S11S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S12S115P018P014N069P067(0) <='1';
          else
          cVar1S12S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND E( 8)='0' AND D( 8)='1' )then
          cVar1S13S115P018P014N069P067(0) <='1';
          else
          cVar1S13S115P018P014N069P067(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='0' )then
          cVar1S14S115P018P014P007P064(0) <='1';
          else
          cVar1S14S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='0' )then
          cVar1S15S115P018P014P007P064(0) <='1';
          else
          cVar1S15S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='0' )then
          cVar1S16S115P018P014P007P064(0) <='1';
          else
          cVar1S16S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='1' )then
          cVar1S17S115P018P014P007P064(0) <='1';
          else
          cVar1S17S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='1' )then
          cVar1S18S115P018P014P007P064(0) <='1';
          else
          cVar1S18S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='0' AND E( 1)='1' )then
          cVar1S19S115P018P014P007P064(0) <='1';
          else
          cVar1S19S115P018P014P007P064(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='1' )then
          cVar1S20S115P018P014P007P037(0) <='1';
          else
          cVar1S20S115P018P014P007P037(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='1' )then
          cVar1S21S115P018P014P007P037(0) <='1';
          else
          cVar1S21S115P018P014P007P037(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='1' )then
          cVar1S22S115P018P014P007P037(0) <='1';
          else
          cVar1S22S115P018P014P007P037(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='0' )then
          cVar1S23S115P018P014P007N037(0) <='1';
          else
          cVar1S23S115P018P014P007N037(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='0' )then
          cVar1S24S115P018P014P007N037(0) <='1';
          else
          cVar1S24S115P018P014P007N037(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A( 6)='1' AND B( 0)='0' )then
          cVar1S25S115P018P014P007N037(0) <='1';
          else
          cVar1S25S115P018P014P007N037(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='0' AND D( 6)='0' )then
          cVar1S26S115P018P062P066P042(0) <='1';
          else
          cVar1S26S115P018P062P066P042(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='0' AND D( 6)='0' )then
          cVar1S27S115P018P062P066P042(0) <='1';
          else
          cVar1S27S115P018P062P066P042(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='0' AND D( 6)='0' )then
          cVar1S28S115P018P062P066P042(0) <='1';
          else
          cVar1S28S115P018P062P066P042(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='1' AND E( 0)='1' )then
          cVar1S29S115P018P062P066P068(0) <='1';
          else
          cVar1S29S115P018P062P066P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='1' AND E( 0)='1' )then
          cVar1S30S115P018P062P066P068(0) <='1';
          else
          cVar1S30S115P018P062P066P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='1' AND E( 0)='0' )then
          cVar1S31S115P018P062P066N068(0) <='1';
          else
          cVar1S31S115P018P062P066N068(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='1' AND D( 0)='1' AND E( 0)='0' )then
          cVar1S32S115P018P062P066N068(0) <='1';
          else
          cVar1S32S115P018P062P066N068(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='1' AND D(13)='1' )then
          cVar1S33S115P018N062P007P047(0) <='1';
          else
          cVar1S33S115P018N062P007P047(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='1' AND D(13)='1' )then
          cVar1S34S115P018N062P007P047(0) <='1';
          else
          cVar1S34S115P018N062P007P047(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='1' AND D(13)='0' )then
          cVar1S35S115P018N062P007N047(0) <='1';
          else
          cVar1S35S115P018N062P007N047(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='1' AND D(13)='0' )then
          cVar1S36S115P018N062P007N047(0) <='1';
          else
          cVar1S36S115P018N062P007N047(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='1' AND D(13)='0' )then
          cVar1S37S115P018N062P007N047(0) <='1';
          else
          cVar1S37S115P018N062P007N047(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='0' AND B(10)='1' )then
          cVar1S38S115P018N062N007P034(0) <='1';
          else
          cVar1S38S115P018N062N007P034(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='0' AND B(10)='1' )then
          cVar1S39S115P018N062N007P034(0) <='1';
          else
          cVar1S39S115P018N062N007P034(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='0' AND B(10)='1' )then
          cVar1S40S115P018N062N007P034(0) <='1';
          else
          cVar1S40S115P018N062N007P034(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='0' AND B(10)='0' )then
          cVar1S41S115P018N062N007N034(0) <='1';
          else
          cVar1S41S115P018N062N007N034(0) <='0';
          end if;
        if(A(10)='1' AND D( 1)='0' AND A( 6)='0' AND B(10)='0' )then
          cVar1S42S115P018N062N007N034(0) <='1';
          else
          cVar1S42S115P018N062N007N034(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='1' AND D(10)='0' )then
          cVar1S0S116P018P063P049P059(0) <='1';
          else
          cVar1S0S116P018P063P049P059(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='1' AND D(10)='0' )then
          cVar1S1S116P018P063P049P059(0) <='1';
          else
          cVar1S1S116P018P063P049P059(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='1' AND D(10)='0' )then
          cVar1S2S116P018P063P049P059(0) <='1';
          else
          cVar1S2S116P018P063P049P059(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='1' )then
          cVar1S3S116P018P063N049P066(0) <='1';
          else
          cVar1S3S116P018P063N049P066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='1' )then
          cVar1S4S116P018P063N049P066(0) <='1';
          else
          cVar1S4S116P018P063N049P066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='1' )then
          cVar1S5S116P018P063N049P066(0) <='1';
          else
          cVar1S5S116P018P063N049P066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='0' )then
          cVar1S6S116P018P063N049N066(0) <='1';
          else
          cVar1S6S116P018P063N049N066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='0' )then
          cVar1S7S116P018P063N049N066(0) <='1';
          else
          cVar1S7S116P018P063N049N066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='0' )then
          cVar1S8S116P018P063N049N066(0) <='1';
          else
          cVar1S8S116P018P063N049N066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='0' AND E(13)='0' AND D( 0)='0' )then
          cVar1S9S116P018P063N049N066(0) <='1';
          else
          cVar1S9S116P018P063N049N066(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='1' AND E( 3)='1' )then
          cVar1S10S116P018P063P031P056(0) <='1';
          else
          cVar1S10S116P018P063P031P056(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='1' AND E( 3)='1' )then
          cVar1S11S116P018P063P031P056(0) <='1';
          else
          cVar1S11S116P018P063P031P056(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='1' AND E( 3)='0' )then
          cVar1S12S116P018P063P031N056(0) <='1';
          else
          cVar1S12S116P018P063P031N056(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='1' )then
          cVar1S13S116P018P063N031P033(0) <='1';
          else
          cVar1S13S116P018P063N031P033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='1' )then
          cVar1S14S116P018P063N031P033(0) <='1';
          else
          cVar1S14S116P018P063N031P033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='1' )then
          cVar1S15S116P018P063N031P033(0) <='1';
          else
          cVar1S15S116P018P063N031P033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='1' )then
          cVar1S16S116P018P063N031P033(0) <='1';
          else
          cVar1S16S116P018P063N031P033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='0' )then
          cVar1S17S116P018P063N031N033(0) <='1';
          else
          cVar1S17S116P018P063N031N033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='0' )then
          cVar1S18S116P018P063N031N033(0) <='1';
          else
          cVar1S18S116P018P063N031N033(0) <='0';
          end if;
        if(A(10)='1' AND D( 9)='1' AND B( 3)='0' AND B( 2)='0' )then
          cVar1S19S116P018P063N031N033(0) <='1';
          else
          cVar1S19S116P018P063N031N033(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S20S116N018P069P064P019(0) <='1';
          else
          cVar1S20S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S21S116N018P069P064P019(0) <='1';
          else
          cVar1S21S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S22S116N018P069P064P019(0) <='1';
          else
          cVar1S22S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='0' )then
          cVar1S23S116N018P069P064P019(0) <='1';
          else
          cVar1S23S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S24S116N018P069P064P019(0) <='1';
          else
          cVar1S24S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S25S116N018P069P064P019(0) <='1';
          else
          cVar1S25S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='1' AND A( 0)='1' )then
          cVar1S26S116N018P069P064P019(0) <='1';
          else
          cVar1S26S116N018P069P064P019(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='0' AND E( 9)='0' )then
          cVar1S27S116N018P069N064P065(0) <='1';
          else
          cVar1S27S116N018P069N064P065(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='0' AND E( 9)='0' )then
          cVar1S28S116N018P069N064P065(0) <='1';
          else
          cVar1S28S116N018P069N064P065(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='0' AND E( 9)='0' )then
          cVar1S29S116N018P069N064P065(0) <='1';
          else
          cVar1S29S116N018P069N064P065(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='0' AND E( 9)='1' )then
          cVar1S30S116N018P069N064P065(0) <='1';
          else
          cVar1S30S116N018P069N064P065(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND E( 1)='0' AND E( 9)='1' )then
          cVar1S31S116N018P069N064P065(0) <='1';
          else
          cVar1S31S116N018P069N064P065(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='1' AND A(13)='1' )then
          cVar1S32S116N018N069P056P012(0) <='1';
          else
          cVar1S32S116N018N069P056P012(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='1' AND A(13)='1' )then
          cVar1S33S116N018N069P056P012(0) <='1';
          else
          cVar1S33S116N018N069P056P012(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='1' AND A(13)='1' )then
          cVar1S34S116N018N069P056P012(0) <='1';
          else
          cVar1S34S116N018N069P056P012(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='1' AND A(13)='0' )then
          cVar1S35S116N018N069P056N012(0) <='1';
          else
          cVar1S35S116N018N069P056N012(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='1' )then
          cVar1S36S116N018N069N056P013(0) <='1';
          else
          cVar1S36S116N018N069N056P013(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='1' )then
          cVar1S37S116N018N069N056P013(0) <='1';
          else
          cVar1S37S116N018N069N056P013(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='1' )then
          cVar1S38S116N018N069N056P013(0) <='1';
          else
          cVar1S38S116N018N069N056P013(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='1' )then
          cVar1S39S116N018N069N056P013(0) <='1';
          else
          cVar1S39S116N018N069N056P013(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='0' )then
          cVar1S40S116N018N069N056N013(0) <='1';
          else
          cVar1S40S116N018N069N056N013(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND E( 3)='0' AND A( 3)='0' )then
          cVar1S41S116N018N069N056N013(0) <='1';
          else
          cVar1S41S116N018N069N056N013(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='0' AND D( 8)='1' )then
          cVar1S0S117P066P069P063P067(0) <='1';
          else
          cVar1S0S117P066P069P063P067(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='0' AND D( 8)='1' )then
          cVar1S1S117P066P069P063P067(0) <='1';
          else
          cVar1S1S117P066P069P063P067(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='0' AND D( 8)='0' )then
          cVar1S2S117P066P069P063N067(0) <='1';
          else
          cVar1S2S117P066P069P063N067(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='0' AND D( 8)='0' )then
          cVar1S3S117P066P069P063N067(0) <='1';
          else
          cVar1S3S117P066P069P063N067(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='1' AND E(10)='0' )then
          cVar1S4S117P066P069P063P061(0) <='1';
          else
          cVar1S4S117P066P069P063P061(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='1' AND E(10)='0' )then
          cVar1S5S117P066P069P063P061(0) <='1';
          else
          cVar1S5S117P066P069P063P061(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='1' AND D( 9)='1' AND E(10)='1' )then
          cVar1S6S117P066P069P063P061(0) <='1';
          else
          cVar1S6S117P066P069P063P061(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='1' )then
          cVar1S7S117P066N069P068P047(0) <='1';
          else
          cVar1S7S117P066N069P068P047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='1' )then
          cVar1S8S117P066N069P068P047(0) <='1';
          else
          cVar1S8S117P066N069P068P047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='1' )then
          cVar1S9S117P066N069P068P047(0) <='1';
          else
          cVar1S9S117P066N069P068P047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='0' )then
          cVar1S10S117P066N069P068N047(0) <='1';
          else
          cVar1S10S117P066N069P068N047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='0' )then
          cVar1S11S117P066N069P068N047(0) <='1';
          else
          cVar1S11S117P066N069P068N047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='0' )then
          cVar1S12S117P066N069P068N047(0) <='1';
          else
          cVar1S12S117P066N069P068N047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='0' AND D(13)='0' )then
          cVar1S13S117P066N069P068N047(0) <='1';
          else
          cVar1S13S117P066N069P068N047(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='1' AND E( 1)='1' )then
          cVar1S14S117P066N069P068P064(0) <='1';
          else
          cVar1S14S117P066N069P068P064(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='1' AND E( 1)='1' )then
          cVar1S15S117P066N069P068P064(0) <='1';
          else
          cVar1S15S117P066N069P068P064(0) <='0';
          end if;
        if(D( 0)='0' AND E( 8)='0' AND E( 0)='1' AND E( 1)='0' )then
          cVar1S16S117P066N069P068N064(0) <='1';
          else
          cVar1S16S117P066N069P068N064(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='0' )then
          cVar1S17S117P066P018P006P047(0) <='1';
          else
          cVar1S17S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='0' )then
          cVar1S18S117P066P018P006P047(0) <='1';
          else
          cVar1S18S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='0' )then
          cVar1S19S117P066P018P006P047(0) <='1';
          else
          cVar1S19S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='0' )then
          cVar1S20S117P066P018P006P047(0) <='1';
          else
          cVar1S20S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='1' )then
          cVar1S21S117P066P018P006P047(0) <='1';
          else
          cVar1S21S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='0' AND D(13)='1' )then
          cVar1S22S117P066P018P006P047(0) <='1';
          else
          cVar1S22S117P066P018P006P047(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='1' AND B(15)='1' )then
          cVar1S23S117P066P018P006P024(0) <='1';
          else
          cVar1S23S117P066P018P006P024(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='1' AND B(15)='1' )then
          cVar1S24S117P066P018P006P024(0) <='1';
          else
          cVar1S24S117P066P018P006P024(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='1' AND B(15)='0' )then
          cVar1S25S117P066P018P006N024(0) <='1';
          else
          cVar1S25S117P066P018P006N024(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='0' AND A(16)='1' AND B(15)='0' )then
          cVar1S26S117P066P018P006N024(0) <='1';
          else
          cVar1S26S117P066P018P006N024(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='1' AND D(12)='1' )then
          cVar1S27S117P066P018P049P051nsss(0) <='1';
          else
          cVar1S27S117P066P018P049P051nsss(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='1' AND D(12)='0' )then
          cVar1S28S117P066P018P049N051(0) <='1';
          else
          cVar1S28S117P066P018P049N051(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='1' AND D(12)='0' )then
          cVar1S29S117P066P018P049N051(0) <='1';
          else
          cVar1S29S117P066P018P049N051(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='0' )then
          cVar1S30S117P066P018N049P067(0) <='1';
          else
          cVar1S30S117P066P018N049P067(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='0' )then
          cVar1S31S117P066P018N049P067(0) <='1';
          else
          cVar1S31S117P066P018N049P067(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='0' )then
          cVar1S32S117P066P018N049P067(0) <='1';
          else
          cVar1S32S117P066P018N049P067(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='1' )then
          cVar1S33S117P066P018N049P067(0) <='1';
          else
          cVar1S33S117P066P018N049P067(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='1' )then
          cVar1S34S117P066P018N049P067(0) <='1';
          else
          cVar1S34S117P066P018N049P067(0) <='0';
          end if;
        if(D( 0)='1' AND A(10)='1' AND E(13)='0' AND D( 8)='1' )then
          cVar1S35S117P066P018N049P067(0) <='1';
          else
          cVar1S35S117P066P018N049P067(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='0' AND E( 5)='1' )then
          cVar1S0S118P035P033P002P048(0) <='1';
          else
          cVar1S0S118P035P033P002P048(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S1S118P035P033P002N048(0) <='1';
          else
          cVar1S1S118P035P033P002N048(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S2S118P035P033P002N048(0) <='1';
          else
          cVar1S2S118P035P033P002N048(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='0' AND E( 5)='0' )then
          cVar1S3S118P035P033P002N048(0) <='1';
          else
          cVar1S3S118P035P033P002N048(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='1' AND A(10)='1' )then
          cVar1S4S118P035P033P002P018(0) <='1';
          else
          cVar1S4S118P035P033P002P018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='1' AND A(10)='0' )then
          cVar1S5S118P035P033P002N018(0) <='1';
          else
          cVar1S5S118P035P033P002N018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='1' AND A(18)='1' AND A(10)='0' )then
          cVar1S6S118P035P033P002N018(0) <='1';
          else
          cVar1S6S118P035P033P002N018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='0' )then
          cVar1S7S118P035N033P019P069(0) <='1';
          else
          cVar1S7S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='0' )then
          cVar1S8S118P035N033P019P069(0) <='1';
          else
          cVar1S8S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='0' )then
          cVar1S9S118P035N033P019P069(0) <='1';
          else
          cVar1S9S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='0' )then
          cVar1S10S118P035N033P019P069(0) <='1';
          else
          cVar1S10S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='1' )then
          cVar1S11S118P035N033P019P069(0) <='1';
          else
          cVar1S11S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='1' )then
          cVar1S12S118P035N033P019P069(0) <='1';
          else
          cVar1S12S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='0' AND E( 8)='1' )then
          cVar1S13S118P035N033P019P069(0) <='1';
          else
          cVar1S13S118P035N033P019P069(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='1' )then
          cVar1S14S118P035N033P019P018(0) <='1';
          else
          cVar1S14S118P035N033P019P018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='1' )then
          cVar1S15S118P035N033P019P018(0) <='1';
          else
          cVar1S15S118P035N033P019P018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='1' )then
          cVar1S16S118P035N033P019P018(0) <='1';
          else
          cVar1S16S118P035N033P019P018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar1S17S118P035N033P019N018(0) <='1';
          else
          cVar1S17S118P035N033P019N018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar1S18S118P035N033P019N018(0) <='1';
          else
          cVar1S18S118P035N033P019N018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar1S19S118P035N033P019N018(0) <='1';
          else
          cVar1S19S118P035N033P019N018(0) <='0';
          end if;
        if(B( 1)='0' AND B( 2)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar1S20S118P035N033P019N018(0) <='1';
          else
          cVar1S20S118P035N033P019N018(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='1' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S21S118P035P046P058P033(0) <='1';
          else
          cVar1S21S118P035P046P058P033(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='1' AND D( 2)='0' AND B( 2)='0' )then
          cVar1S22S118P035P046P058P033(0) <='1';
          else
          cVar1S22S118P035P046P058P033(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='0' )then
          cVar1S23S118P035N046P022P034(0) <='1';
          else
          cVar1S23S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='0' )then
          cVar1S24S118P035N046P022P034(0) <='1';
          else
          cVar1S24S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='0' )then
          cVar1S25S118P035N046P022P034(0) <='1';
          else
          cVar1S25S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='1' )then
          cVar1S26S118P035N046P022P034(0) <='1';
          else
          cVar1S26S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='1' )then
          cVar1S27S118P035N046P022P034(0) <='1';
          else
          cVar1S27S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='0' AND B(10)='1' )then
          cVar1S28S118P035N046P022P034(0) <='1';
          else
          cVar1S28S118P035N046P022P034(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='1' AND E( 9)='1' )then
          cVar1S29S118P035N046P022P065nsss(0) <='1';
          else
          cVar1S29S118P035N046P022P065nsss(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='1' AND E( 9)='0' )then
          cVar1S30S118P035N046P022N065(0) <='1';
          else
          cVar1S30S118P035N046P022N065(0) <='0';
          end if;
        if(B( 1)='1' AND D( 5)='0' AND B(16)='1' AND E( 9)='0' )then
          cVar1S31S118P035N046P022N065(0) <='1';
          else
          cVar1S31S118P035N046P022N065(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='0' AND B(11)='0' )then
          cVar1S0S119P065P027P010P032(0) <='1';
          else
          cVar1S0S119P065P027P010P032(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='0' AND B(11)='0' )then
          cVar1S1S119P065P027P010P032(0) <='1';
          else
          cVar1S1S119P065P027P010P032(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='0' AND B(11)='1' )then
          cVar1S2S119P065P027P010P032(0) <='1';
          else
          cVar1S2S119P065P027P010P032(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='1' AND B( 3)='0' )then
          cVar1S3S119P065P027P010P031(0) <='1';
          else
          cVar1S3S119P065P027P010P031(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='1' AND B( 3)='0' )then
          cVar1S4S119P065P027P010P031(0) <='1';
          else
          cVar1S4S119P065P027P010P031(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='1' AND A(14)='1' AND B( 3)='0' )then
          cVar1S5S119P065P027P010P031(0) <='1';
          else
          cVar1S5S119P065P027P010P031(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='1' )then
          cVar1S6S119P065N027P037P016(0) <='1';
          else
          cVar1S6S119P065N027P037P016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='1' )then
          cVar1S7S119P065N027P037P016(0) <='1';
          else
          cVar1S7S119P065N027P037P016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='1' )then
          cVar1S8S119P065N027P037P016(0) <='1';
          else
          cVar1S8S119P065N027P037P016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='0' )then
          cVar1S9S119P065N027P037N016(0) <='1';
          else
          cVar1S9S119P065N027P037N016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='0' )then
          cVar1S10S119P065N027P037N016(0) <='1';
          else
          cVar1S10S119P065N027P037N016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='0' AND A(11)='0' )then
          cVar1S11S119P065N027P037N016(0) <='1';
          else
          cVar1S11S119P065N027P037N016(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='1' )then
          cVar1S12S119P065N027P037P008(0) <='1';
          else
          cVar1S12S119P065N027P037P008(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='1' )then
          cVar1S13S119P065N027P037P008(0) <='1';
          else
          cVar1S13S119P065N027P037P008(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='1' )then
          cVar1S14S119P065N027P037P008(0) <='1';
          else
          cVar1S14S119P065N027P037P008(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='1' )then
          cVar1S15S119P065N027P037P008(0) <='1';
          else
          cVar1S15S119P065N027P037P008(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='0' )then
          cVar1S16S119P065N027P037N008(0) <='1';
          else
          cVar1S16S119P065N027P037N008(0) <='0';
          end if;
        if(E( 9)='0' AND B( 5)='0' AND B( 0)='1' AND A(15)='0' )then
          cVar1S17S119P065N027P037N008(0) <='1';
          else
          cVar1S17S119P065N027P037N008(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='0' AND E( 8)='0' )then
          cVar1S18S119P065P008P064P069(0) <='1';
          else
          cVar1S18S119P065P008P064P069(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='0' AND E( 8)='0' )then
          cVar1S19S119P065P008P064P069(0) <='1';
          else
          cVar1S19S119P065P008P064P069(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='0' AND E( 8)='0' )then
          cVar1S20S119P065P008P064P069(0) <='1';
          else
          cVar1S20S119P065P008P064P069(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='0' AND E( 8)='1' )then
          cVar1S21S119P065P008P064P069(0) <='1';
          else
          cVar1S21S119P065P008P064P069(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='0' AND E( 8)='1' )then
          cVar1S22S119P065P008P064P069(0) <='1';
          else
          cVar1S22S119P065P008P064P069(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='1' )then
          cVar1S23S119P065P008P064P014(0) <='1';
          else
          cVar1S23S119P065P008P064P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='1' )then
          cVar1S24S119P065P008P064P014(0) <='1';
          else
          cVar1S24S119P065P008P064P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='1' )then
          cVar1S25S119P065P008P064P014(0) <='1';
          else
          cVar1S25S119P065P008P064P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='0' )then
          cVar1S26S119P065P008P064N014(0) <='1';
          else
          cVar1S26S119P065P008P064N014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='0' )then
          cVar1S27S119P065P008P064N014(0) <='1';
          else
          cVar1S27S119P065P008P064N014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='0' )then
          cVar1S28S119P065P008P064N014(0) <='1';
          else
          cVar1S28S119P065P008P064N014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='0' AND E( 1)='1' AND A(12)='0' )then
          cVar1S29S119P065P008P064N014(0) <='1';
          else
          cVar1S29S119P065P008P064N014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='1' AND A(12)='0' )then
          cVar1S30S119P065P008P011P014(0) <='1';
          else
          cVar1S30S119P065P008P011P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='1' AND A(12)='0' )then
          cVar1S31S119P065P008P011P014(0) <='1';
          else
          cVar1S31S119P065P008P011P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='1' AND A(12)='1' )then
          cVar1S32S119P065P008P011P014(0) <='1';
          else
          cVar1S32S119P065P008P011P014(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='0' AND E( 3)='1' )then
          cVar1S33S119P065P008N011P056nsss(0) <='1';
          else
          cVar1S33S119P065P008N011P056nsss(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='0' AND E( 3)='0' )then
          cVar1S34S119P065P008N011N056(0) <='1';
          else
          cVar1S34S119P065P008N011N056(0) <='0';
          end if;
        if(E( 9)='1' AND A(15)='1' AND A( 4)='0' AND E( 3)='0' )then
          cVar1S35S119P065P008N011N056(0) <='1';
          else
          cVar1S35S119P065P008N011N056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='1' )then
          cVar1S0S120P037P001P032P018(0) <='1';
          else
          cVar1S0S120P037P001P032P018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='1' )then
          cVar1S1S120P037P001P032P018(0) <='1';
          else
          cVar1S1S120P037P001P032P018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='1' )then
          cVar1S2S120P037P001P032P018(0) <='1';
          else
          cVar1S2S120P037P001P032P018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='1' )then
          cVar1S3S120P037P001P032P018(0) <='1';
          else
          cVar1S3S120P037P001P032P018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='0' )then
          cVar1S4S120P037P001P032N018(0) <='1';
          else
          cVar1S4S120P037P001P032N018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='1' AND A(10)='0' )then
          cVar1S5S120P037P001P032N018(0) <='1';
          else
          cVar1S5S120P037P001P032N018(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='1' )then
          cVar1S6S120P037P001N032P056(0) <='1';
          else
          cVar1S6S120P037P001N032P056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='1' )then
          cVar1S7S120P037P001N032P056(0) <='1';
          else
          cVar1S7S120P037P001N032P056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='1' )then
          cVar1S8S120P037P001N032P056(0) <='1';
          else
          cVar1S8S120P037P001N032P056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='1' )then
          cVar1S9S120P037P001N032P056(0) <='1';
          else
          cVar1S9S120P037P001N032P056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='0' )then
          cVar1S10S120P037P001N032N056(0) <='1';
          else
          cVar1S10S120P037P001N032N056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='0' )then
          cVar1S11S120P037P001N032N056(0) <='1';
          else
          cVar1S11S120P037P001N032N056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='0' AND B(11)='0' AND E( 3)='0' )then
          cVar1S12S120P037P001N032N056(0) <='1';
          else
          cVar1S12S120P037P001N032N056(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='1' AND B( 9)='0' AND A( 0)='1' )then
          cVar1S13S120P037P001P036P019(0) <='1';
          else
          cVar1S13S120P037P001P036P019(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='1' AND B( 9)='0' AND A( 0)='1' )then
          cVar1S14S120P037P001P036P019(0) <='1';
          else
          cVar1S14S120P037P001P036P019(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='1' AND B( 9)='0' AND A( 0)='1' )then
          cVar1S15S120P037P001P036P019(0) <='1';
          else
          cVar1S15S120P037P001P036P019(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='1' AND B( 9)='0' AND A( 0)='0' )then
          cVar1S16S120P037P001P036N019(0) <='1';
          else
          cVar1S16S120P037P001P036N019(0) <='0';
          end if;
        if(B( 0)='1' AND A( 9)='1' AND B( 9)='1' AND A(15)='0' )then
          cVar1S17S120P037P001P036P008(0) <='1';
          else
          cVar1S17S120P037P001P036P008(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='1' )then
          cVar1S18S120N037P036P065P017(0) <='1';
          else
          cVar1S18S120N037P036P065P017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='1' )then
          cVar1S19S120N037P036P065P017(0) <='1';
          else
          cVar1S19S120N037P036P065P017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='1' )then
          cVar1S20S120N037P036P065P017(0) <='1';
          else
          cVar1S20S120N037P036P065P017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='0' )then
          cVar1S21S120N037P036P065N017(0) <='1';
          else
          cVar1S21S120N037P036P065N017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='0' )then
          cVar1S22S120N037P036P065N017(0) <='1';
          else
          cVar1S22S120N037P036P065N017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='0' AND A( 1)='0' )then
          cVar1S23S120N037P036P065N017(0) <='1';
          else
          cVar1S23S120N037P036P065N017(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='1' AND A(11)='0' )then
          cVar1S24S120N037P036P065P016(0) <='1';
          else
          cVar1S24S120N037P036P065P016(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='1' AND A(11)='0' )then
          cVar1S25S120N037P036P065P016(0) <='1';
          else
          cVar1S25S120N037P036P065P016(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='1' AND E( 9)='1' AND A(11)='1' )then
          cVar1S26S120N037P036P065P016(0) <='1';
          else
          cVar1S26S120N037P036P065P016(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='0' )then
          cVar1S27S120N037N036P034P050(0) <='1';
          else
          cVar1S27S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='0' )then
          cVar1S28S120N037N036P034P050(0) <='1';
          else
          cVar1S28S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='0' )then
          cVar1S29S120N037N036P034P050(0) <='1';
          else
          cVar1S29S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='0' )then
          cVar1S30S120N037N036P034P050(0) <='1';
          else
          cVar1S30S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='1' )then
          cVar1S31S120N037N036P034P050(0) <='1';
          else
          cVar1S31S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='1' AND D( 4)='1' )then
          cVar1S32S120N037N036P034P050(0) <='1';
          else
          cVar1S32S120N037N036P034P050(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='0' AND E( 9)='0' )then
          cVar1S33S120N037N036N034P065(0) <='1';
          else
          cVar1S33S120N037N036N034P065(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='0' AND E( 9)='0' )then
          cVar1S34S120N037N036N034P065(0) <='1';
          else
          cVar1S34S120N037N036N034P065(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='0' AND E( 9)='0' )then
          cVar1S35S120N037N036N034P065(0) <='1';
          else
          cVar1S35S120N037N036N034P065(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='0' AND E( 9)='1' )then
          cVar1S36S120N037N036N034P065(0) <='1';
          else
          cVar1S36S120N037N036N034P065(0) <='0';
          end if;
        if(B( 0)='0' AND B( 9)='0' AND B(10)='0' AND E( 9)='1' )then
          cVar1S37S120N037N036N034P065(0) <='1';
          else
          cVar1S37S120N037N036N034P065(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='0' AND A( 5)='1' )then
          cVar1S0S121P065P052P034P009(0) <='1';
          else
          cVar1S0S121P065P052P034P009(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='0' AND A( 5)='1' )then
          cVar1S1S121P065P052P034P009(0) <='1';
          else
          cVar1S1S121P065P052P034P009(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='0' AND A( 5)='1' )then
          cVar1S2S121P065P052P034P009(0) <='1';
          else
          cVar1S2S121P065P052P034P009(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='0' AND A( 5)='0' )then
          cVar1S3S121P065P052P034N009(0) <='1';
          else
          cVar1S3S121P065P052P034N009(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='0' AND A( 5)='0' )then
          cVar1S4S121P065P052P034N009(0) <='1';
          else
          cVar1S4S121P065P052P034N009(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='1' AND A( 4)='1' )then
          cVar1S5S121P065P052P034P011(0) <='1';
          else
          cVar1S5S121P065P052P034P011(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='1' AND B(10)='1' AND A( 4)='0' )then
          cVar1S6S121P065P052P034N011(0) <='1';
          else
          cVar1S6S121P065P052P034N011(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='1' )then
          cVar1S7S121P065N052P050P046(0) <='1';
          else
          cVar1S7S121P065N052P050P046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='1' )then
          cVar1S8S121P065N052P050P046(0) <='1';
          else
          cVar1S8S121P065N052P050P046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='1' )then
          cVar1S9S121P065N052P050P046(0) <='1';
          else
          cVar1S9S121P065N052P050P046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='0' )then
          cVar1S10S121P065N052P050N046(0) <='1';
          else
          cVar1S10S121P065N052P050N046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='0' )then
          cVar1S11S121P065N052P050N046(0) <='1';
          else
          cVar1S11S121P065N052P050N046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='0' AND D( 5)='0' )then
          cVar1S12S121P065N052P050N046(0) <='1';
          else
          cVar1S12S121P065N052P050N046(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='1' )then
          cVar1S13S121P065N052P050P060(0) <='1';
          else
          cVar1S13S121P065N052P050P060(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='1' )then
          cVar1S14S121P065N052P050P060(0) <='1';
          else
          cVar1S14S121P065N052P050P060(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='1' )then
          cVar1S15S121P065N052P050P060(0) <='1';
          else
          cVar1S15S121P065N052P050P060(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='0' )then
          cVar1S16S121P065N052P050N060(0) <='1';
          else
          cVar1S16S121P065N052P050N060(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='0' )then
          cVar1S17S121P065N052P050N060(0) <='1';
          else
          cVar1S17S121P065N052P050N060(0) <='0';
          end if;
        if(E( 9)='0' AND E( 4)='0' AND D( 4)='1' AND E( 2)='0' )then
          cVar1S18S121P065N052P050N060(0) <='1';
          else
          cVar1S18S121P065N052P050N060(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='0' AND B(12)='1' )then
          cVar1S19S121P065P036P024P030(0) <='1';
          else
          cVar1S19S121P065P036P024P030(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='0' AND B(12)='0' )then
          cVar1S20S121P065P036P024N030(0) <='1';
          else
          cVar1S20S121P065P036P024N030(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='0' AND B(12)='0' )then
          cVar1S21S121P065P036P024N030(0) <='1';
          else
          cVar1S21S121P065P036P024N030(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='0' AND B(12)='0' )then
          cVar1S22S121P065P036P024N030(0) <='1';
          else
          cVar1S22S121P065P036P024N030(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='0' AND B(12)='0' )then
          cVar1S23S121P065P036P024N030(0) <='1';
          else
          cVar1S23S121P065P036P024N030(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='1' AND B(15)='1' AND B(10)='0' )then
          cVar1S24S121P065P036P024P034(0) <='1';
          else
          cVar1S24S121P065P036P024P034(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='0' AND E(15)='0' )then
          cVar1S25S121P065N036P008P041(0) <='1';
          else
          cVar1S25S121P065N036P008P041(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='0' AND E(15)='0' )then
          cVar1S26S121P065N036P008P041(0) <='1';
          else
          cVar1S26S121P065N036P008P041(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='0' AND E(15)='0' )then
          cVar1S27S121P065N036P008P041(0) <='1';
          else
          cVar1S27S121P065N036P008P041(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='0' AND E(15)='1' )then
          cVar1S28S121P065N036P008P041(0) <='1';
          else
          cVar1S28S121P065N036P008P041(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='1' AND B( 0)='1' )then
          cVar1S29S121P065N036P008P037(0) <='1';
          else
          cVar1S29S121P065N036P008P037(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='1' AND B( 0)='1' )then
          cVar1S30S121P065N036P008P037(0) <='1';
          else
          cVar1S30S121P065N036P008P037(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='1' AND B( 0)='0' )then
          cVar1S31S121P065N036P008N037(0) <='1';
          else
          cVar1S31S121P065N036P008N037(0) <='0';
          end if;
        if(E( 9)='1' AND B( 9)='0' AND A(15)='1' AND B( 0)='0' )then
          cVar1S32S121P065N036P008N037(0) <='1';
          else
          cVar1S32S121P065N036P008N037(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='1' AND E( 3)='1' )then
          cVar1S0S122P052P009P056nsss(0) <='1';
          else
          cVar1S0S122P052P009P056nsss(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='1' AND E( 3)='0' AND A(14)='1' )then
          cVar1S1S122P052P009N056P010(0) <='1';
          else
          cVar1S1S122P052P009N056P010(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='1' AND E( 3)='0' AND A(14)='0' )then
          cVar1S2S122P052P009N056N010(0) <='1';
          else
          cVar1S2S122P052P009N056N010(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='1' AND E( 3)='0' AND A(14)='0' )then
          cVar1S3S122P052P009N056N010(0) <='1';
          else
          cVar1S3S122P052P009N056N010(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S4S122P052N009P056P046(0) <='1';
          else
          cVar1S4S122P052N009P056P046(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S5S122P052N009P056P046(0) <='1';
          else
          cVar1S5S122P052N009P056P046(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S6S122P052N009P056P046(0) <='1';
          else
          cVar1S6S122P052N009P056P046(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='0' AND D( 5)='1' )then
          cVar1S7S122P052N009P056P046(0) <='1';
          else
          cVar1S7S122P052N009P056P046(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='1' AND A( 2)='1' )then
          cVar1S8S122P052N009P056P015nsss(0) <='1';
          else
          cVar1S8S122P052N009P056P015nsss(0) <='0';
          end if;
        if(E( 4)='1' AND A( 5)='0' AND E( 3)='1' AND A( 2)='0' )then
          cVar1S9S122P052N009P056N015(0) <='1';
          else
          cVar1S9S122P052N009P056N015(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='0' AND D( 6)='0' )then
          cVar1S10S122N052P046P050P042(0) <='1';
          else
          cVar1S10S122N052P046P050P042(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='0' AND D( 6)='0' )then
          cVar1S11S122N052P046P050P042(0) <='1';
          else
          cVar1S11S122N052P046P050P042(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='0' AND D( 6)='0' )then
          cVar1S12S122N052P046P050P042(0) <='1';
          else
          cVar1S12S122N052P046P050P042(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='0' AND D( 6)='0' )then
          cVar1S13S122N052P046P050P042(0) <='1';
          else
          cVar1S13S122N052P046P050P042(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='0' AND D( 6)='1' )then
          cVar1S14S122N052P046P050P042(0) <='1';
          else
          cVar1S14S122N052P046P050P042(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='1' AND D( 4)='1' AND A(16)='1' )then
          cVar1S15S122N052P046P050P006nsss(0) <='1';
          else
          cVar1S15S122N052P046P050P006nsss(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='1' AND A(15)='0' )then
          cVar1S16S122N052N046P065P008(0) <='1';
          else
          cVar1S16S122N052N046P065P008(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='1' AND A(15)='0' )then
          cVar1S17S122N052N046P065P008(0) <='1';
          else
          cVar1S17S122N052N046P065P008(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='1' AND A(15)='0' )then
          cVar1S18S122N052N046P065P008(0) <='1';
          else
          cVar1S18S122N052N046P065P008(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='1' AND A(15)='1' )then
          cVar1S19S122N052N046P065P008(0) <='1';
          else
          cVar1S19S122N052N046P065P008(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='1' AND A(15)='1' )then
          cVar1S20S122N052N046P065P008(0) <='1';
          else
          cVar1S20S122N052N046P065P008(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='0' AND E(13)='1' )then
          cVar1S21S122N052N046N065P049(0) <='1';
          else
          cVar1S21S122N052N046N065P049(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='0' AND E(13)='1' )then
          cVar1S22S122N052N046N065P049(0) <='1';
          else
          cVar1S22S122N052N046N065P049(0) <='0';
          end if;
        if(E( 4)='0' AND D( 5)='0' AND E( 9)='0' AND E(13)='0' )then
          cVar1S23S122N052N046N065N049(0) <='1';
          else
          cVar1S23S122N052N046N065N049(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='0' )then
          cVar1S0S123P017P036P016P021(0) <='1';
          else
          cVar1S0S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='0' )then
          cVar1S1S123P017P036P016P021(0) <='1';
          else
          cVar1S1S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='0' )then
          cVar1S2S123P017P036P016P021(0) <='1';
          else
          cVar1S2S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='0' )then
          cVar1S3S123P017P036P016P021(0) <='1';
          else
          cVar1S3S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='1' )then
          cVar1S4S123P017P036P016P021(0) <='1';
          else
          cVar1S4S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='1' AND B( 8)='1' )then
          cVar1S5S123P017P036P016P021(0) <='1';
          else
          cVar1S5S123P017P036P016P021(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='0' )then
          cVar1S6S123P017P036N016P034(0) <='1';
          else
          cVar1S6S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='0' )then
          cVar1S7S123P017P036N016P034(0) <='1';
          else
          cVar1S7S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='0' )then
          cVar1S8S123P017P036N016P034(0) <='1';
          else
          cVar1S8S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='1' )then
          cVar1S9S123P017P036N016P034(0) <='1';
          else
          cVar1S9S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='1' )then
          cVar1S10S123P017P036N016P034(0) <='1';
          else
          cVar1S10S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='0' AND A(11)='0' AND B(10)='1' )then
          cVar1S11S123P017P036N016P034(0) <='1';
          else
          cVar1S11S123P017P036N016P034(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='1' AND E( 4)='0' )then
          cVar1S12S123P017P036P056P052(0) <='1';
          else
          cVar1S12S123P017P036P056P052(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='1' AND E( 4)='0' )then
          cVar1S13S123P017P036P056P052(0) <='1';
          else
          cVar1S13S123P017P036P056P052(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='1' AND E( 4)='0' )then
          cVar1S14S123P017P036P056P052(0) <='1';
          else
          cVar1S14S123P017P036P056P052(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='0' AND E( 9)='1' )then
          cVar1S15S123P017P036N056P065(0) <='1';
          else
          cVar1S15S123P017P036N056P065(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='0' AND E( 9)='1' )then
          cVar1S16S123P017P036N056P065(0) <='1';
          else
          cVar1S16S123P017P036N056P065(0) <='0';
          end if;
        if(A( 1)='0' AND B( 9)='1' AND E( 3)='0' AND E( 9)='0' )then
          cVar1S17S123P017P036N056N065(0) <='1';
          else
          cVar1S17S123P017P036N056N065(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='0' )then
          cVar1S18S123P017P036P065P019(0) <='1';
          else
          cVar1S18S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='0' )then
          cVar1S19S123P017P036P065P019(0) <='1';
          else
          cVar1S19S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='0' )then
          cVar1S20S123P017P036P065P019(0) <='1';
          else
          cVar1S20S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='0' )then
          cVar1S21S123P017P036P065P019(0) <='1';
          else
          cVar1S21S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='1' )then
          cVar1S22S123P017P036P065P019(0) <='1';
          else
          cVar1S22S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='1' )then
          cVar1S23S123P017P036P065P019(0) <='1';
          else
          cVar1S23S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='1' )then
          cVar1S24S123P017P036P065P019(0) <='1';
          else
          cVar1S24S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='0' AND A( 0)='1' )then
          cVar1S25S123P017P036P065P019(0) <='1';
          else
          cVar1S25S123P017P036P065P019(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='1' AND D( 9)='1' )then
          cVar1S26S123P017P036P065P063(0) <='1';
          else
          cVar1S26S123P017P036P065P063(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='1' AND D( 9)='1' )then
          cVar1S27S123P017P036P065P063(0) <='1';
          else
          cVar1S27S123P017P036P065P063(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='1' AND D( 9)='1' )then
          cVar1S28S123P017P036P065P063(0) <='1';
          else
          cVar1S28S123P017P036P065P063(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='1' AND D( 9)='1' )then
          cVar1S29S123P017P036P065P063(0) <='1';
          else
          cVar1S29S123P017P036P065P063(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='1' AND E( 9)='1' AND D( 9)='0' )then
          cVar1S30S123P017P036P065N063(0) <='1';
          else
          cVar1S30S123P017P036P065N063(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='1' )then
          cVar1S31S123P017N036P060P069(0) <='1';
          else
          cVar1S31S123P017N036P060P069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='1' )then
          cVar1S32S123P017N036P060P069(0) <='1';
          else
          cVar1S32S123P017N036P060P069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='1' )then
          cVar1S33S123P017N036P060P069(0) <='1';
          else
          cVar1S33S123P017N036P060P069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='0' )then
          cVar1S34S123P017N036P060N069(0) <='1';
          else
          cVar1S34S123P017N036P060N069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='0' )then
          cVar1S35S123P017N036P060N069(0) <='1';
          else
          cVar1S35S123P017N036P060N069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='1' AND E( 8)='0' )then
          cVar1S36S123P017N036P060N069(0) <='1';
          else
          cVar1S36S123P017N036P060N069(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='1' )then
          cVar1S37S123P017N036N060P037(0) <='1';
          else
          cVar1S37S123P017N036N060P037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='1' )then
          cVar1S38S123P017N036N060P037(0) <='1';
          else
          cVar1S38S123P017N036N060P037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='1' )then
          cVar1S39S123P017N036N060P037(0) <='1';
          else
          cVar1S39S123P017N036N060P037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='1' )then
          cVar1S40S123P017N036N060P037(0) <='1';
          else
          cVar1S40S123P017N036N060P037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='0' )then
          cVar1S41S123P017N036N060N037(0) <='1';
          else
          cVar1S41S123P017N036N060N037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='0' )then
          cVar1S42S123P017N036N060N037(0) <='1';
          else
          cVar1S42S123P017N036N060N037(0) <='0';
          end if;
        if(A( 1)='1' AND B( 9)='0' AND E( 2)='0' AND B( 0)='0' )then
          cVar1S43S123P017N036N060N037(0) <='1';
          else
          cVar1S43S123P017N036N060N037(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='0' AND A( 0)='0' )then
          cVar1S0S124P036P065P032P019(0) <='1';
          else
          cVar1S0S124P036P065P032P019(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='0' AND A( 0)='0' )then
          cVar1S1S124P036P065P032P019(0) <='1';
          else
          cVar1S1S124P036P065P032P019(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='0' AND A( 0)='0' )then
          cVar1S2S124P036P065P032P019(0) <='1';
          else
          cVar1S2S124P036P065P032P019(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='0' AND A( 0)='1' )then
          cVar1S3S124P036P065P032P019(0) <='1';
          else
          cVar1S3S124P036P065P032P019(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='0' AND A( 0)='1' )then
          cVar1S4S124P036P065P032P019(0) <='1';
          else
          cVar1S4S124P036P065P032P019(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='1' AND D(11)='0' )then
          cVar1S5S124P036P065P032P055(0) <='1';
          else
          cVar1S5S124P036P065P032P055(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='0' AND B(11)='1' AND D(11)='0' )then
          cVar1S6S124P036P065P032P055(0) <='1';
          else
          cVar1S6S124P036P065P032P055(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='1' )then
          cVar1S7S124P036P065P024P063(0) <='1';
          else
          cVar1S7S124P036P065P024P063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='1' )then
          cVar1S8S124P036P065P024P063(0) <='1';
          else
          cVar1S8S124P036P065P024P063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='1' )then
          cVar1S9S124P036P065P024P063(0) <='1';
          else
          cVar1S9S124P036P065P024P063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='1' )then
          cVar1S10S124P036P065P024P063(0) <='1';
          else
          cVar1S10S124P036P065P024P063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='0' )then
          cVar1S11S124P036P065P024N063(0) <='1';
          else
          cVar1S11S124P036P065P024N063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='0' )then
          cVar1S12S124P036P065P024N063(0) <='1';
          else
          cVar1S12S124P036P065P024N063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='0' AND D( 9)='0' )then
          cVar1S13S124P036P065P024N063(0) <='1';
          else
          cVar1S13S124P036P065P024N063(0) <='0';
          end if;
        if(B( 9)='1' AND E( 9)='1' AND B(15)='1' AND B(10)='0' )then
          cVar1S14S124P036P065P024P034(0) <='1';
          else
          cVar1S14S124P036P065P024P034(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='1' AND D(14)='1' )then
          cVar1S15S124N036P017P034P043nsss(0) <='1';
          else
          cVar1S15S124N036P017P034P043nsss(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='1' AND D(14)='0' )then
          cVar1S16S124N036P017P034N043(0) <='1';
          else
          cVar1S16S124N036P017P034N043(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='1' AND D(14)='0' )then
          cVar1S17S124N036P017P034N043(0) <='1';
          else
          cVar1S17S124N036P017P034N043(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='1' AND D(14)='0' )then
          cVar1S18S124N036P017P034N043(0) <='1';
          else
          cVar1S18S124N036P017P034N043(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='1' AND D(14)='0' )then
          cVar1S19S124N036P017P034N043(0) <='1';
          else
          cVar1S19S124N036P017P034N043(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='0' AND A(18)='0' )then
          cVar1S20S124N036P017N034P002(0) <='1';
          else
          cVar1S20S124N036P017N034P002(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='0' AND A(18)='0' )then
          cVar1S21S124N036P017N034P002(0) <='1';
          else
          cVar1S21S124N036P017N034P002(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='0' AND A(18)='1' )then
          cVar1S22S124N036P017N034P002(0) <='1';
          else
          cVar1S22S124N036P017N034P002(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='1' AND B(10)='0' AND A(18)='1' )then
          cVar1S23S124N036P017N034P002(0) <='1';
          else
          cVar1S23S124N036P017N034P002(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='1' AND B( 3)='0' )then
          cVar1S24S124N036N017P032P031(0) <='1';
          else
          cVar1S24S124N036N017P032P031(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='1' AND B( 3)='0' )then
          cVar1S25S124N036N017P032P031(0) <='1';
          else
          cVar1S25S124N036N017P032P031(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='1' AND B( 3)='1' )then
          cVar1S26S124N036N017P032P031(0) <='1';
          else
          cVar1S26S124N036N017P032P031(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='1' AND B( 3)='1' )then
          cVar1S27S124N036N017P032P031(0) <='1';
          else
          cVar1S27S124N036N017P032P031(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='0' AND D( 5)='1' )then
          cVar1S28S124N036N017N032P046(0) <='1';
          else
          cVar1S28S124N036N017N032P046(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='0' AND D( 5)='1' )then
          cVar1S29S124N036N017N032P046(0) <='1';
          else
          cVar1S29S124N036N017N032P046(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='0' AND D( 5)='0' )then
          cVar1S30S124N036N017N032N046(0) <='1';
          else
          cVar1S30S124N036N017N032N046(0) <='0';
          end if;
        if(B( 9)='0' AND A( 1)='0' AND B(11)='0' AND D( 5)='0' )then
          cVar1S31S124N036N017N032N046(0) <='1';
          else
          cVar1S31S124N036N017N032N046(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='0' AND B(16)='0' )then
          cVar1S0S125P032P064P050P022(0) <='1';
          else
          cVar1S0S125P032P064P050P022(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='0' AND B(16)='0' )then
          cVar1S1S125P032P064P050P022(0) <='1';
          else
          cVar1S1S125P032P064P050P022(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='0' AND B(16)='0' )then
          cVar1S2S125P032P064P050P022(0) <='1';
          else
          cVar1S2S125P032P064P050P022(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='0' AND B(16)='1' )then
          cVar1S3S125P032P064P050P022(0) <='1';
          else
          cVar1S3S125P032P064P050P022(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='0' AND B(16)='1' )then
          cVar1S4S125P032P064P050P022(0) <='1';
          else
          cVar1S4S125P032P064P050P022(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='1' AND B( 5)='1' )then
          cVar1S5S125P032P064P050P027(0) <='1';
          else
          cVar1S5S125P032P064P050P027(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S6S125P032P064P050N027(0) <='1';
          else
          cVar1S6S125P032P064P050N027(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S7S125P032P064P050N027(0) <='1';
          else
          cVar1S7S125P032P064P050N027(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='1' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S8S125P032P064P050N027(0) <='1';
          else
          cVar1S8S125P032P064P050N027(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='1' )then
          cVar1S9S125P032N064P037P068(0) <='1';
          else
          cVar1S9S125P032N064P037P068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='1' )then
          cVar1S10S125P032N064P037P068(0) <='1';
          else
          cVar1S10S125P032N064P037P068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='1' )then
          cVar1S11S125P032N064P037P068(0) <='1';
          else
          cVar1S11S125P032N064P037P068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='0' )then
          cVar1S12S125P032N064P037N068(0) <='1';
          else
          cVar1S12S125P032N064P037N068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='0' )then
          cVar1S13S125P032N064P037N068(0) <='1';
          else
          cVar1S13S125P032N064P037N068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='0' AND E( 0)='0' )then
          cVar1S14S125P032N064P037N068(0) <='1';
          else
          cVar1S14S125P032N064P037N068(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='1' )then
          cVar1S15S125P032N064P037P056(0) <='1';
          else
          cVar1S15S125P032N064P037P056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='1' )then
          cVar1S16S125P032N064P037P056(0) <='1';
          else
          cVar1S16S125P032N064P037P056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='1' )then
          cVar1S17S125P032N064P037P056(0) <='1';
          else
          cVar1S17S125P032N064P037P056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='1' )then
          cVar1S18S125P032N064P037P056(0) <='1';
          else
          cVar1S18S125P032N064P037P056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='0' )then
          cVar1S19S125P032N064P037N056(0) <='1';
          else
          cVar1S19S125P032N064P037N056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='0' )then
          cVar1S20S125P032N064P037N056(0) <='1';
          else
          cVar1S20S125P032N064P037N056(0) <='0';
          end if;
        if(B(11)='0' AND E( 1)='0' AND B( 0)='1' AND E( 3)='0' )then
          cVar1S21S125P032N064P037N056(0) <='1';
          else
          cVar1S21S125P032N064P037N056(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='1' AND A(11)='0' )then
          cVar1S22S125P032P037P063P016(0) <='1';
          else
          cVar1S22S125P032P037P063P016(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='1' AND A(11)='0' )then
          cVar1S23S125P032P037P063P016(0) <='1';
          else
          cVar1S23S125P032P037P063P016(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='1' AND A(11)='1' )then
          cVar1S24S125P032P037P063P016(0) <='1';
          else
          cVar1S24S125P032P037P063P016(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='0' AND A(13)='1' )then
          cVar1S25S125P032P037N063P012(0) <='1';
          else
          cVar1S25S125P032P037N063P012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='0' AND A(13)='1' )then
          cVar1S26S125P032P037N063P012(0) <='1';
          else
          cVar1S26S125P032P037N063P012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='0' AND A(13)='0' )then
          cVar1S27S125P032P037N063N012(0) <='1';
          else
          cVar1S27S125P032P037N063N012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='1' AND D( 9)='0' AND A(13)='0' )then
          cVar1S28S125P032P037N063N012(0) <='1';
          else
          cVar1S28S125P032P037N063N012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='0' AND E( 0)='1' )then
          cVar1S29S125P032N037P031P068(0) <='1';
          else
          cVar1S29S125P032N037P031P068(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='0' AND E( 0)='1' )then
          cVar1S30S125P032N037P031P068(0) <='1';
          else
          cVar1S30S125P032N037P031P068(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='0' AND E( 0)='1' )then
          cVar1S31S125P032N037P031P068(0) <='1';
          else
          cVar1S31S125P032N037P031P068(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='0' AND E( 0)='0' )then
          cVar1S32S125P032N037P031N068(0) <='1';
          else
          cVar1S32S125P032N037P031N068(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='0' AND E( 0)='0' )then
          cVar1S33S125P032N037P031N068(0) <='1';
          else
          cVar1S33S125P032N037P031N068(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='1' AND A(13)='0' )then
          cVar1S34S125P032N037P031P012(0) <='1';
          else
          cVar1S34S125P032N037P031P012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='1' AND A(13)='0' )then
          cVar1S35S125P032N037P031P012(0) <='1';
          else
          cVar1S35S125P032N037P031P012(0) <='0';
          end if;
        if(B(11)='1' AND B( 0)='0' AND B( 3)='1' AND A(13)='1' )then
          cVar1S36S125P032N037P031P012(0) <='1';
          else
          cVar1S36S125P032N037P031P012(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='1' AND E( 1)='1' )then
          cVar1S0S126P069P018P026P064nsss(0) <='1';
          else
          cVar1S0S126P069P018P026P064nsss(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='1' AND E( 1)='0' )then
          cVar1S1S126P069P018P026N064(0) <='1';
          else
          cVar1S1S126P069P018P026N064(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='1' AND E( 1)='0' )then
          cVar1S2S126P069P018P026N064(0) <='1';
          else
          cVar1S2S126P069P018P026N064(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='0' AND B( 3)='1' )then
          cVar1S3S126P069P018N026P031(0) <='1';
          else
          cVar1S3S126P069P018N026P031(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='0' AND B( 3)='0' )then
          cVar1S4S126P069P018N026N031(0) <='1';
          else
          cVar1S4S126P069P018N026N031(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='0' AND B( 3)='0' )then
          cVar1S5S126P069P018N026N031(0) <='1';
          else
          cVar1S5S126P069P018N026N031(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='0' AND B( 3)='0' )then
          cVar1S6S126P069P018N026N031(0) <='1';
          else
          cVar1S6S126P069P018N026N031(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='0' AND B(14)='0' AND B( 3)='0' )then
          cVar1S7S126P069P018N026N031(0) <='1';
          else
          cVar1S7S126P069P018N026N031(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='0' AND D( 8)='1' )then
          cVar1S8S126P069P018P068P067(0) <='1';
          else
          cVar1S8S126P069P018P068P067(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='0' AND D( 8)='1' )then
          cVar1S9S126P069P018P068P067(0) <='1';
          else
          cVar1S9S126P069P018P068P067(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='0' AND D( 8)='1' )then
          cVar1S10S126P069P018P068P067(0) <='1';
          else
          cVar1S10S126P069P018P068P067(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='0' AND D( 8)='0' )then
          cVar1S11S126P069P018P068N067(0) <='1';
          else
          cVar1S11S126P069P018P068N067(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='0' AND D( 8)='0' )then
          cVar1S12S126P069P018P068N067(0) <='1';
          else
          cVar1S12S126P069P018P068N067(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='1' AND E( 7)='1' )then
          cVar1S13S126P069P018P068P040nsss(0) <='1';
          else
          cVar1S13S126P069P018P068P040nsss(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='1' AND E( 7)='0' )then
          cVar1S14S126P069P018P068N040(0) <='1';
          else
          cVar1S14S126P069P018P068N040(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='1' AND E( 7)='0' )then
          cVar1S15S126P069P018P068N040(0) <='1';
          else
          cVar1S15S126P069P018P068N040(0) <='0';
          end if;
        if(E( 8)='1' AND A(10)='1' AND E( 0)='1' AND E( 7)='0' )then
          cVar1S16S126P069P018P068N040(0) <='1';
          else
          cVar1S16S126P069P018P068N040(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='1' AND B(11)='0' )then
          cVar1S17S126N069P018P049P032(0) <='1';
          else
          cVar1S17S126N069P018P049P032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='1' AND B(11)='0' )then
          cVar1S18S126N069P018P049P032(0) <='1';
          else
          cVar1S18S126N069P018P049P032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='1' AND B(11)='0' )then
          cVar1S19S126N069P018P049P032(0) <='1';
          else
          cVar1S19S126N069P018P049P032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='0' AND B(11)='1' )then
          cVar1S20S126N069P018N049P032(0) <='1';
          else
          cVar1S20S126N069P018N049P032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='0' AND B(11)='0' )then
          cVar1S21S126N069P018N049N032(0) <='1';
          else
          cVar1S21S126N069P018N049N032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='0' AND B(11)='0' )then
          cVar1S22S126N069P018N049N032(0) <='1';
          else
          cVar1S22S126N069P018N049N032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND E(13)='0' AND B(11)='0' )then
          cVar1S23S126N069P018N049N032(0) <='1';
          else
          cVar1S23S126N069P018N049N032(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='0' )then
          cVar1S24S126N069N018P066P064(0) <='1';
          else
          cVar1S24S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='0' )then
          cVar1S25S126N069N018P066P064(0) <='1';
          else
          cVar1S25S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='0' )then
          cVar1S26S126N069N018P066P064(0) <='1';
          else
          cVar1S26S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='1' )then
          cVar1S27S126N069N018P066P064(0) <='1';
          else
          cVar1S27S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='1' )then
          cVar1S28S126N069N018P066P064(0) <='1';
          else
          cVar1S28S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='1' )then
          cVar1S29S126N069N018P066P064(0) <='1';
          else
          cVar1S29S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='0' AND E( 1)='1' )then
          cVar1S30S126N069N018P066P064(0) <='1';
          else
          cVar1S30S126N069N018P066P064(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='0' )then
          cVar1S31S126N069N018P066P006(0) <='1';
          else
          cVar1S31S126N069N018P066P006(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='0' )then
          cVar1S32S126N069N018P066P006(0) <='1';
          else
          cVar1S32S126N069N018P066P006(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='1' )then
          cVar1S33S126N069N018P066P006(0) <='1';
          else
          cVar1S33S126N069N018P066P006(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='1' )then
          cVar1S34S126N069N018P066P006(0) <='1';
          else
          cVar1S34S126N069N018P066P006(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='1' )then
          cVar1S35S126N069N018P066P006(0) <='1';
          else
          cVar1S35S126N069N018P066P006(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND D( 0)='1' AND A(16)='1' )then
          cVar1S36S126N069N018P066P006(0) <='1';
          else
          cVar1S36S126N069N018P066P006(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='0' )then
          cVar1S0S127P064P069P034P016(0) <='1';
          else
          cVar1S0S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='0' )then
          cVar1S1S127P064P069P034P016(0) <='1';
          else
          cVar1S1S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='1' )then
          cVar1S2S127P064P069P034P016(0) <='1';
          else
          cVar1S2S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='1' )then
          cVar1S3S127P064P069P034P016(0) <='1';
          else
          cVar1S3S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='1' )then
          cVar1S4S127P064P069P034P016(0) <='1';
          else
          cVar1S4S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='0' AND A(11)='1' )then
          cVar1S5S127P064P069P034P016(0) <='1';
          else
          cVar1S5S127P064P069P034P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='1' AND A(15)='0' )then
          cVar1S6S127P064P069P034P008(0) <='1';
          else
          cVar1S6S127P064P069P034P008(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='1' AND A(15)='0' )then
          cVar1S7S127P064P069P034P008(0) <='1';
          else
          cVar1S7S127P064P069P034P008(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='1' AND A(15)='0' )then
          cVar1S8S127P064P069P034P008(0) <='1';
          else
          cVar1S8S127P064P069P034P008(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='1' AND A(15)='1' )then
          cVar1S9S127P064P069P034P008(0) <='1';
          else
          cVar1S9S127P064P069P034P008(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='0' AND B(10)='1' AND A(15)='1' )then
          cVar1S10S127P064P069P034P008(0) <='1';
          else
          cVar1S10S127P064P069P034P008(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='1' AND A(11)='0' )then
          cVar1S11S127P064P069P037P016(0) <='1';
          else
          cVar1S11S127P064P069P037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='1' AND A(11)='0' )then
          cVar1S12S127P064P069P037P016(0) <='1';
          else
          cVar1S12S127P064P069P037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='1' AND A(11)='0' )then
          cVar1S13S127P064P069P037P016(0) <='1';
          else
          cVar1S13S127P064P069P037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='1' AND A(11)='1' )then
          cVar1S14S127P064P069P037P016(0) <='1';
          else
          cVar1S14S127P064P069P037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='1' )then
          cVar1S15S127P064P069N037P016(0) <='1';
          else
          cVar1S15S127P064P069N037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='1' )then
          cVar1S16S127P064P069N037P016(0) <='1';
          else
          cVar1S16S127P064P069N037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='1' )then
          cVar1S17S127P064P069N037P016(0) <='1';
          else
          cVar1S17S127P064P069N037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='1' )then
          cVar1S18S127P064P069N037P016(0) <='1';
          else
          cVar1S18S127P064P069N037P016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='0' )then
          cVar1S19S127P064P069N037N016(0) <='1';
          else
          cVar1S19S127P064P069N037N016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='0' )then
          cVar1S20S127P064P069N037N016(0) <='1';
          else
          cVar1S20S127P064P069N037N016(0) <='0';
          end if;
        if(E( 1)='0' AND E( 8)='1' AND B( 0)='0' AND A(11)='0' )then
          cVar1S21S127P064P069N037N016(0) <='1';
          else
          cVar1S21S127P064P069N037N016(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='0' )then
          cVar1S22S127P064P018P054P035(0) <='1';
          else
          cVar1S22S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='0' )then
          cVar1S23S127P064P018P054P035(0) <='1';
          else
          cVar1S23S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='0' )then
          cVar1S24S127P064P018P054P035(0) <='1';
          else
          cVar1S24S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='1' )then
          cVar1S25S127P064P018P054P035(0) <='1';
          else
          cVar1S25S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='1' )then
          cVar1S26S127P064P018P054P035(0) <='1';
          else
          cVar1S26S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='1' )then
          cVar1S27S127P064P018P054P035(0) <='1';
          else
          cVar1S27S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='0' AND B( 1)='1' )then
          cVar1S28S127P064P018P054P035(0) <='1';
          else
          cVar1S28S127P064P018P054P035(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='1' AND E( 9)='1' )then
          cVar1S29S127P064P018P054P065nsss(0) <='1';
          else
          cVar1S29S127P064P018P054P065nsss(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='1' AND E( 9)='0' )then
          cVar1S30S127P064P018P054N065(0) <='1';
          else
          cVar1S30S127P064P018P054N065(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='1' AND D( 3)='1' AND E( 9)='0' )then
          cVar1S31S127P064P018P054N065(0) <='1';
          else
          cVar1S31S127P064P018P054N065(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='0' AND E( 5)='0' )then
          cVar1S32S127P064N018P050P048(0) <='1';
          else
          cVar1S32S127P064N018P050P048(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='0' AND E( 5)='0' )then
          cVar1S33S127P064N018P050P048(0) <='1';
          else
          cVar1S33S127P064N018P050P048(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='0' AND E( 5)='0' )then
          cVar1S34S127P064N018P050P048(0) <='1';
          else
          cVar1S34S127P064N018P050P048(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='0' AND E( 5)='1' )then
          cVar1S35S127P064N018P050P048(0) <='1';
          else
          cVar1S35S127P064N018P050P048(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='1' AND B( 5)='1' )then
          cVar1S36S127P064N018P050P027nsss(0) <='1';
          else
          cVar1S36S127P064N018P050P027nsss(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S37S127P064N018P050N027(0) <='1';
          else
          cVar1S37S127P064N018P050N027(0) <='0';
          end if;
        if(E( 1)='1' AND A(10)='0' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S38S127P064N018P050N027(0) <='1';
          else
          cVar1S38S127P064N018P050N027(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV2 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar1S0S0P069P019P067P064(0)='1' AND  D( 1)='1' AND A( 4)='0' )then
          cVar2S0S0P062P011nsss(0) <='1';
          else
          cVar2S0S0P062P011nsss(0) <='0';
          end if;
        if(cVar1S1S0P069P019P067P064(0)='1' AND  D( 1)='1' AND A( 4)='1' AND A(12)='0' )then
          cVar2S1S0P062P011P014nsss(0) <='1';
          else
          cVar2S1S0P062P011P014nsss(0) <='0';
          end if;
        if(cVar1S2S0P069P019P067P064(0)='1' AND  D( 1)='0' AND D( 0)='1' )then
          cVar2S2S0N062P066nsss(0) <='1';
          else
          cVar2S2S0N062P066nsss(0) <='0';
          end if;
        if(cVar1S3S0P069P019P067N064(0)='1' AND  D( 2)='1' AND B( 2)='1' )then
          cVar2S3S0P058P033nsss(0) <='1';
          else
          cVar2S3S0P058P033nsss(0) <='0';
          end if;
        if(cVar1S4S0P069P019P067N064(0)='1' AND  D( 2)='1' AND B( 2)='0' AND A( 3)='0' )then
          cVar2S4S0P058N033P013nsss(0) <='1';
          else
          cVar2S4S0P058N033P013nsss(0) <='0';
          end if;
        if(cVar1S5S0P069P019P067N064(0)='1' AND  D( 2)='0' AND E( 0)='1' AND D( 0)='1' )then
          cVar2S5S0N058P068P066nsss(0) <='1';
          else
          cVar2S5S0N058P068P066nsss(0) <='0';
          end if;
        if(cVar1S6S0P069P019P067N064(0)='1' AND  D( 2)='0' AND E( 0)='0' AND D( 3)='1' )then
          cVar2S6S0N058N068P054nsss(0) <='1';
          else
          cVar2S6S0N058N068P054nsss(0) <='0';
          end if;
        if(cVar1S7S0P069P019N067P063(0)='1' AND  B( 9)='1' AND A( 1)='0' )then
          cVar2S7S0P036P017nsss(0) <='1';
          else
          cVar2S7S0P036P017nsss(0) <='0';
          end if;
        if(cVar1S8S0P069P019N067P063(0)='1' AND  B( 9)='0' AND E( 9)='1' AND E( 0)='1' )then
          cVar2S8S0N036P065P068nsss(0) <='1';
          else
          cVar2S8S0N036P065P068nsss(0) <='0';
          end if;
        if(cVar1S9S0P069N019P036P017(0)='1' AND  D( 1)='1' )then
          cVar2S9S0P062nsss(0) <='1';
          else
          cVar2S9S0P062nsss(0) <='0';
          end if;
        if(cVar1S10S0P069N019P036P017(0)='1' AND  D( 1)='0' AND E( 0)='1' AND D( 8)='1' )then
          cVar2S10S0N062P068P067nsss(0) <='1';
          else
          cVar2S10S0N062P068P067nsss(0) <='0';
          end if;
        if(cVar1S11S0P069N019P036P017(0)='1' AND  D( 1)='0' AND E( 0)='0' AND E( 2)='1' )then
          cVar2S11S0N062N068P060nsss(0) <='1';
          else
          cVar2S11S0N062N068P060nsss(0) <='0';
          end if;
        if(cVar1S12S0P069N019P036N017(0)='1' AND  A(10)='1' AND D( 1)='1' )then
          cVar2S12S0P018P062nsss(0) <='1';
          else
          cVar2S12S0P018P062nsss(0) <='0';
          end if;
        if(cVar1S13S0P069N019P036N017(0)='1' AND  A(10)='1' AND D( 1)='0' AND E( 0)='1' )then
          cVar2S13S0P018N062P068nsss(0) <='1';
          else
          cVar2S13S0P018N062P068nsss(0) <='0';
          end if;
        if(cVar1S14S0P069N019P036N017(0)='1' AND  A(10)='0' AND A(11)='1' AND D( 2)='1' )then
          cVar2S14S0N018P016P058nsss(0) <='1';
          else
          cVar2S14S0N018P016P058nsss(0) <='0';
          end if;
        if(cVar1S15S0P069N019N036P018(0)='1' AND  E( 0)='1' AND D( 0)='1' AND A(13)='0' )then
          cVar2S15S0P068P066P012nsss(0) <='1';
          else
          cVar2S15S0P068P066P012nsss(0) <='0';
          end if;
        if(cVar1S16S0P069N019N036P018(0)='1' AND  E( 0)='0' AND D( 8)='1' AND D( 1)='1' )then
          cVar2S16S0N068P067P062nsss(0) <='1';
          else
          cVar2S16S0N068P067P062nsss(0) <='0';
          end if;
        if(cVar1S17S0P069N019N036N018(0)='1' AND  E( 2)='1' AND B( 2)='1' )then
          cVar2S17S0P060P033nsss(0) <='1';
          else
          cVar2S17S0P060P033nsss(0) <='0';
          end if;
        if(cVar1S18S0N069P063P065P017(0)='1' AND  E( 0)='1' AND D( 0)='1' )then
          cVar2S18S0P068P066nsss(0) <='1';
          else
          cVar2S18S0P068P066nsss(0) <='0';
          end if;
        if(cVar1S19S0N069P063P065P017(0)='1' AND  E( 0)='1' AND D( 0)='0' AND A( 0)='0' )then
          cVar2S19S0P068N066P019nsss(0) <='1';
          else
          cVar2S19S0P068N066P019nsss(0) <='0';
          end if;
        if(cVar1S20S0N069P063P065P017(0)='1' AND  E( 0)='0' AND E( 1)='1' )then
          cVar2S20S0N068P064nsss(0) <='1';
          else
          cVar2S20S0N068P064nsss(0) <='0';
          end if;
        if(cVar1S21S0N069P063P065P017(0)='1' AND  E( 0)='0' AND E( 1)='0' AND E( 2)='1' )then
          cVar2S21S0N068N064P060nsss(0) <='1';
          else
          cVar2S21S0N068N064P060nsss(0) <='0';
          end if;
        if(cVar1S22S0N069P063P065N017(0)='1' AND  E( 1)='1' AND A(11)='1' )then
          cVar2S22S0P064P016nsss(0) <='1';
          else
          cVar2S22S0P064P016nsss(0) <='0';
          end if;
        if(cVar1S23S0N069P063P065N017(0)='1' AND  E( 1)='1' AND A(11)='0' AND B( 0)='1' )then
          cVar2S23S0P064N016P037nsss(0) <='1';
          else
          cVar2S23S0P064N016P037nsss(0) <='0';
          end if;
        if(cVar1S24S0N069P063P065N017(0)='1' AND  E( 1)='0' AND E( 0)='1' AND A(10)='1' )then
          cVar2S24S0N064P068P018nsss(0) <='1';
          else
          cVar2S24S0N064P068P018nsss(0) <='0';
          end if;
        if(cVar1S25S0N069P063P065N017(0)='1' AND  E( 1)='0' AND E( 0)='0' AND E( 2)='1' )then
          cVar2S25S0N064N068P060nsss(0) <='1';
          else
          cVar2S25S0N064N068P060nsss(0) <='0';
          end if;
        if(cVar1S26S0N069P063N065P061(0)='1' AND  B(10)='1' AND D( 1)='1' )then
          cVar2S26S0P034P062nsss(0) <='1';
          else
          cVar2S26S0P034P062nsss(0) <='0';
          end if;
        if(cVar1S27S0N069P063N065P061(0)='1' AND  B(10)='1' AND D( 1)='0' AND E( 0)='1' )then
          cVar2S27S0P034N062P068nsss(0) <='1';
          else
          cVar2S27S0P034N062P068nsss(0) <='0';
          end if;
        if(cVar1S28S0N069N063P061P059(0)='1' AND  A( 2)='1' AND B(11)='1' )then
          cVar2S28S0P015P032nsss(0) <='1';
          else
          cVar2S28S0P015P032nsss(0) <='0';
          end if;
        if(cVar1S29S0N069N063P061P059(0)='1' AND  A( 2)='1' AND B(11)='0' AND E( 1)='1' )then
          cVar2S29S0P015N032P064nsss(0) <='1';
          else
          cVar2S29S0P015N032P064nsss(0) <='0';
          end if;
        if(cVar1S30S0N069N063P061P059(0)='1' AND  A( 2)='0' AND D( 0)='1' )then
          cVar2S30S0N015P066nsss(0) <='1';
          else
          cVar2S30S0N015P066nsss(0) <='0';
          end if;
        if(cVar1S31S0N069N063P061P059(0)='1' AND  A( 2)='0' AND D( 0)='0' AND D( 1)='1' )then
          cVar2S31S0N015N066P062nsss(0) <='1';
          else
          cVar2S31S0N015N066P062nsss(0) <='0';
          end if;
        if(cVar1S32S0N069N063N061P055(0)='1' AND  A( 3)='1' AND B(12)='1' )then
          cVar2S32S0P013P030nsss(0) <='1';
          else
          cVar2S32S0P013P030nsss(0) <='0';
          end if;
        if(cVar1S33S0N069N063N061P055(0)='1' AND  A( 3)='1' AND B(12)='0' AND D( 0)='1' )then
          cVar2S33S0P013N030P066nsss(0) <='1';
          else
          cVar2S33S0P013N030P066nsss(0) <='0';
          end if;
        if(cVar1S34S0N069N063N061P055(0)='1' AND  A( 3)='0' AND E( 0)='1' AND A(10)='1' )then
          cVar2S34S0N013P068P018nsss(0) <='1';
          else
          cVar2S34S0N013P068P018nsss(0) <='0';
          end if;
        if(cVar1S35S0N069N063N061P055(0)='1' AND  A( 3)='0' AND E( 0)='0' AND E( 1)='1' )then
          cVar2S35S0N013N068P064nsss(0) <='1';
          else
          cVar2S35S0N013N068P064nsss(0) <='0';
          end if;
        if(cVar1S36S0N069N063N061N055(0)='1' AND  D(12)='1' AND B(13)='1' AND D( 0)='1' )then
          cVar2S36S0P051P028P066nsss(0) <='1';
          else
          cVar2S36S0P051P028P066nsss(0) <='0';
          end if;
        if(cVar1S37S0N069N063N061N055(0)='1' AND  D(12)='0' AND D(13)='1' AND E( 0)='1' )then
          cVar2S37S0N051P047P068nsss(0) <='1';
          else
          cVar2S37S0N051P047P068nsss(0) <='0';
          end if;
        if(cVar1S0S1P052P050P010P068(0)='1' AND  D( 1)='0' )then
          cVar2S0S1P062nsss(0) <='1';
          else
          cVar2S0S1P062nsss(0) <='0';
          end if;
        if(cVar1S1S1P052P050P010P068(0)='1' AND  D( 1)='1' AND B( 4)='1' )then
          cVar2S1S1P062P029nsss(0) <='1';
          else
          cVar2S1S1P062P029nsss(0) <='0';
          end if;
        if(cVar1S2S1P052P050P010P068(0)='1' AND  B( 4)='1' )then
          cVar2S2S1P029nsss(0) <='1';
          else
          cVar2S2S1P029nsss(0) <='0';
          end if;
        if(cVar1S3S1P052P050P010P068(0)='1' AND  B( 4)='0' AND B(13)='1' )then
          cVar2S3S1N029P028nsss(0) <='1';
          else
          cVar2S3S1N029P028nsss(0) <='0';
          end if;
        if(cVar1S4S1P052P050N010P069(0)='1' AND  D( 0)='0' )then
          cVar2S4S1P066nsss(0) <='1';
          else
          cVar2S4S1P066nsss(0) <='0';
          end if;
        if(cVar1S5S1P052P050N010P069(0)='1' AND  D( 0)='1' AND B( 9)='0' AND A( 0)='0' )then
          cVar2S5S1P066P036P019nsss(0) <='1';
          else
          cVar2S5S1P066P036P019nsss(0) <='0';
          end if;
        if(cVar1S6S1P052P050N010N069(0)='1' AND  A(15)='1' AND E( 1)='0' )then
          cVar2S6S1P008P064nsss(0) <='1';
          else
          cVar2S6S1P008P064nsss(0) <='0';
          end if;
        if(cVar1S7S1P052P050N010N069(0)='1' AND  A(15)='0' )then
          cVar2S7S1N008psss(0) <='1';
          else
          cVar2S7S1N008psss(0) <='0';
          end if;
        if(cVar1S9S1P052N050N029P028(0)='1' AND  D( 3)='1' )then
          cVar2S9S1P054nsss(0) <='1';
          else
          cVar2S9S1P054nsss(0) <='0';
          end if;
        if(cVar1S10S1P052N050N029N028(0)='1' AND  E(13)='1' )then
          cVar2S10S1P049nsss(0) <='1';
          else
          cVar2S10S1P049nsss(0) <='0';
          end if;
        if(cVar1S11S1N052P056P031P063(0)='1' AND  D( 1)='0' )then
          cVar2S11S1P062nsss(0) <='1';
          else
          cVar2S11S1P062nsss(0) <='0';
          end if;
        if(cVar1S12S1N052P056P031P063(0)='1' AND  D( 1)='1' AND A(11)='0' )then
          cVar2S12S1P062P016nsss(0) <='1';
          else
          cVar2S12S1P062P016nsss(0) <='0';
          end if;
        if(cVar1S14S1N052P056N031P029(0)='1' AND  A( 8)='0' )then
          cVar2S14S1P003nsss(0) <='1';
          else
          cVar2S14S1P003nsss(0) <='0';
          end if;
        if(cVar1S15S1N052P056N031N029(0)='1' AND  B(12)='1' AND A(13)='1' AND E( 1)='0' )then
          cVar2S15S1P030P012P064nsss(0) <='1';
          else
          cVar2S15S1P030P012P064nsss(0) <='0';
          end if;
        if(cVar1S16S1N052P056N031N029(0)='1' AND  B(12)='1' AND A(13)='0' AND D( 3)='1' )then
          cVar2S16S1P030N012P054nsss(0) <='1';
          else
          cVar2S16S1P030N012P054nsss(0) <='0';
          end if;
        if(cVar1S17S1N052P056N031N029(0)='1' AND  B(12)='0' AND B(13)='1' )then
          cVar2S17S1N030P028nsss(0) <='1';
          else
          cVar2S17S1N030P028nsss(0) <='0';
          end if;
        if(cVar1S18S1N052P056N031N029(0)='1' AND  B(12)='0' AND B(13)='0' AND B( 5)='1' )then
          cVar2S18S1N030N028P027nsss(0) <='1';
          else
          cVar2S18S1N030N028P027nsss(0) <='0';
          end if;
        if(cVar1S19S1N052N056P060P065(0)='1' AND  B( 2)='1' AND E( 8)='0' )then
          cVar2S19S1P033P069nsss(0) <='1';
          else
          cVar2S19S1P033P069nsss(0) <='0';
          end if;
        if(cVar1S20S1N052N056P060P065(0)='1' AND  B( 2)='1' AND E( 8)='1' AND A(10)='1' )then
          cVar2S20S1P033P069P018nsss(0) <='1';
          else
          cVar2S20S1P033P069P018nsss(0) <='0';
          end if;
        if(cVar1S21S1N052N056P060P065(0)='1' AND  B( 2)='0' AND B( 1)='1' )then
          cVar2S21S1N033P035nsss(0) <='1';
          else
          cVar2S21S1N033P035nsss(0) <='0';
          end if;
        if(cVar1S22S1N052N056P060P065(0)='1' AND  B( 2)='0' AND B( 1)='0' AND B(11)='1' )then
          cVar2S22S1N033N035P032nsss(0) <='1';
          else
          cVar2S22S1N033N035P032nsss(0) <='0';
          end if;
        if(cVar1S23S1N052N056P060P065(0)='1' AND  B( 1)='1' AND D( 2)='1' AND E( 1)='1' )then
          cVar2S23S1P035P058P064nsss(0) <='1';
          else
          cVar2S23S1P035P058P064nsss(0) <='0';
          end if;
        if(cVar1S24S1N052N056P060P065(0)='1' AND  B( 1)='1' AND D( 2)='0' AND A( 0)='1' )then
          cVar2S24S1P035N058P019nsss(0) <='1';
          else
          cVar2S24S1P035N058P019nsss(0) <='0';
          end if;
        if(cVar1S25S1N052N056P060P065(0)='1' AND  B( 1)='0' AND A(12)='1' AND B(11)='1' )then
          cVar2S25S1N035P014P032nsss(0) <='1';
          else
          cVar2S25S1N035P014P032nsss(0) <='0';
          end if;
        if(cVar1S26S1N052N056N060P046(0)='1' AND  A(16)='1' )then
          cVar2S26S1P006nsss(0) <='1';
          else
          cVar2S26S1P006nsss(0) <='0';
          end if;
        if(cVar1S27S1N052N056N060P046(0)='1' AND  A(16)='0' AND A(15)='1' )then
          cVar2S27S1N006P008nsss(0) <='1';
          else
          cVar2S27S1N006P008nsss(0) <='0';
          end if;
        if(cVar1S28S1N052N056N060P046(0)='1' AND  A(16)='0' AND A(15)='0' AND B( 5)='1' )then
          cVar2S28S1N006N008P027nsss(0) <='1';
          else
          cVar2S28S1N006N008P027nsss(0) <='0';
          end if;
        if(cVar1S29S1N052N056N060N046(0)='1' AND  E( 1)='1' AND D(12)='1' )then
          cVar2S29S1P064P051nsss(0) <='1';
          else
          cVar2S29S1P064P051nsss(0) <='0';
          end if;
        if(cVar1S30S1N052N056N060N046(0)='1' AND  E( 1)='1' AND D(12)='0' AND B( 1)='1' )then
          cVar2S30S1P064N051P035nsss(0) <='1';
          else
          cVar2S30S1P064N051P035nsss(0) <='0';
          end if;
        if(cVar1S31S1N052N056N060N046(0)='1' AND  E( 1)='0' AND E( 0)='0' AND E( 8)='1' )then
          cVar2S31S1N064N068P069nsss(0) <='1';
          else
          cVar2S31S1N064N068P069nsss(0) <='0';
          end if;
        if(cVar1S0S2P068P067P066P035(0)='1' AND  D(14)='1' AND B(16)='1' )then
          cVar2S0S2P043P022nsss(0) <='1';
          else
          cVar2S0S2P043P022nsss(0) <='0';
          end if;
        if(cVar1S1S2P068P067P066P035(0)='1' AND  D(14)='1' AND B(16)='0' AND E(14)='1' )then
          cVar2S1S2P043N022P045nsss(0) <='1';
          else
          cVar2S1S2P043N022P045nsss(0) <='0';
          end if;
        if(cVar1S2S2P068P067P066P035(0)='1' AND  D(14)='0' AND D(13)='0' )then
          cVar2S2S2N043P047nsss(0) <='1';
          else
          cVar2S2S2N043P047nsss(0) <='0';
          end if;
        if(cVar1S3S2P068P067P066P035(0)='1' AND  D(14)='0' AND D(13)='1' AND E(13)='1' )then
          cVar2S3S2N043P047P049nsss(0) <='1';
          else
          cVar2S3S2N043P047P049nsss(0) <='0';
          end if;
        if(cVar1S4S2P068P067P066P035(0)='1' AND  E( 1)='0' AND A( 2)='1' )then
          cVar2S4S2P064P015nsss(0) <='1';
          else
          cVar2S4S2P064P015nsss(0) <='0';
          end if;
        if(cVar1S5S2P068P067P066P035(0)='1' AND  E( 1)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar2S5S2P064N015P017nsss(0) <='1';
          else
          cVar2S5S2P064N015P017nsss(0) <='0';
          end if;
        if(cVar1S6S2P068P067P066P035(0)='1' AND  E( 1)='1' AND D(10)='0' AND D( 1)='1' )then
          cVar2S6S2P064P059P062nsss(0) <='1';
          else
          cVar2S6S2P064P059P062nsss(0) <='0';
          end if;
        if(cVar1S7S2P068P067N066P063(0)='1' AND  E( 1)='0' AND A( 0)='1' )then
          cVar2S7S2P064P019nsss(0) <='1';
          else
          cVar2S7S2P064P019nsss(0) <='0';
          end if;
        if(cVar1S8S2P068P067N066P063(0)='1' AND  E( 1)='0' AND A( 0)='0' AND A(13)='1' )then
          cVar2S8S2P064N019P012nsss(0) <='1';
          else
          cVar2S8S2P064N019P012nsss(0) <='0';
          end if;
        if(cVar1S9S2P068P067N066N063(0)='1' AND  B(13)='1' AND A(10)='0' )then
          cVar2S9S2P028P018nsss(0) <='1';
          else
          cVar2S9S2P028P018nsss(0) <='0';
          end if;
        if(cVar1S10S2P068P067N066N063(0)='1' AND  B(13)='0' AND D(15)='1' )then
          cVar2S10S2N028P039nsss(0) <='1';
          else
          cVar2S10S2N028P039nsss(0) <='0';
          end if;
        if(cVar1S11S2P068P067P035P016(0)='1' AND  A(10)='0' AND A( 0)='0' AND D( 2)='0' )then
          cVar2S11S2P018P019P058nsss(0) <='1';
          else
          cVar2S11S2P018P019P058nsss(0) <='0';
          end if;
        if(cVar1S12S2P068P067P035P016(0)='1' AND  A(10)='0' AND A( 0)='1' )then
          cVar2S12S2P018P019psss(0) <='1';
          else
          cVar2S12S2P018P019psss(0) <='0';
          end if;
        if(cVar1S13S2P068P067P035P016(0)='1' AND  A(10)='1' AND D( 0)='0' )then
          cVar2S13S2P018P066nsss(0) <='1';
          else
          cVar2S13S2P018P066nsss(0) <='0';
          end if;
        if(cVar1S14S2P068P067P035N016(0)='1' AND  A(10)='1' AND E( 8)='0' AND E( 9)='0' )then
          cVar2S14S2P018P069P065nsss(0) <='1';
          else
          cVar2S14S2P018P069P065nsss(0) <='0';
          end if;
        if(cVar1S15S2P068P067P035N016(0)='1' AND  A(10)='1' AND E( 8)='1' )then
          cVar2S15S2P018P069psss(0) <='1';
          else
          cVar2S15S2P018P069psss(0) <='0';
          end if;
        if(cVar1S16S2P068P067P035N016(0)='1' AND  A(10)='0' AND E( 6)='1' )then
          cVar2S16S2N018P044nsss(0) <='1';
          else
          cVar2S16S2N018P044nsss(0) <='0';
          end if;
        if(cVar1S18S2P068P067P035N031(0)='1' AND  A(16)='0' AND A(12)='1' AND D( 1)='1' )then
          cVar2S18S2P006P014P062nsss(0) <='1';
          else
          cVar2S18S2P006P014P062nsss(0) <='0';
          end if;
        if(cVar1S19S2N068P063P062P065(0)='1' AND  E( 2)='0' AND E( 8)='0' AND E( 1)='0' )then
          cVar2S19S2P060P069P064nsss(0) <='1';
          else
          cVar2S19S2P060P069P064nsss(0) <='0';
          end if;
        if(cVar1S20S2N068P063P062P065(0)='1' AND  E( 2)='0' AND E( 8)='1' )then
          cVar2S20S2P060P069psss(0) <='1';
          else
          cVar2S20S2P060P069psss(0) <='0';
          end if;
        if(cVar1S21S2N068P063P062P065(0)='1' AND  E( 2)='1' AND D( 2)='1' AND B( 2)='1' )then
          cVar2S21S2P060P058P033nsss(0) <='1';
          else
          cVar2S21S2P060P058P033nsss(0) <='0';
          end if;
        if(cVar1S22S2N068P063P062N065(0)='1' AND  E( 1)='1' AND A(10)='1' )then
          cVar2S22S2P064P018nsss(0) <='1';
          else
          cVar2S22S2P064P018nsss(0) <='0';
          end if;
        if(cVar1S23S2N068P063P062N065(0)='1' AND  E( 1)='0' AND E( 2)='1' AND E(10)='1' )then
          cVar2S23S2N064P060P061nsss(0) <='1';
          else
          cVar2S23S2N064P060P061nsss(0) <='0';
          end if;
        if(cVar1S24S2N068P063P062P035(0)='1' AND  D( 0)='0' AND A(14)='0' )then
          cVar2S24S2P066P010nsss(0) <='1';
          else
          cVar2S24S2P066P010nsss(0) <='0';
          end if;
        if(cVar1S25S2N068P063P062P035(0)='1' AND  E( 1)='0' AND A(12)='1' )then
          cVar2S25S2P064P014nsss(0) <='1';
          else
          cVar2S25S2P064P014nsss(0) <='0';
          end if;
        if(cVar1S26S2N068P063P062P035(0)='1' AND  E( 1)='0' AND A(12)='0' AND E( 2)='0' )then
          cVar2S26S2P064N014P060nsss(0) <='1';
          else
          cVar2S26S2P064N014P060nsss(0) <='0';
          end if;
        if(cVar1S27S2N068P063P062P035(0)='1' AND  E( 1)='1' AND A( 1)='0' AND A(12)='1' )then
          cVar2S27S2P064P017P014nsss(0) <='1';
          else
          cVar2S27S2P064P017P014nsss(0) <='0';
          end if;
        if(cVar1S28S2N068P063P062P035(0)='1' AND  E( 1)='1' AND A( 1)='1' AND B(12)='1' )then
          cVar2S28S2P064P017P030nsss(0) <='1';
          else
          cVar2S28S2P064P017P030nsss(0) <='0';
          end if;
        if(cVar1S30S2N068N063P051N028(0)='1' AND  B(14)='1' )then
          cVar2S30S2P026nsss(0) <='1';
          else
          cVar2S30S2P026nsss(0) <='0';
          end if;
        if(cVar1S31S2N068N063P051N028(0)='1' AND  B(14)='0' AND B( 4)='1' )then
          cVar2S31S2N026P029nsss(0) <='1';
          else
          cVar2S31S2N026P029nsss(0) <='0';
          end if;
        if(cVar1S32S2N068N063P051N028(0)='1' AND  B(14)='0' AND B( 4)='0' AND B( 5)='1' )then
          cVar2S32S2N026N029P027nsss(0) <='1';
          else
          cVar2S32S2N026N029P027nsss(0) <='0';
          end if;
        if(cVar1S33S2N068N063N051P067(0)='1' AND  D( 4)='1' AND E( 4)='1' )then
          cVar2S33S2P050P052nsss(0) <='1';
          else
          cVar2S33S2P050P052nsss(0) <='0';
          end if;
        if(cVar1S34S2N068N063N051P067(0)='1' AND  D( 4)='1' AND E( 4)='0' AND B( 5)='1' )then
          cVar2S34S2P050N052P027nsss(0) <='1';
          else
          cVar2S34S2P050N052P027nsss(0) <='0';
          end if;
        if(cVar1S35S2N068N063N051P067(0)='1' AND  D( 4)='0' AND D( 5)='1' )then
          cVar2S35S2N050P046nsss(0) <='1';
          else
          cVar2S35S2N050P046nsss(0) <='0';
          end if;
        if(cVar1S36S2N068N063N051P067(0)='1' AND  D( 4)='0' AND D( 5)='0' AND E( 2)='1' )then
          cVar2S36S2N050N046P060nsss(0) <='1';
          else
          cVar2S36S2N050N046P060nsss(0) <='0';
          end if;
        if(cVar1S37S2N068N063N051N067(0)='1' AND  E( 1)='1' AND B( 0)='1' AND B( 1)='0' )then
          cVar2S37S2P064P037P035nsss(0) <='1';
          else
          cVar2S37S2P064P037P035nsss(0) <='0';
          end if;
        if(cVar1S38S2N068N063N051N067(0)='1' AND  E( 1)='1' AND B( 0)='0' AND E(13)='1' )then
          cVar2S38S2P064N037P049nsss(0) <='1';
          else
          cVar2S38S2P064N037P049nsss(0) <='0';
          end if;
        if(cVar1S39S2N068N063N051N067(0)='1' AND  E( 1)='0' AND D(10)='1' )then
          cVar2S39S2N064P059nsss(0) <='1';
          else
          cVar2S39S2N064P059nsss(0) <='0';
          end if;
        if(cVar1S40S2N068N063N051N067(0)='1' AND  E( 1)='0' AND D(10)='0' AND D(11)='1' )then
          cVar2S40S2N064N059P055nsss(0) <='1';
          else
          cVar2S40S2N064N059P055nsss(0) <='0';
          end if;
        if(cVar1S1S3P043N022P007P015(0)='1' AND  B(15)='1' )then
          cVar2S1S3P024nsss(0) <='1';
          else
          cVar2S1S3P024nsss(0) <='0';
          end if;
        if(cVar1S2S3P043N022P007P015(0)='1' AND  B(15)='0' AND E( 8)='0' )then
          cVar2S2S3N024P069nsss(0) <='1';
          else
          cVar2S2S3N024P069nsss(0) <='0';
          end if;
        if(cVar1S4S3P043N022N007P049(0)='1' AND  B(15)='1' AND E(14)='1' )then
          cVar2S4S3P024P045nsss(0) <='1';
          else
          cVar2S4S3P024P045nsss(0) <='0';
          end if;
        if(cVar1S5S3P043N022N007P049(0)='1' AND  B(15)='0' AND B( 7)='1' )then
          cVar2S5S3N024P023nsss(0) <='1';
          else
          cVar2S5S3N024P023nsss(0) <='0';
          end if;
        if(cVar1S6S3P043N022N007P049(0)='1' AND  B(15)='0' AND B( 7)='0' AND A(11)='1' )then
          cVar2S6S3N024N023P016nsss(0) <='1';
          else
          cVar2S6S3N024N023P016nsss(0) <='0';
          end if;
        if(cVar1S7S3N043P067P068P060(0)='1' AND  E( 9)='0' )then
          cVar2S7S3P065nsss(0) <='1';
          else
          cVar2S7S3P065nsss(0) <='0';
          end if;
        if(cVar1S8S3N043P067P068P060(0)='1' AND  E( 9)='1' AND A(11)='1' AND E( 8)='1' )then
          cVar2S8S3P065P016P069nsss(0) <='1';
          else
          cVar2S8S3P065P016P069nsss(0) <='0';
          end if;
        if(cVar1S9S3N043P067P068P060(0)='1' AND  E( 9)='1' AND A(11)='0' AND B(13)='1' )then
          cVar2S9S3P065N016P028nsss(0) <='1';
          else
          cVar2S9S3P065N016P028nsss(0) <='0';
          end if;
        if(cVar1S10S3N043P067P068P060(0)='1' AND  A(12)='1' AND A( 1)='0' AND A(14)='0' )then
          cVar2S10S3P014P017P010nsss(0) <='1';
          else
          cVar2S10S3P014P017P010nsss(0) <='0';
          end if;
        if(cVar1S11S3N043P067P068P016(0)='1' AND  D( 1)='0' AND A( 0)='0' )then
          cVar2S11S3P062P019nsss(0) <='1';
          else
          cVar2S11S3P062P019nsss(0) <='0';
          end if;
        if(cVar1S12S3N043P067P068P016(0)='1' AND  D( 1)='0' AND A( 0)='1' AND A(10)='1' )then
          cVar2S12S3P062P019P018nsss(0) <='1';
          else
          cVar2S12S3P062P019P018nsss(0) <='0';
          end if;
        if(cVar1S13S3N043P067P068N016(0)='1' AND  A(10)='0' AND E( 8)='1' AND D( 3)='0' )then
          cVar2S13S3P018P069P054nsss(0) <='1';
          else
          cVar2S13S3P018P069P054nsss(0) <='0';
          end if;
        if(cVar1S14S3N043P067P068N016(0)='1' AND  A(10)='1' AND E( 8)='0' AND D( 0)='1' )then
          cVar2S14S3P018P069P066nsss(0) <='1';
          else
          cVar2S14S3P018P069P066nsss(0) <='0';
          end if;
        if(cVar1S15S3N043P067P068N016(0)='1' AND  A(10)='1' AND E( 8)='1' AND B(10)='1' )then
          cVar2S15S3P018P069P034nsss(0) <='1';
          else
          cVar2S15S3P018P069P034nsss(0) <='0';
          end if;
        if(cVar1S16S3N043N067P034P062(0)='1' AND  E( 9)='1' AND E( 8)='0' )then
          cVar2S16S3P065P069nsss(0) <='1';
          else
          cVar2S16S3P065P069nsss(0) <='0';
          end if;
        if(cVar1S17S3N043N067P034P062(0)='1' AND  E( 9)='1' AND E( 8)='1' AND A( 1)='1' )then
          cVar2S17S3P065P069P017nsss(0) <='1';
          else
          cVar2S17S3P065P069P017nsss(0) <='0';
          end if;
        if(cVar1S18S3N043N067P034P062(0)='1' AND  E( 9)='0' AND E(10)='1' AND B(11)='0' )then
          cVar2S18S3N065P061P032nsss(0) <='1';
          else
          cVar2S18S3N065P061P032nsss(0) <='0';
          end if;
        if(cVar1S19S3N043N067P034P062(0)='1' AND  E( 9)='0' AND E(10)='0' AND E(13)='1' )then
          cVar2S19S3N065N061P049nsss(0) <='1';
          else
          cVar2S19S3N065N061P049nsss(0) <='0';
          end if;
        if(cVar1S20S3N043N067P034P062(0)='1' AND  E( 9)='0' AND E( 1)='1' AND A(11)='1' )then
          cVar2S20S3P065P064P016nsss(0) <='1';
          else
          cVar2S20S3P065P064P016nsss(0) <='0';
          end if;
        if(cVar1S21S3N043N067P034P062(0)='1' AND  E( 9)='1' AND A(11)='0' AND E( 0)='0' )then
          cVar2S21S3P065P016P068nsss(0) <='1';
          else
          cVar2S21S3P065P016P068nsss(0) <='0';
          end if;
        if(cVar1S22S3N043N067N034P051(0)='1' AND  A( 5)='1' )then
          cVar2S22S3P009nsss(0) <='1';
          else
          cVar2S22S3P009nsss(0) <='0';
          end if;
        if(cVar1S23S3N043N067N034P051(0)='1' AND  A( 5)='0' AND A( 4)='1' )then
          cVar2S23S3N009P011nsss(0) <='1';
          else
          cVar2S23S3N009P011nsss(0) <='0';
          end if;
        if(cVar1S24S3N043N067N034P051(0)='1' AND  A( 5)='0' AND A( 4)='0' AND E( 3)='1' )then
          cVar2S24S3N009N011P056nsss(0) <='1';
          else
          cVar2S24S3N009N011P056nsss(0) <='0';
          end if;
        if(cVar1S25S3N043N067N034N051(0)='1' AND  D(15)='1' AND E(15)='1' )then
          cVar2S25S3P039P041nsss(0) <='1';
          else
          cVar2S25S3P039P041nsss(0) <='0';
          end if;
        if(cVar1S26S3N043N067N034N051(0)='1' AND  D(15)='1' AND E(15)='0' AND B(17)='1' )then
          cVar2S26S3P039N041P020nsss(0) <='1';
          else
          cVar2S26S3P039N041P020nsss(0) <='0';
          end if;
        if(cVar1S27S3N043N067N034N051(0)='1' AND  D(15)='0' AND D(13)='1' AND E( 0)='0' )then
          cVar2S27S3N039P047P068nsss(0) <='1';
          else
          cVar2S27S3N039P047P068nsss(0) <='0';
          end if;
        if(cVar1S2S4P044P023N006N004(0)='1' AND  D( 5)='0' )then
          cVar2S2S4P046nsss(0) <='1';
          else
          cVar2S2S4P046nsss(0) <='0';
          end if;
        if(cVar1S3S4P044N023P025P018(0)='1' AND  A( 1)='1' )then
          cVar2S3S4P017nsss(0) <='1';
          else
          cVar2S3S4P017nsss(0) <='0';
          end if;
        if(cVar1S4S4P044N023P025P018(0)='1' AND  A( 1)='0' AND E( 5)='0' )then
          cVar2S4S4N017P048nsss(0) <='1';
          else
          cVar2S4S4N017P048nsss(0) <='0';
          end if;
        if(cVar1S6S4P044N023N025P022(0)='1' AND  D( 6)='1' )then
          cVar2S6S4P042nsss(0) <='1';
          else
          cVar2S6S4P042nsss(0) <='0';
          end if;
        if(cVar1S7S4P044N023N025N022(0)='1' AND  A( 4)='0' AND B(15)='1' )then
          cVar2S7S4P011P024nsss(0) <='1';
          else
          cVar2S7S4P011P024nsss(0) <='0';
          end if;
        if(cVar1S8S4P044N023N025N022(0)='1' AND  A( 4)='0' AND B(15)='0' AND B( 8)='1' )then
          cVar2S8S4P011N024P021nsss(0) <='1';
          else
          cVar2S8S4P011N024P021nsss(0) <='0';
          end if;
        if(cVar1S9S4N044P037P008P067(0)='1' AND  B(10)='0' AND A(12)='0' )then
          cVar2S9S4P034P014nsss(0) <='1';
          else
          cVar2S9S4P034P014nsss(0) <='0';
          end if;
        if(cVar1S10S4N044P037P008P067(0)='1' AND  B(10)='0' AND A(12)='1' AND B( 2)='1' )then
          cVar2S10S4P034P014P033nsss(0) <='1';
          else
          cVar2S10S4P034P014P033nsss(0) <='0';
          end if;
        if(cVar1S11S4N044P037P008P067(0)='1' AND  B(10)='1' AND A( 2)='1' )then
          cVar2S11S4P034P015nsss(0) <='1';
          else
          cVar2S11S4P034P015nsss(0) <='0';
          end if;
        if(cVar1S12S4N044P037P008P067(0)='1' AND  A(11)='1' AND A(14)='0' AND A( 8)='0' )then
          cVar2S12S4P016P010P003nsss(0) <='1';
          else
          cVar2S12S4P016P010P003nsss(0) <='0';
          end if;
        if(cVar1S13S4N044P037P008P067(0)='1' AND  A(11)='0' AND A( 1)='1' )then
          cVar2S13S4N016P017nsss(0) <='1';
          else
          cVar2S13S4N016P017nsss(0) <='0';
          end if;
        if(cVar1S14S4N044P037P008P050(0)='1' AND  B( 9)='0' AND A( 2)='0' )then
          cVar2S14S4P036P015nsss(0) <='1';
          else
          cVar2S14S4P036P015nsss(0) <='0';
          end if;
        if(cVar1S15S4N044P037P008N050(0)='1' AND  A( 4)='0' AND B( 2)='0' AND E( 8)='1' )then
          cVar2S15S4P011P033P069nsss(0) <='1';
          else
          cVar2S15S4P011P033P069nsss(0) <='0';
          end if;
        if(cVar1S16S4N044P037P008N050(0)='1' AND  A( 4)='1' AND A( 6)='0' AND B(14)='1' )then
          cVar2S16S4P011P007P026nsss(0) <='1';
          else
          cVar2S16S4P011P007P026nsss(0) <='0';
          end if;
        if(cVar1S17S4N044N037P031P066(0)='1' AND  A(13)='1' AND B(12)='0' )then
          cVar2S17S4P012P030nsss(0) <='1';
          else
          cVar2S17S4P012P030nsss(0) <='0';
          end if;
        if(cVar1S18S4N044N037P031P066(0)='1' AND  A(13)='1' AND B(12)='1' AND A( 3)='0' )then
          cVar2S18S4P012P030P013nsss(0) <='1';
          else
          cVar2S18S4P012P030P013nsss(0) <='0';
          end if;
        if(cVar1S19S4N044N037P031P066(0)='1' AND  A(13)='0' AND E( 1)='1' AND D( 1)='1' )then
          cVar2S19S4N012P064P062nsss(0) <='1';
          else
          cVar2S19S4N012P064P062nsss(0) <='0';
          end if;
        if(cVar1S20S4N044N037P031P066(0)='1' AND  A(13)='0' AND E( 1)='0' )then
          cVar2S20S4N012N064psss(0) <='1';
          else
          cVar2S20S4N012N064psss(0) <='0';
          end if;
        if(cVar1S21S4N044N037P031P066(0)='1' AND  A(12)='0' AND B( 1)='0' AND E( 3)='0' )then
          cVar2S21S4P014P035P056nsss(0) <='1';
          else
          cVar2S21S4P014P035P056nsss(0) <='0';
          end if;
        if(cVar1S22S4N044N037N031P036(0)='1' AND  E( 8)='0' AND D( 9)='1' )then
          cVar2S22S4P069P063nsss(0) <='1';
          else
          cVar2S22S4P069P063nsss(0) <='0';
          end if;
        if(cVar1S23S4N044N037N031P036(0)='1' AND  E( 8)='0' AND D( 9)='0' AND E( 1)='1' )then
          cVar2S23S4P069N063P064nsss(0) <='1';
          else
          cVar2S23S4P069N063P064nsss(0) <='0';
          end if;
        if(cVar1S24S4N044N037N031P036(0)='1' AND  E( 8)='1' AND B( 4)='1' )then
          cVar2S24S4P069P029nsss(0) <='1';
          else
          cVar2S24S4P069P029nsss(0) <='0';
          end if;
        if(cVar1S25S4N044N037N031P036(0)='1' AND  E( 8)='1' AND B( 4)='0' AND D(10)='1' )then
          cVar2S25S4P069N029P059nsss(0) <='1';
          else
          cVar2S25S4P069N029P059nsss(0) <='0';
          end if;
        if(cVar1S26S4N044N037N031N036(0)='1' AND  B( 2)='1' AND E( 8)='0' )then
          cVar2S26S4P033P069nsss(0) <='1';
          else
          cVar2S26S4P033P069nsss(0) <='0';
          end if;
        if(cVar1S27S4N044N037N031N036(0)='1' AND  B( 2)='0' AND B( 1)='1' AND D( 8)='0' )then
          cVar2S27S4N033P035P067nsss(0) <='1';
          else
          cVar2S27S4N033P035P067nsss(0) <='0';
          end if;
        if(cVar1S28S4N044N037N031N036(0)='1' AND  B( 2)='0' AND B( 1)='0' AND B(12)='1' )then
          cVar2S28S4N033N035P030nsss(0) <='1';
          else
          cVar2S28S4N033N035P030nsss(0) <='0';
          end if;
        if(cVar1S1S5P027P048P052N050(0)='1' AND  A(15)='1' )then
          cVar2S1S5P008nsss(0) <='1';
          else
          cVar2S1S5P008nsss(0) <='0';
          end if;
        if(cVar1S2S5P027P048P052N050(0)='1' AND  A(15)='0' AND A( 0)='1' )then
          cVar2S2S5N008P019nsss(0) <='1';
          else
          cVar2S2S5N008P019nsss(0) <='0';
          end if;
        if(cVar1S3S5P027P048P052N050(0)='1' AND  A(15)='0' AND A( 0)='0' AND D( 5)='1' )then
          cVar2S3S5N008N019P046nsss(0) <='1';
          else
          cVar2S3S5N008N019P046nsss(0) <='0';
          end if;
        if(cVar1S6S5P027N048P050N008(0)='1' AND  E(12)='0' AND A(11)='0' )then
          cVar2S6S5P053P016nsss(0) <='1';
          else
          cVar2S6S5P053P016nsss(0) <='0';
          end if;
        if(cVar1S7S5P027N048P050N008(0)='1' AND  E(12)='0' AND A(11)='1' AND B(10)='1' )then
          cVar2S7S5P053P016P034nsss(0) <='1';
          else
          cVar2S7S5P053P016P034nsss(0) <='0';
          end if;
        if(cVar1S8S5P027N048P050N008(0)='1' AND  E(12)='1' AND A(10)='1' )then
          cVar2S8S5P053P018nsss(0) <='1';
          else
          cVar2S8S5P053P018nsss(0) <='0';
          end if;
        if(cVar1S9S5P027N048N050P049(0)='1' AND  B( 9)='0' )then
          cVar2S9S5P036nsss(0) <='1';
          else
          cVar2S9S5P036nsss(0) <='0';
          end if;
        if(cVar1S10S5P027N048N050N049(0)='1' AND  D( 7)='1' )then
          cVar2S10S5P038nsss(0) <='1';
          else
          cVar2S10S5P038nsss(0) <='0';
          end if;
        if(cVar1S11S5P027N048N050N049(0)='1' AND  D( 7)='0' AND A(13)='1' AND A( 8)='0' )then
          cVar2S11S5N038P012P003nsss(0) <='1';
          else
          cVar2S11S5N038P012P003nsss(0) <='0';
          end if;
        if(cVar1S12S5P027N048N050N049(0)='1' AND  D( 7)='0' AND A(13)='0' AND D(12)='1' )then
          cVar2S12S5N038N012P051nsss(0) <='1';
          else
          cVar2S12S5N038N012P051nsss(0) <='0';
          end if;
        if(cVar1S14S5N027P043N022P007(0)='1' AND  D( 9)='0' )then
          cVar2S14S5P063nsss(0) <='1';
          else
          cVar2S14S5P063nsss(0) <='0';
          end if;
        if(cVar1S15S5N027P043N022N007(0)='1' AND  B( 9)='1' AND D( 0)='1' )then
          cVar2S15S5P036P066nsss(0) <='1';
          else
          cVar2S15S5P036P066nsss(0) <='0';
          end if;
        if(cVar1S16S5N027P043N022N007(0)='1' AND  B( 9)='1' AND D( 0)='0' AND E( 8)='1' )then
          cVar2S16S5P036N066P069nsss(0) <='1';
          else
          cVar2S16S5P036N066P069nsss(0) <='0';
          end if;
        if(cVar1S17S5N027P043N022N007(0)='1' AND  B( 9)='0' AND A(10)='1' AND A( 1)='0' )then
          cVar2S17S5N036P018P017nsss(0) <='1';
          else
          cVar2S17S5N036P018P017nsss(0) <='0';
          end if;
        if(cVar1S18S5N027P043N022N007(0)='1' AND  B( 9)='0' AND A(10)='0' AND D(15)='1' )then
          cVar2S18S5N036N018P039nsss(0) <='1';
          else
          cVar2S18S5N036N018P039nsss(0) <='0';
          end if;
        if(cVar1S19S5N027N043P036P015(0)='1' AND  E( 3)='1' AND A( 0)='0' AND E( 0)='0' )then
          cVar2S19S5P056P019P068nsss(0) <='1';
          else
          cVar2S19S5P056P019P068nsss(0) <='0';
          end if;
        if(cVar1S20S5N027N043P036P015(0)='1' AND  E( 3)='1' AND A( 0)='1' AND E( 9)='1' )then
          cVar2S20S5P056P019P065nsss(0) <='1';
          else
          cVar2S20S5P056P019P065nsss(0) <='0';
          end if;
        if(cVar1S21S5N027N043P036P015(0)='1' AND  E( 3)='0' AND A( 0)='1' )then
          cVar2S21S5N056P019nsss(0) <='1';
          else
          cVar2S21S5N056P019nsss(0) <='0';
          end if;
        if(cVar1S22S5N027N043P036P015(0)='1' AND  E( 3)='0' AND A( 0)='0' AND A(11)='1' )then
          cVar2S22S5N056N019P016nsss(0) <='1';
          else
          cVar2S22S5N056N019P016nsss(0) <='0';
          end if;
        if(cVar1S23S5N027N043P036P015(0)='1' AND  A(11)='0' AND A( 3)='0' AND A( 4)='0' )then
          cVar2S23S5P016P013P011nsss(0) <='1';
          else
          cVar2S23S5P016P013P011nsss(0) <='0';
          end if;
        if(cVar1S24S5N027N043P036P015(0)='1' AND  A(11)='1' AND B(12)='1' AND B( 0)='0' )then
          cVar2S24S5P016P030P037nsss(0) <='1';
          else
          cVar2S24S5P016P030P037nsss(0) <='0';
          end if;
        if(cVar1S25S5N027N043P036P015(0)='1' AND  A(11)='1' AND B(12)='0' AND D(12)='1' )then
          cVar2S25S5P016N030P051nsss(0) <='1';
          else
          cVar2S25S5P016N030P051nsss(0) <='0';
          end if;
        if(cVar1S26S5N027N043N036P068(0)='1' AND  E( 9)='0' AND A(10)='1' )then
          cVar2S26S5P065P018nsss(0) <='1';
          else
          cVar2S26S5P065P018nsss(0) <='0';
          end if;
        if(cVar1S27S5N027N043N036P068(0)='1' AND  E( 9)='0' AND A(10)='0' AND E(11)='1' )then
          cVar2S27S5P065N018P057nsss(0) <='1';
          else
          cVar2S27S5P065N018P057nsss(0) <='0';
          end if;
        if(cVar1S28S5N027N043N036P068(0)='1' AND  E( 9)='1' AND A( 4)='0' AND E( 1)='0' )then
          cVar2S28S5P065P011P064nsss(0) <='1';
          else
          cVar2S28S5P065P011P064nsss(0) <='0';
          end if;
        if(cVar1S29S5N027N043N036N068(0)='1' AND  B( 4)='1' AND A(14)='1' )then
          cVar2S29S5P029P010nsss(0) <='1';
          else
          cVar2S29S5P029P010nsss(0) <='0';
          end if;
        if(cVar1S30S5N027N043N036N068(0)='1' AND  B( 4)='1' AND A(14)='0' AND D(12)='0' )then
          cVar2S30S5P029N010P051nsss(0) <='1';
          else
          cVar2S30S5P029N010P051nsss(0) <='0';
          end if;
        if(cVar1S31S5N027N043N036N068(0)='1' AND  B( 4)='0' AND E( 1)='1' AND A(11)='1' )then
          cVar2S31S5N029P064P016nsss(0) <='1';
          else
          cVar2S31S5N029P064P016nsss(0) <='0';
          end if;
        if(cVar1S32S5N027N043N036N068(0)='1' AND  B( 4)='0' AND E( 1)='0' AND D( 6)='1' )then
          cVar2S32S5N029N064P042nsss(0) <='1';
          else
          cVar2S32S5N029N064P042nsss(0) <='0';
          end if;
        if(cVar1S2S6P040N021P023N018(0)='1' AND  A( 7)='0' )then
          cVar2S2S6P005nsss(0) <='1';
          else
          cVar2S2S6P005nsss(0) <='0';
          end if;
        if(cVar1S3S6P040N021N023P020(0)='1' AND  A(10)='1' )then
          cVar2S3S6P018nsss(0) <='1';
          else
          cVar2S3S6P018nsss(0) <='0';
          end if;
        if(cVar1S4S6P040N021N023P020(0)='1' AND  A(10)='0' AND D( 7)='1' )then
          cVar2S4S6N018P038nsss(0) <='1';
          else
          cVar2S4S6N018P038nsss(0) <='0';
          end if;
        if(cVar1S5S6P040N021N023N020(0)='1' AND  B( 2)='1' AND A( 0)='1' )then
          cVar2S5S6P033P019nsss(0) <='1';
          else
          cVar2S5S6P033P019nsss(0) <='0';
          end if;
        if(cVar1S6S6P040N021N023N020(0)='1' AND  B( 2)='0' AND E(12)='1' )then
          cVar2S6S6N033P053nsss(0) <='1';
          else
          cVar2S6S6N033P053nsss(0) <='0';
          end if;
        if(cVar1S7S6N040P025P046P016(0)='1' AND  D( 6)='0' )then
          cVar2S7S6P042nsss(0) <='1';
          else
          cVar2S7S6P042nsss(0) <='0';
          end if;
        if(cVar1S8S6N040P025P046P016(0)='1' AND  E( 5)='1' )then
          cVar2S8S6P048nsss(0) <='1';
          else
          cVar2S8S6P048nsss(0) <='0';
          end if;
        if(cVar1S10S6N040P025N046N044(0)='1' AND  D( 2)='1' AND B(10)='0' )then
          cVar2S10S6P058P034nsss(0) <='1';
          else
          cVar2S10S6P058P034nsss(0) <='0';
          end if;
        if(cVar1S11S6N040P025N046N044(0)='1' AND  D( 2)='0' AND E(14)='1' )then
          cVar2S11S6N058P045nsss(0) <='1';
          else
          cVar2S11S6N058P045nsss(0) <='0';
          end if;
        if(cVar1S12S6N040P025N046N044(0)='1' AND  D( 2)='0' AND E(14)='0' AND D(13)='1' )then
          cVar2S12S6N058N045P047nsss(0) <='1';
          else
          cVar2S12S6N058N045P047nsss(0) <='0';
          end if;
        if(cVar1S13S6N040N025P056P055(0)='1' AND  A( 0)='0' )then
          cVar2S13S6P019nsss(0) <='1';
          else
          cVar2S13S6P019nsss(0) <='0';
          end if;
        if(cVar1S14S6N040N025P056P055(0)='1' AND  A( 0)='1' AND E( 8)='0' )then
          cVar2S14S6P019P069nsss(0) <='1';
          else
          cVar2S14S6P019P069nsss(0) <='0';
          end if;
        if(cVar1S15S6N040N025P056P055(0)='1' AND  A( 0)='1' AND E( 8)='1' AND D( 0)='1' )then
          cVar2S15S6P019P069P066nsss(0) <='1';
          else
          cVar2S15S6P019P069P066nsss(0) <='0';
          end if;
        if(cVar1S16S6N040N025P056P055(0)='1' AND  A(13)='1' AND A( 4)='1' )then
          cVar2S16S6P012P011nsss(0) <='1';
          else
          cVar2S16S6P012P011nsss(0) <='0';
          end if;
        if(cVar1S17S6N040N025P056P055(0)='1' AND  A(13)='1' AND A( 4)='0' AND B( 3)='1' )then
          cVar2S17S6P012N011P031nsss(0) <='1';
          else
          cVar2S17S6P012N011P031nsss(0) <='0';
          end if;
        if(cVar1S18S6N040N025P056P055(0)='1' AND  A(13)='0' AND B(13)='1' AND A(14)='1' )then
          cVar2S18S6N012P028P010nsss(0) <='1';
          else
          cVar2S18S6N012P028P010nsss(0) <='0';
          end if;
        if(cVar1S19S6N040N025P056P055(0)='1' AND  A(13)='0' AND B(13)='0' AND B( 1)='1' )then
          cVar2S19S6N012N028P035nsss(0) <='1';
          else
          cVar2S19S6N012N028P035nsss(0) <='0';
          end if;
        if(cVar1S20S6N040N025N056P060(0)='1' AND  D( 0)='0' AND D( 2)='1' )then
          cVar2S20S6P066P058nsss(0) <='1';
          else
          cVar2S20S6P066P058nsss(0) <='0';
          end if;
        if(cVar1S21S6N040N025N056P060(0)='1' AND  D( 0)='0' AND D( 2)='0' AND E(10)='0' )then
          cVar2S21S6P066N058P061nsss(0) <='1';
          else
          cVar2S21S6P066N058P061nsss(0) <='0';
          end if;
        if(cVar1S22S6N040N025N056P060(0)='1' AND  D( 0)='1' AND A( 0)='1' AND A(10)='0' )then
          cVar2S22S6P066P019P018nsss(0) <='1';
          else
          cVar2S22S6P066P019P018nsss(0) <='0';
          end if;
        if(cVar1S23S6N040N025N056N060(0)='1' AND  E(10)='1' AND D(10)='1' )then
          cVar2S23S6P061P059nsss(0) <='1';
          else
          cVar2S23S6P061P059nsss(0) <='0';
          end if;
        if(cVar1S24S6N040N025N056N060(0)='1' AND  E(10)='1' AND D(10)='0' AND D(12)='1' )then
          cVar2S24S6P061N059P051nsss(0) <='1';
          else
          cVar2S24S6P061N059P051nsss(0) <='0';
          end if;
        if(cVar1S25S6N040N025N056N060(0)='1' AND  E(10)='0' AND D( 4)='1' )then
          cVar2S25S6N061P050nsss(0) <='1';
          else
          cVar2S25S6N061P050nsss(0) <='0';
          end if;
        if(cVar1S26S6N040N025N056N060(0)='1' AND  E(10)='0' AND D( 4)='0' AND D( 0)='1' )then
          cVar2S26S6N061N050P066nsss(0) <='1';
          else
          cVar2S26S6N061N050P066nsss(0) <='0';
          end if;
        if(cVar1S2S7P066P028N055N053(0)='1' AND  A(14)='1' AND E( 4)='1' )then
          cVar2S2S7P010P052nsss(0) <='1';
          else
          cVar2S2S7P010P052nsss(0) <='0';
          end if;
        if(cVar1S3S7P066P028N055N053(0)='1' AND  A(14)='1' AND E( 4)='0' AND D( 3)='1' )then
          cVar2S3S7P010N052P054nsss(0) <='1';
          else
          cVar2S3S7P010N052P054nsss(0) <='0';
          end if;
        if(cVar1S4S7P066P028N055N053(0)='1' AND  A(14)='0' AND B( 6)='1' )then
          cVar2S4S7N010P025nsss(0) <='1';
          else
          cVar2S4S7N010P025nsss(0) <='0';
          end if;
        if(cVar1S5S7P066P028N055N053(0)='1' AND  A(14)='0' AND B( 6)='0' AND B(10)='1' )then
          cVar2S5S7N010N025P034nsss(0) <='1';
          else
          cVar2S5S7N010N025P034nsss(0) <='0';
          end if;
        if(cVar1S7S7P066N028P044N023(0)='1' AND  B( 6)='1' AND A( 1)='1' )then
          cVar2S7S7P025P017nsss(0) <='1';
          else
          cVar2S7S7P025P017nsss(0) <='0';
          end if;
        if(cVar1S8S7P066N028P044N023(0)='1' AND  B( 6)='1' AND A( 1)='0' AND A(10)='0' )then
          cVar2S8S7P025N017P018nsss(0) <='1';
          else
          cVar2S8S7P025N017P018nsss(0) <='0';
          end if;
        if(cVar1S9S7P066N028P044N023(0)='1' AND  B( 6)='0' AND A(16)='1' )then
          cVar2S9S7N025P006nsss(0) <='1';
          else
          cVar2S9S7N025P006nsss(0) <='0';
          end if;
        if(cVar1S10S7P066N028P044N023(0)='1' AND  B( 6)='0' AND A(16)='0' AND A(14)='0' )then
          cVar2S10S7N025N006P010nsss(0) <='1';
          else
          cVar2S10S7N025N006P010nsss(0) <='0';
          end if;
        if(cVar1S11S7P066N028N044P040(0)='1' AND  B( 8)='1' )then
          cVar2S11S7P021nsss(0) <='1';
          else
          cVar2S11S7P021nsss(0) <='0';
          end if;
        if(cVar1S12S7P066N028N044P040(0)='1' AND  B( 8)='0' AND B( 7)='1' )then
          cVar2S12S7N021P023nsss(0) <='1';
          else
          cVar2S12S7N021P023nsss(0) <='0';
          end if;
        if(cVar1S13S7P066N028N044P040(0)='1' AND  B( 8)='0' AND B( 7)='0' AND A( 3)='0' )then
          cVar2S13S7N021N023P013nsss(0) <='1';
          else
          cVar2S13S7N021N023P013nsss(0) <='0';
          end if;
        if(cVar1S14S7P066N028N044N040(0)='1' AND  E( 8)='1' AND A(19)='0' )then
          cVar2S14S7P069P000nsss(0) <='1';
          else
          cVar2S14S7P069P000nsss(0) <='0';
          end if;
        if(cVar1S15S7P066N028N044N040(0)='1' AND  E( 8)='0' AND B( 3)='1' )then
          cVar2S15S7N069P031nsss(0) <='1';
          else
          cVar2S15S7N069P031nsss(0) <='0';
          end if;
        if(cVar1S16S7P066N028N044N040(0)='1' AND  E( 8)='0' AND B( 3)='0' AND E( 5)='1' )then
          cVar2S16S7N069N031P048nsss(0) <='1';
          else
          cVar2S16S7N069N031P048nsss(0) <='0';
          end if;
        if(cVar1S17S7P066P065P003P067(0)='1' AND  E(15)='1' )then
          cVar2S17S7P041nsss(0) <='1';
          else
          cVar2S17S7P041nsss(0) <='0';
          end if;
        if(cVar1S18S7P066P065P003P067(0)='1' AND  E(15)='0' AND B(17)='0' AND D( 9)='1' )then
          cVar2S18S7N041P020P063nsss(0) <='1';
          else
          cVar2S18S7N041P020P063nsss(0) <='0';
          end if;
        if(cVar1S19S7P066P065P003P067(0)='1' AND  D(12)='1' AND A(15)='1' )then
          cVar2S19S7P051P008nsss(0) <='1';
          else
          cVar2S19S7P051P008nsss(0) <='0';
          end if;
        if(cVar1S20S7P066P065P003P067(0)='1' AND  D(12)='1' AND A(15)='0' AND B( 0)='1' )then
          cVar2S20S7P051N008P037nsss(0) <='1';
          else
          cVar2S20S7P051N008P037nsss(0) <='0';
          end if;
        if(cVar1S22S7P066P065P003N041(0)='1' AND  B(16)='1' )then
          cVar2S22S7P022nsss(0) <='1';
          else
          cVar2S22S7P022nsss(0) <='0';
          end if;
        if(cVar1S23S7P066P065P068P018(0)='1' AND  E( 1)='1' AND B( 1)='0' )then
          cVar2S23S7P064P035nsss(0) <='1';
          else
          cVar2S23S7P064P035nsss(0) <='0';
          end if;
        if(cVar1S24S7P066P065P068N018(0)='1' AND  A( 1)='1' AND A( 0)='0' )then
          cVar2S24S7P017P019nsss(0) <='1';
          else
          cVar2S24S7P017P019nsss(0) <='0';
          end if;
        if(cVar1S25S7P066P065P068N018(0)='1' AND  A( 1)='0' AND B( 0)='1' AND A( 0)='1' )then
          cVar2S25S7N017P037P019nsss(0) <='1';
          else
          cVar2S25S7N017P037P019nsss(0) <='0';
          end if;
        if(cVar1S26S7P066P065P068P018(0)='1' AND  A( 1)='0' AND E( 1)='0' AND D( 9)='1' )then
          cVar2S26S7P017P064P063nsss(0) <='1';
          else
          cVar2S26S7P017P064P063nsss(0) <='0';
          end if;
        if(cVar1S27S7P066P065P068P018(0)='1' AND  A( 1)='1' AND E( 8)='1' AND A(11)='1' )then
          cVar2S27S7P017P069P016nsss(0) <='1';
          else
          cVar2S27S7P017P069P016nsss(0) <='0';
          end if;
        if(cVar1S28S7P066P065P068P018(0)='1' AND  A(11)='0' AND A( 1)='0' AND B( 1)='1' )then
          cVar2S28S7P016N017P035nsss(0) <='1';
          else
          cVar2S28S7P016N017P035nsss(0) <='0';
          end if;
        if(cVar1S29S7P066P065P068P018(0)='1' AND  A(11)='1' AND D( 8)='1' AND B(10)='1' )then
          cVar2S29S7P016P067P034nsss(0) <='1';
          else
          cVar2S29S7P016P067P034nsss(0) <='0';
          end if;
        if(cVar1S1S8P043P045N064P031(0)='1' AND  E( 6)='0' AND D(13)='0' )then
          cVar2S1S8P044P047nsss(0) <='1';
          else
          cVar2S1S8P044P047nsss(0) <='0';
          end if;
        if(cVar1S2S8P043P045N064P031(0)='1' AND  E( 6)='1' AND A( 7)='1' )then
          cVar2S2S8P044P005nsss(0) <='1';
          else
          cVar2S2S8P044P005nsss(0) <='0';
          end if;
        if(cVar1S3S8P043P045N064P031(0)='1' AND  E( 6)='1' AND A( 7)='0' AND D( 5)='0' )then
          cVar2S3S8P044N005P046nsss(0) <='1';
          else
          cVar2S3S8P044N005P046nsss(0) <='0';
          end if;
        if(cVar1S5S8P043N045P005N022(0)='1' AND  A(10)='0' )then
          cVar2S5S8P018nsss(0) <='1';
          else
          cVar2S5S8P018nsss(0) <='0';
          end if;
        if(cVar1S6S8P043N045N005P022(0)='1' AND  E(15)='1' )then
          cVar2S6S8P041nsss(0) <='1';
          else
          cVar2S6S8P041nsss(0) <='0';
          end if;
        if(cVar1S7S8P043N045N005N022(0)='1' AND  E( 0)='1' AND D( 0)='1' AND A( 4)='0' )then
          cVar2S7S8P068P066P011nsss(0) <='1';
          else
          cVar2S7S8P068P066P011nsss(0) <='0';
          end if;
        if(cVar1S8S8P043N045N005N022(0)='1' AND  E( 0)='0' AND A(12)='1' AND A(10)='1' )then
          cVar2S8S8N068P014P018nsss(0) <='1';
          else
          cVar2S8S8N068P014P018nsss(0) <='0';
          end if;
        if(cVar1S10S8N043P003P040N021(0)='1' AND  A(17)='1' )then
          cVar2S10S8P004nsss(0) <='1';
          else
          cVar2S10S8P004nsss(0) <='0';
          end if;
        if(cVar1S11S8N043P003P040N021(0)='1' AND  A(17)='0' AND A( 1)='1' AND B( 0)='0' )then
          cVar2S11S8N004P017P037nsss(0) <='1';
          else
          cVar2S11S8N004P017P037nsss(0) <='0';
          end if;
        if(cVar1S12S8N043P003P040N021(0)='1' AND  A(17)='0' AND A( 1)='0' AND E(10)='1' )then
          cVar2S12S8N004N017P061nsss(0) <='1';
          else
          cVar2S12S8N004N017P061nsss(0) <='0';
          end if;
        if(cVar1S13S8N043P003N040P026(0)='1' AND  E(13)='1' )then
          cVar2S13S8P049nsss(0) <='1';
          else
          cVar2S13S8P049nsss(0) <='0';
          end if;
        if(cVar1S14S8N043P003N040P026(0)='1' AND  E(13)='0' AND D(12)='1' AND E(12)='1' )then
          cVar2S14S8N049P051P053nsss(0) <='1';
          else
          cVar2S14S8N049P051P053nsss(0) <='0';
          end if;
        if(cVar1S15S8N043P003N040P026(0)='1' AND  E(13)='0' AND D(12)='0' AND E( 3)='1' )then
          cVar2S15S8N049N051P056nsss(0) <='1';
          else
          cVar2S15S8N049N051P056nsss(0) <='0';
          end if;
        if(cVar1S16S8N043P003N040N026(0)='1' AND  E(11)='1' AND E(13)='0' AND D(11)='1' )then
          cVar2S16S8P057P049P055nsss(0) <='1';
          else
          cVar2S16S8P057P049P055nsss(0) <='0';
          end if;
        if(cVar1S17S8N043P003N040N026(0)='1' AND  E(11)='0' AND B( 6)='1' )then
          cVar2S17S8N057P025nsss(0) <='1';
          else
          cVar2S17S8N057P025nsss(0) <='0';
          end if;
        if(cVar1S18S8N043P003N040N026(0)='1' AND  E(11)='0' AND B( 6)='0' AND E( 1)='1' )then
          cVar2S18S8N057N025P064nsss(0) <='1';
          else
          cVar2S18S8N057N025P064nsss(0) <='0';
          end if;
        if(cVar1S20S8N043P003P039N020(0)='1' AND  A(11)='1' )then
          cVar2S20S8P016nsss(0) <='1';
          else
          cVar2S20S8P016nsss(0) <='0';
          end if;
        if(cVar1S21S8N043P003P039N020(0)='1' AND  A(11)='0' AND B( 8)='1' )then
          cVar2S21S8N016P021nsss(0) <='1';
          else
          cVar2S21S8N016P021nsss(0) <='0';
          end if;
        if(cVar1S22S8N043P003N039P036(0)='1' AND  A( 9)='0' AND A(14)='0' AND D( 2)='1' )then
          cVar2S22S8P001P010P058nsss(0) <='1';
          else
          cVar2S22S8P001P010P058nsss(0) <='0';
          end if;
        if(cVar1S23S8N043P003N039N036(0)='1' AND  E( 6)='1' AND A(10)='1' )then
          cVar2S23S8P044P018nsss(0) <='1';
          else
          cVar2S23S8P044P018nsss(0) <='0';
          end if;
        if(cVar1S24S8N043P003N039N036(0)='1' AND  E( 6)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar2S24S8N044P021P040nsss(0) <='1';
          else
          cVar2S24S8N044P021P040nsss(0) <='0';
          end if;
        if(cVar1S0S9P032P015P062P059(0)='1' AND  D( 0)='0' AND E( 8)='0' )then
          cVar2S0S9P066P069nsss(0) <='1';
          else
          cVar2S0S9P066P069nsss(0) <='0';
          end if;
        if(cVar1S1S9P032P015P062P059(0)='1' AND  D( 0)='0' AND E( 8)='1' AND E( 2)='0' )then
          cVar2S1S9P066P069P060nsss(0) <='1';
          else
          cVar2S1S9P066P069P060nsss(0) <='0';
          end if;
        if(cVar1S2S9P032P015P062P059(0)='1' AND  D( 0)='1' AND A(10)='1' )then
          cVar2S2S9P066P018nsss(0) <='1';
          else
          cVar2S2S9P066P018nsss(0) <='0';
          end if;
        if(cVar1S3S9P032P015P062P059(0)='1' AND  D( 0)='1' AND A(10)='0' AND E( 8)='1' )then
          cVar2S3S9P066N018P069nsss(0) <='1';
          else
          cVar2S3S9P066N018P069nsss(0) <='0';
          end if;
        if(cVar1S4S9P032P015P062N059(0)='1' AND  D( 2)='1' AND D( 8)='0' )then
          cVar2S4S9P058P067nsss(0) <='1';
          else
          cVar2S4S9P058P067nsss(0) <='0';
          end if;
        if(cVar1S5S9P032P015P062N059(0)='1' AND  D( 2)='1' AND D( 8)='1' AND B( 9)='1' )then
          cVar2S5S9P058P067P036nsss(0) <='1';
          else
          cVar2S5S9P058P067P036nsss(0) <='0';
          end if;
        if(cVar1S6S9P032P015P062N059(0)='1' AND  D( 2)='0' AND E(11)='1' )then
          cVar2S6S9N058P057nsss(0) <='1';
          else
          cVar2S6S9N058P057nsss(0) <='0';
          end if;
        if(cVar1S7S9P032P015P062N059(0)='1' AND  D( 2)='0' AND E(11)='0' AND D( 4)='1' )then
          cVar2S7S9N058N057P050nsss(0) <='1';
          else
          cVar2S7S9N058N057P050nsss(0) <='0';
          end if;
        if(cVar1S8S9P032P015P062P055(0)='1' AND  A(16)='0' AND E( 9)='1' )then
          cVar2S8S9P006P065nsss(0) <='1';
          else
          cVar2S8S9P006P065nsss(0) <='0';
          end if;
        if(cVar1S9S9P032P015P062P055(0)='1' AND  A(16)='0' AND E( 9)='0' AND E( 2)='0' )then
          cVar2S9S9P006N065P060nsss(0) <='1';
          else
          cVar2S9S9P006N065P060nsss(0) <='0';
          end if;
        if(cVar1S11S9P032P015P063N059(0)='1' AND  E( 0)='0' AND A(11)='1' )then
          cVar2S11S9P068P016nsss(0) <='1';
          else
          cVar2S11S9P068P016nsss(0) <='0';
          end if;
        if(cVar1S12S9P032P015N063P068(0)='1' AND  D(10)='1' AND E( 1)='0' )then
          cVar2S12S9P059P064nsss(0) <='1';
          else
          cVar2S12S9P059P064nsss(0) <='0';
          end if;
        if(cVar1S13S9P032P015N063P068(0)='1' AND  D(10)='0' AND D( 2)='1' )then
          cVar2S13S9N059P058nsss(0) <='1';
          else
          cVar2S13S9N059P058nsss(0) <='0';
          end if;
        if(cVar1S14S9P032P015N063N068(0)='1' AND  E( 1)='1' AND A( 1)='0' )then
          cVar2S14S9P064P017nsss(0) <='1';
          else
          cVar2S14S9P064P017nsss(0) <='0';
          end if;
        if(cVar1S15S9P032P015N063N068(0)='1' AND  E( 1)='1' AND A( 1)='1' AND A( 3)='1' )then
          cVar2S15S9P064P017P013nsss(0) <='1';
          else
          cVar2S15S9P064P017P013nsss(0) <='0';
          end if;
        if(cVar1S16S9P032P015N063N068(0)='1' AND  E( 1)='0' AND E(10)='0' AND A( 0)='0' )then
          cVar2S16S9N064P061P019nsss(0) <='1';
          else
          cVar2S16S9N064P061P019nsss(0) <='0';
          end if;
        if(cVar1S17S9P032P015N063N068(0)='1' AND  E( 1)='0' AND E(10)='1' AND E( 8)='1' )then
          cVar2S17S9N064P061P069nsss(0) <='1';
          else
          cVar2S17S9N064P061P069nsss(0) <='0';
          end if;
        if(cVar1S19S9N032P043P045N062(0)='1' AND  B(16)='1' )then
          cVar2S19S9P022nsss(0) <='1';
          else
          cVar2S19S9P022nsss(0) <='0';
          end if;
        if(cVar1S20S9N032P043P045N062(0)='1' AND  B(16)='0' AND E(13)='0' )then
          cVar2S20S9N022P049nsss(0) <='1';
          else
          cVar2S20S9N022P049nsss(0) <='0';
          end if;
        if(cVar1S22S9N032P043N045N005(0)='1' AND  E( 0)='1' AND A(13)='0' )then
          cVar2S22S9P068P012nsss(0) <='1';
          else
          cVar2S22S9P068P012nsss(0) <='0';
          end if;
        if(cVar1S23S9N032P043N045N005(0)='1' AND  E( 0)='0' AND E(15)='1' AND A( 3)='0' )then
          cVar2S23S9N068P041P013nsss(0) <='1';
          else
          cVar2S23S9N068P041P013nsss(0) <='0';
          end if;
        if(cVar1S24S9N032P043N045N005(0)='1' AND  E( 0)='0' AND E(15)='0' AND B(10)='1' )then
          cVar2S24S9N068N041P034nsss(0) <='1';
          else
          cVar2S24S9N068N041P034nsss(0) <='0';
          end if;
        if(cVar1S26S9N032N043P044N023(0)='1' AND  B( 6)='1' )then
          cVar2S26S9P025nsss(0) <='1';
          else
          cVar2S26S9P025nsss(0) <='0';
          end if;
        if(cVar1S27S9N032N043P044N023(0)='1' AND  B( 6)='0' AND B(16)='1' )then
          cVar2S27S9N025P022nsss(0) <='1';
          else
          cVar2S27S9N025P022nsss(0) <='0';
          end if;
        if(cVar1S28S9N032N043P044N023(0)='1' AND  B( 6)='0' AND B(16)='0' AND A( 5)='0' )then
          cVar2S28S9N025N022P009nsss(0) <='1';
          else
          cVar2S28S9N025N022P009nsss(0) <='0';
          end if;
        if(cVar1S29S9N032N043N044P040(0)='1' AND  B( 8)='1' )then
          cVar2S29S9P021nsss(0) <='1';
          else
          cVar2S29S9P021nsss(0) <='0';
          end if;
        if(cVar1S30S9N032N043N044P040(0)='1' AND  B( 8)='0' AND B( 7)='1' )then
          cVar2S30S9N021P023nsss(0) <='1';
          else
          cVar2S30S9N021P023nsss(0) <='0';
          end if;
        if(cVar1S31S9N032N043N044P040(0)='1' AND  B( 8)='0' AND B( 7)='0' AND E(15)='1' )then
          cVar2S31S9N021N023P041nsss(0) <='1';
          else
          cVar2S31S9N021N023P041nsss(0) <='0';
          end if;
        if(cVar1S32S9N032N043N044N040(0)='1' AND  A( 8)='0' AND B( 2)='1' AND B(10)='0' )then
          cVar2S32S9P003P033P034nsss(0) <='1';
          else
          cVar2S32S9P003P033P034nsss(0) <='0';
          end if;
        if(cVar1S33S9N032N043N044N040(0)='1' AND  A( 8)='0' AND B( 2)='0' )then
          cVar2S33S9P003N033psss(0) <='1';
          else
          cVar2S33S9P003N033psss(0) <='0';
          end if;
        if(cVar1S34S9N032N043N044N040(0)='1' AND  A( 8)='1' AND D(15)='1' AND B(17)='1' )then
          cVar2S34S9P003P039P020nsss(0) <='1';
          else
          cVar2S34S9P003P039P020nsss(0) <='0';
          end if;
        if(cVar1S35S9N032N043N044N040(0)='1' AND  A( 8)='1' AND D(15)='0' AND B( 9)='1' )then
          cVar2S35S9P003N039P036nsss(0) <='1';
          else
          cVar2S35S9P003N039P036nsss(0) <='0';
          end if;
        if(cVar1S0S10P032P015P062P061(0)='1' AND  D( 0)='0' AND E( 8)='0' )then
          cVar2S0S10P066P069nsss(0) <='1';
          else
          cVar2S0S10P066P069nsss(0) <='0';
          end if;
        if(cVar1S1S10P032P015P062P061(0)='1' AND  D( 0)='0' AND E( 8)='1' AND D( 2)='0' )then
          cVar2S1S10P066P069P058nsss(0) <='1';
          else
          cVar2S1S10P066P069P058nsss(0) <='0';
          end if;
        if(cVar1S2S10P032P015P062P061(0)='1' AND  D( 0)='1' AND E( 8)='1' )then
          cVar2S2S10P066P069nsss(0) <='1';
          else
          cVar2S2S10P066P069nsss(0) <='0';
          end if;
        if(cVar1S3S10P032P015P062P061(0)='1' AND  D( 0)='1' AND E( 8)='0' AND A(12)='1' )then
          cVar2S3S10P066N069P014nsss(0) <='1';
          else
          cVar2S3S10P066N069P014nsss(0) <='0';
          end if;
        if(cVar1S4S10P032P015P062N061(0)='1' AND  B( 2)='0' AND D(13)='1' )then
          cVar2S4S10P033P047nsss(0) <='1';
          else
          cVar2S4S10P033P047nsss(0) <='0';
          end if;
        if(cVar1S5S10P032P015P062N061(0)='1' AND  B( 2)='0' AND D(13)='0' AND A(12)='1' )then
          cVar2S5S10P033N047P014nsss(0) <='1';
          else
          cVar2S5S10P033N047P014nsss(0) <='0';
          end if;
        if(cVar1S6S10P032P015P062P055(0)='1' AND  A(16)='0' AND E( 9)='1' )then
          cVar2S6S10P006P065nsss(0) <='1';
          else
          cVar2S6S10P006P065nsss(0) <='0';
          end if;
        if(cVar1S7S10P032P015P062P055(0)='1' AND  A(16)='0' AND E( 9)='0' AND E(10)='0' )then
          cVar2S7S10P006N065P061nsss(0) <='1';
          else
          cVar2S7S10P006N065P061nsss(0) <='0';
          end if;
        if(cVar1S8S10P032P015P063P057(0)='1' AND  D(10)='1' )then
          cVar2S8S10P059nsss(0) <='1';
          else
          cVar2S8S10P059nsss(0) <='0';
          end if;
        if(cVar1S9S10P032P015P063P057(0)='1' AND  D(10)='0' AND A(11)='1' )then
          cVar2S9S10N059P016nsss(0) <='1';
          else
          cVar2S9S10N059P016nsss(0) <='0';
          end if;
        if(cVar1S10S10P032P015P063P057(0)='1' AND  D(10)='0' AND A(11)='0' AND A( 1)='0' )then
          cVar2S10S10N059N016P017nsss(0) <='1';
          else
          cVar2S10S10N059N016P017nsss(0) <='0';
          end if;
        if(cVar1S11S10P032P015N063P018(0)='1' AND  D(10)='1' AND A( 4)='0' )then
          cVar2S11S10P059P011nsss(0) <='1';
          else
          cVar2S11S10P059P011nsss(0) <='0';
          end if;
        if(cVar1S12S10P032P015N063P018(0)='1' AND  D(10)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar2S12S10N059P060P017nsss(0) <='1';
          else
          cVar2S12S10N059P060P017nsss(0) <='0';
          end if;
        if(cVar1S13S10P032P015N063N018(0)='1' AND  E(10)='0' AND D( 0)='0' )then
          cVar2S13S10P061P066nsss(0) <='1';
          else
          cVar2S13S10P061P066nsss(0) <='0';
          end if;
        if(cVar1S14S10P032P015N063N018(0)='1' AND  E(10)='1' AND E( 0)='1' )then
          cVar2S14S10P061P068nsss(0) <='1';
          else
          cVar2S14S10P061P068nsss(0) <='0';
          end if;
        if(cVar1S15S10P032P015N063N018(0)='1' AND  E(10)='1' AND E( 0)='0' AND E( 1)='1' )then
          cVar2S15S10P061N068P064nsss(0) <='1';
          else
          cVar2S15S10P061N068P064nsss(0) <='0';
          end if;
        if(cVar1S17S10N032P040N021P010(0)='1' AND  B( 9)='1' AND A( 1)='1' )then
          cVar2S17S10P036P017nsss(0) <='1';
          else
          cVar2S17S10P036P017nsss(0) <='0';
          end if;
        if(cVar1S18S10N032P040N021P010(0)='1' AND  B( 9)='1' AND A( 1)='0' AND E( 0)='0' )then
          cVar2S18S10P036N017P068nsss(0) <='1';
          else
          cVar2S18S10P036N017P068nsss(0) <='0';
          end if;
        if(cVar1S19S10N032P040N021P010(0)='1' AND  B( 9)='0' AND E( 6)='0' AND A( 8)='0' )then
          cVar2S19S10N036P044P003nsss(0) <='1';
          else
          cVar2S19S10N036P044P003nsss(0) <='0';
          end if;
        if(cVar1S20S10N032P040N021P010(0)='1' AND  B( 9)='0' AND E( 6)='1' AND D( 6)='0' )then
          cVar2S20S10N036P044P042nsss(0) <='1';
          else
          cVar2S20S10N036P044P042nsss(0) <='0';
          end if;
        if(cVar1S21S10N032P040N021P010(0)='1' AND  B( 9)='0' AND D( 6)='1' )then
          cVar2S21S10P036P042nsss(0) <='1';
          else
          cVar2S21S10P036P042nsss(0) <='0';
          end if;
        if(cVar1S22S10N032P040N021P010(0)='1' AND  B( 9)='0' AND D( 6)='0' AND A(10)='1' )then
          cVar2S22S10P036N042P018nsss(0) <='1';
          else
          cVar2S22S10P036N042P018nsss(0) <='0';
          end if;
        if(cVar1S23S10N032N040P043P062(0)='1' AND  E(14)='1' )then
          cVar2S23S10P045nsss(0) <='1';
          else
          cVar2S23S10P045nsss(0) <='0';
          end if;
        if(cVar1S24S10N032N040P043P062(0)='1' AND  E(14)='0' AND A( 0)='1' )then
          cVar2S24S10N045P019nsss(0) <='1';
          else
          cVar2S24S10N045P019nsss(0) <='0';
          end if;
        if(cVar1S25S10N032N040P043N062(0)='1' AND  B(16)='1' AND A( 6)='1' )then
          cVar2S25S10P022P007nsss(0) <='1';
          else
          cVar2S25S10P022P007nsss(0) <='0';
          end if;
        if(cVar1S26S10N032N040P043N062(0)='1' AND  B(16)='1' AND A( 6)='0' AND A( 7)='1' )then
          cVar2S26S10P022N007P005nsss(0) <='1';
          else
          cVar2S26S10P022N007P005nsss(0) <='0';
          end if;
        if(cVar1S27S10N032N040P043N062(0)='1' AND  B(16)='0' AND B(15)='1' AND D(13)='0' )then
          cVar2S27S10N022P024P047nsss(0) <='1';
          else
          cVar2S27S10N022P024P047nsss(0) <='0';
          end if;
        if(cVar1S28S10N032N040P043N062(0)='1' AND  B(16)='0' AND B(15)='0' AND B( 7)='1' )then
          cVar2S28S10N022N024P023nsss(0) <='1';
          else
          cVar2S28S10N022N024P023nsss(0) <='0';
          end if;
        if(cVar1S29S10N032N040N043P033(0)='1' AND  D( 2)='1' AND A(12)='1' )then
          cVar2S29S10P058P014nsss(0) <='1';
          else
          cVar2S29S10P058P014nsss(0) <='0';
          end if;
        if(cVar1S30S10N032N040N043P033(0)='1' AND  D( 2)='1' AND A(12)='0' AND A(13)='1' )then
          cVar2S30S10P058N014P012nsss(0) <='1';
          else
          cVar2S30S10P058N014P012nsss(0) <='0';
          end if;
        if(cVar1S31S10N032N040N043P033(0)='1' AND  D( 2)='0' AND D(10)='1' AND A( 2)='1' )then
          cVar2S31S10N058P059P015nsss(0) <='1';
          else
          cVar2S31S10N058P059P015nsss(0) <='0';
          end if;
        if(cVar1S32S10N032N040N043N033(0)='1' AND  E( 6)='1' AND B( 7)='1' )then
          cVar2S32S10P044P023nsss(0) <='1';
          else
          cVar2S32S10P044P023nsss(0) <='0';
          end if;
        if(cVar1S33S10N032N040N043N033(0)='1' AND  E( 6)='1' AND B( 7)='0' AND A(11)='0' )then
          cVar2S33S10P044N023P016nsss(0) <='1';
          else
          cVar2S33S10P044N023P016nsss(0) <='0';
          end if;
        if(cVar1S34S10N032N040N043N033(0)='1' AND  E( 6)='0' AND D(13)='1' AND E( 0)='0' )then
          cVar2S34S10N044P047P068nsss(0) <='1';
          else
          cVar2S34S10N044P047P068nsss(0) <='0';
          end if;
        if(cVar1S35S10N032N040N043N033(0)='1' AND  E( 6)='0' AND D(13)='0' AND B(13)='1' )then
          cVar2S35S10N044N047P028nsss(0) <='1';
          else
          cVar2S35S10N044N047P028nsss(0) <='0';
          end if;
        if(cVar1S2S11P027P008N046N050(0)='1' AND  E( 8)='0' AND B( 0)='1' )then
          cVar2S2S11P069P037nsss(0) <='1';
          else
          cVar2S2S11P069P037nsss(0) <='0';
          end if;
        if(cVar1S3S11P027N008P050P052(0)='1' AND  D( 5)='0' )then
          cVar2S3S11P046nsss(0) <='1';
          else
          cVar2S3S11P046nsss(0) <='0';
          end if;
        if(cVar1S4S11P027N008P050P052(0)='1' AND  A(14)='1' )then
          cVar2S4S11P010nsss(0) <='1';
          else
          cVar2S4S11P010nsss(0) <='0';
          end if;
        if(cVar1S5S11P027N008P050P052(0)='1' AND  A(14)='0' AND E( 5)='0' AND A(16)='1' )then
          cVar2S5S11N010P048P006nsss(0) <='1';
          else
          cVar2S5S11N010P048P006nsss(0) <='0';
          end if;
        if(cVar1S6S11P027N008N050P018(0)='1' AND  E(13)='1' )then
          cVar2S6S11P049nsss(0) <='1';
          else
          cVar2S6S11P049nsss(0) <='0';
          end if;
        if(cVar1S7S11P027N008N050P018(0)='1' AND  E(13)='0' AND D( 1)='0' )then
          cVar2S7S11N049P062nsss(0) <='1';
          else
          cVar2S7S11N049P062nsss(0) <='0';
          end if;
        if(cVar1S8S11P027N008N050N018(0)='1' AND  B(15)='0' AND A( 9)='0' AND E(13)='1' )then
          cVar2S8S11P024P001P049nsss(0) <='1';
          else
          cVar2S8S11P024P001P049nsss(0) <='0';
          end if;
        if(cVar1S10S11N027P039P020N005(0)='1' AND  E(15)='1' AND D( 7)='0' )then
          cVar2S10S11P041P038nsss(0) <='1';
          else
          cVar2S10S11P041P038nsss(0) <='0';
          end if;
        if(cVar1S11S11N027P039N020P013(0)='1' AND  B(16)='1' )then
          cVar2S11S11P022nsss(0) <='1';
          else
          cVar2S11S11P022nsss(0) <='0';
          end if;
        if(cVar1S12S11N027P039N020P013(0)='1' AND  B(16)='0' AND B( 7)='1' )then
          cVar2S12S11N022P023nsss(0) <='1';
          else
          cVar2S12S11N022P023nsss(0) <='0';
          end if;
        if(cVar1S13S11N027P039N020P013(0)='1' AND  B(16)='0' AND B( 7)='0' AND A( 0)='1' )then
          cVar2S13S11N022N023P019nsss(0) <='1';
          else
          cVar2S13S11N022N023P019nsss(0) <='0';
          end if;
        if(cVar1S14S11N027P039N020P013(0)='1' AND  D( 0)='0' AND A( 0)='1' AND A( 2)='0' )then
          cVar2S14S11P066P019P015nsss(0) <='1';
          else
          cVar2S14S11P066P019P015nsss(0) <='0';
          end if;
        if(cVar1S15S11N027N039P020P034(0)='1' AND  B( 1)='0' AND D( 0)='0' )then
          cVar2S15S11P035P066nsss(0) <='1';
          else
          cVar2S15S11P035P066nsss(0) <='0';
          end if;
        if(cVar1S16S11N027N039P020P034(0)='1' AND  B( 1)='0' AND D( 0)='1' AND A( 2)='1' )then
          cVar2S16S11P035P066P015nsss(0) <='1';
          else
          cVar2S16S11P035P066P015nsss(0) <='0';
          end if;
        if(cVar1S17S11N027N039P020N034(0)='1' AND  E( 0)='1' AND E( 9)='0' )then
          cVar2S17S11P068P065nsss(0) <='1';
          else
          cVar2S17S11P068P065nsss(0) <='0';
          end if;
        if(cVar1S18S11N027N039P020N034(0)='1' AND  E( 0)='0' AND D( 3)='1' AND E(11)='0' )then
          cVar2S18S11N068P054P057nsss(0) <='1';
          else
          cVar2S18S11N068P054P057nsss(0) <='0';
          end if;
        if(cVar1S19S11N027N039P020N034(0)='1' AND  E( 0)='0' AND D( 3)='0' AND B( 1)='1' )then
          cVar2S19S11N068N054P035nsss(0) <='1';
          else
          cVar2S19S11N068N054P035nsss(0) <='0';
          end if;
        if(cVar1S20S11N027N039P020P040(0)='1' AND  D( 7)='1' )then
          cVar2S20S11P038nsss(0) <='1';
          else
          cVar2S20S11P038nsss(0) <='0';
          end if;
        if(cVar1S21S11N027N039P020P040(0)='1' AND  D( 7)='0' AND D( 6)='1' )then
          cVar2S21S11N038P042nsss(0) <='1';
          else
          cVar2S21S11N038P042nsss(0) <='0';
          end if;
        if(cVar1S22S11N027N039P020N040(0)='1' AND  A( 3)='0' AND E( 9)='1' AND A( 1)='1' )then
          cVar2S22S11P013P065P017nsss(0) <='1';
          else
          cVar2S22S11P013P065P017nsss(0) <='0';
          end if;
        if(cVar1S23S11N027N039P020N040(0)='1' AND  A( 3)='1' AND B( 3)='1' )then
          cVar2S23S11P013P031nsss(0) <='1';
          else
          cVar2S23S11P013P031nsss(0) <='0';
          end if;
        if(cVar1S0S12P035P068P032P015(0)='1' AND  D( 1)='0' )then
          cVar2S0S12P062nsss(0) <='1';
          else
          cVar2S0S12P062nsss(0) <='0';
          end if;
        if(cVar1S1S12P035P068P032P015(0)='1' AND  D( 1)='1' AND A(10)='1' AND A( 3)='0' )then
          cVar2S1S12P062P018P013nsss(0) <='1';
          else
          cVar2S1S12P062P018P013nsss(0) <='0';
          end if;
        if(cVar1S2S12P035P068P032P015(0)='1' AND  D( 1)='1' AND A(10)='0' AND B( 0)='1' )then
          cVar2S2S12P062N018P037nsss(0) <='1';
          else
          cVar2S2S12P062N018P037nsss(0) <='0';
          end if;
        if(cVar1S3S12P035P068P032P015(0)='1' AND  D( 9)='1' AND E( 8)='0' )then
          cVar2S3S12P063P069nsss(0) <='1';
          else
          cVar2S3S12P063P069nsss(0) <='0';
          end if;
        if(cVar1S4S12P035P068P032P015(0)='1' AND  D( 9)='0' AND D(11)='1' )then
          cVar2S4S12N063P055nsss(0) <='1';
          else
          cVar2S4S12N063P055nsss(0) <='0';
          end if;
        if(cVar1S5S12P035P068P032P015(0)='1' AND  D( 9)='0' AND D(11)='0' AND D( 5)='1' )then
          cVar2S5S12N063N055P046nsss(0) <='1';
          else
          cVar2S5S12N063N055P046nsss(0) <='0';
          end if;
        if(cVar1S6S12P035P068N032P036(0)='1' AND  A(12)='0' AND B(10)='0' )then
          cVar2S6S12P014P034nsss(0) <='1';
          else
          cVar2S6S12P014P034nsss(0) <='0';
          end if;
        if(cVar1S7S12P035P068N032P036(0)='1' AND  A(12)='0' AND B(10)='1' AND E( 5)='0' )then
          cVar2S7S12P014P034P048nsss(0) <='1';
          else
          cVar2S7S12P014P034P048nsss(0) <='0';
          end if;
        if(cVar1S8S12P035P068N032P036(0)='1' AND  A(12)='1' AND E( 3)='1' AND A( 1)='0' )then
          cVar2S8S12P014P056P017nsss(0) <='1';
          else
          cVar2S8S12P014P056P017nsss(0) <='0';
          end if;
        if(cVar1S9S12P035P068N032P036(0)='1' AND  A(12)='1' AND E( 3)='0' AND E( 1)='1' )then
          cVar2S9S12P014N056P064nsss(0) <='1';
          else
          cVar2S9S12P014N056P064nsss(0) <='0';
          end if;
        if(cVar1S10S12P035P068N032N036(0)='1' AND  B(10)='1' AND A( 1)='1' AND E( 2)='0' )then
          cVar2S10S12P034P017P060nsss(0) <='1';
          else
          cVar2S10S12P034P017P060nsss(0) <='0';
          end if;
        if(cVar1S11S12P035P068N032N036(0)='1' AND  B(10)='1' AND A( 1)='0' )then
          cVar2S11S12P034N017psss(0) <='1';
          else
          cVar2S11S12P034N017psss(0) <='0';
          end if;
        if(cVar1S12S12P035P068N032N036(0)='1' AND  B(10)='0' AND B( 0)='1' )then
          cVar2S12S12N034P037nsss(0) <='1';
          else
          cVar2S12S12N034P037nsss(0) <='0';
          end if;
        if(cVar1S13S12P035P068N032N036(0)='1' AND  B(10)='0' AND B( 0)='0' AND B( 2)='1' )then
          cVar2S13S12N034N037P033nsss(0) <='1';
          else
          cVar2S13S12N034N037P033nsss(0) <='0';
          end if;
        if(cVar1S14S12P035P068P028P067(0)='1' AND  A( 3)='0' AND A(13)='0' )then
          cVar2S14S12P013P012nsss(0) <='1';
          else
          cVar2S14S12P013P012nsss(0) <='0';
          end if;
        if(cVar1S15S12P035P068P028P067(0)='1' AND  A( 3)='0' AND A(13)='1' AND A(10)='0' )then
          cVar2S15S12P013P012P018nsss(0) <='1';
          else
          cVar2S15S12P013P012P018nsss(0) <='0';
          end if;
        if(cVar1S16S12P035P068P028P067(0)='1' AND  A( 3)='1' AND D(10)='1' AND A( 2)='1' )then
          cVar2S16S12P013P059P015nsss(0) <='1';
          else
          cVar2S16S12P013P059P015nsss(0) <='0';
          end if;
        if(cVar1S17S12P035P068P028P067(0)='1' AND  A( 3)='1' AND D(10)='0' AND B( 9)='1' )then
          cVar2S17S12P013N059P036nsss(0) <='1';
          else
          cVar2S17S12P013N059P036nsss(0) <='0';
          end if;
        if(cVar1S18S12P035P068P028P067(0)='1' AND  E( 1)='0' AND B( 2)='0' AND A(13)='1' )then
          cVar2S18S12P064P033P012nsss(0) <='1';
          else
          cVar2S18S12P064P033P012nsss(0) <='0';
          end if;
        if(cVar1S19S12P035P068P028P067(0)='1' AND  E( 1)='1' AND A( 1)='0' AND A( 0)='1' )then
          cVar2S19S12P064P017P019nsss(0) <='1';
          else
          cVar2S19S12P064P017P019nsss(0) <='0';
          end if;
        if(cVar1S20S12P035P068P028P018(0)='1' AND  D(11)='1' )then
          cVar2S20S12P055nsss(0) <='1';
          else
          cVar2S20S12P055nsss(0) <='0';
          end if;
        if(cVar1S21S12P035P068P028P018(0)='1' AND  D(11)='0' AND E( 8)='1' AND B( 0)='0' )then
          cVar2S21S12N055P069P037nsss(0) <='1';
          else
          cVar2S21S12N055P069P037nsss(0) <='0';
          end if;
        if(cVar1S22S12P035P068P028P018(0)='1' AND  B( 9)='1' AND D(12)='1' )then
          cVar2S22S12P036P051nsss(0) <='1';
          else
          cVar2S22S12P036P051nsss(0) <='0';
          end if;
        if(cVar1S23S12P035P068P028P018(0)='1' AND  B( 9)='0' AND E(12)='1' AND B( 0)='0' )then
          cVar2S23S12N036P053P037nsss(0) <='1';
          else
          cVar2S23S12N036P053P037nsss(0) <='0';
          end if;
        if(cVar1S24S12P035P067P066P061(0)='1' AND  D( 3)='1' )then
          cVar2S24S12P054nsss(0) <='1';
          else
          cVar2S24S12P054nsss(0) <='0';
          end if;
        if(cVar1S25S12P035P067P066P061(0)='1' AND  D( 3)='0' AND A(13)='0' AND D( 1)='1' )then
          cVar2S25S12N054P012P062nsss(0) <='1';
          else
          cVar2S25S12N054P012P062nsss(0) <='0';
          end if;
        if(cVar1S26S12P035P067P066P061(0)='1' AND  D( 3)='0' AND A(13)='1' AND D( 2)='1' )then
          cVar2S26S12N054P012P058nsss(0) <='1';
          else
          cVar2S26S12N054P012P058nsss(0) <='0';
          end if;
        if(cVar1S27S12P035P067P066P061(0)='1' AND  E( 1)='0' AND A( 8)='0' AND A( 1)='1' )then
          cVar2S27S12P064P003P017nsss(0) <='1';
          else
          cVar2S27S12P064P003P017nsss(0) <='0';
          end if;
        if(cVar1S28S12P035P067P066P061(0)='1' AND  E( 1)='1' AND B(11)='1' AND A( 0)='1' )then
          cVar2S28S12P064P032P019nsss(0) <='1';
          else
          cVar2S28S12P064P032P019nsss(0) <='0';
          end if;
        if(cVar1S29S12P035P067P066P061(0)='1' AND  E( 1)='1' AND B(11)='0' AND D(10)='0' )then
          cVar2S29S12P064N032P059nsss(0) <='1';
          else
          cVar2S29S12P064N032P059nsss(0) <='0';
          end if;
        if(cVar1S30S12P035P067P066P037(0)='1' AND  D(11)='0' AND A(13)='0' AND A( 9)='0' )then
          cVar2S30S12P055P012P001nsss(0) <='1';
          else
          cVar2S30S12P055P012P001nsss(0) <='0';
          end if;
        if(cVar1S31S12P035P067P066P037(0)='1' AND  D(11)='0' AND A(13)='1' AND E( 1)='0' )then
          cVar2S31S12P055P012P064nsss(0) <='1';
          else
          cVar2S31S12P055P012P064nsss(0) <='0';
          end if;
        if(cVar1S32S12P035P067P066N037(0)='1' AND  E( 1)='0' AND B(10)='0' AND A(14)='0' )then
          cVar2S32S12P064P034P010nsss(0) <='1';
          else
          cVar2S32S12P064P034P010nsss(0) <='0';
          end if;
        if(cVar1S33S12P035P067P068P014(0)='1' AND  A( 7)='0' AND A( 5)='0' )then
          cVar2S33S12P005P009nsss(0) <='1';
          else
          cVar2S33S12P005P009nsss(0) <='0';
          end if;
        if(cVar1S34S12P035P067P068P014(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S34S12P016P018nsss(0) <='1';
          else
          cVar2S34S12P016P018nsss(0) <='0';
          end if;
        if(cVar1S35S12P035P067P068P014(0)='1' AND  A(11)='1' AND A(10)='0' )then
          cVar2S35S12P016P018nsss(0) <='1';
          else
          cVar2S35S12P016P018nsss(0) <='0';
          end if;
        if(cVar1S36S12P035P067N068P018(0)='1' AND  A(14)='0' AND B( 9)='0' AND A( 1)='1' )then
          cVar2S36S12P010P036P017nsss(0) <='1';
          else
          cVar2S36S12P010P036P017nsss(0) <='0';
          end if;
        if(cVar1S37S12P035P067N068P018(0)='1' AND  A(14)='0' AND B( 9)='1' AND A( 1)='0' )then
          cVar2S37S12P010P036P017nsss(0) <='1';
          else
          cVar2S37S12P010P036P017nsss(0) <='0';
          end if;
        if(cVar1S38S12P035P067N068P018(0)='1' AND  E( 9)='1' AND E( 1)='0' )then
          cVar2S38S12P065P064nsss(0) <='1';
          else
          cVar2S38S12P065P064nsss(0) <='0';
          end if;
        if(cVar1S0S13P064P037P029P010(0)='1' AND  A(13)='0' )then
          cVar2S0S13P012nsss(0) <='1';
          else
          cVar2S0S13P012nsss(0) <='0';
          end if;
        if(cVar1S1S13P064P037P029P010(0)='1' AND  A(13)='1' AND E( 4)='1' )then
          cVar2S1S13P012P052nsss(0) <='1';
          else
          cVar2S1S13P012P052nsss(0) <='0';
          end if;
        if(cVar1S2S13P064P037P029N010(0)='1' AND  B( 3)='0' AND B(13)='0' )then
          cVar2S2S13P031P028nsss(0) <='1';
          else
          cVar2S2S13P031P028nsss(0) <='0';
          end if;
        if(cVar1S3S13P064P037P029N010(0)='1' AND  B( 3)='0' AND B(13)='1' AND A( 4)='1' )then
          cVar2S3S13P031P028P011nsss(0) <='1';
          else
          cVar2S3S13P031P028P011nsss(0) <='0';
          end if;
        if(cVar1S4S13P064P037P029N010(0)='1' AND  B( 3)='1' AND A(13)='1' )then
          cVar2S4S13P031P012nsss(0) <='1';
          else
          cVar2S4S13P031P012nsss(0) <='0';
          end if;
        if(cVar1S5S13P064P037N029P046(0)='1' AND  E( 5)='1' AND E( 7)='0' )then
          cVar2S5S13P048P040nsss(0) <='1';
          else
          cVar2S5S13P048P040nsss(0) <='0';
          end if;
        if(cVar1S6S13P064P037N029P046(0)='1' AND  E( 5)='0' AND B( 6)='1' )then
          cVar2S6S13N048P025nsss(0) <='1';
          else
          cVar2S6S13N048P025nsss(0) <='0';
          end if;
        if(cVar1S7S13P064P037N029P046(0)='1' AND  E( 5)='0' AND B( 6)='0' AND B( 7)='1' )then
          cVar2S7S13N048N025P023nsss(0) <='1';
          else
          cVar2S7S13N048N025P023nsss(0) <='0';
          end if;
        if(cVar1S8S13P064P037N029N046(0)='1' AND  B(12)='1' AND A(13)='1' AND D( 0)='0' )then
          cVar2S8S13P030P012P066nsss(0) <='1';
          else
          cVar2S8S13P030P012P066nsss(0) <='0';
          end if;
        if(cVar1S9S13P064P037N029N046(0)='1' AND  B(12)='1' AND A(13)='0' AND B( 9)='1' )then
          cVar2S9S13P030N012P036nsss(0) <='1';
          else
          cVar2S9S13P030N012P036nsss(0) <='0';
          end if;
        if(cVar1S10S13P064P037N029N046(0)='1' AND  B(12)='0' )then
          cVar2S10S13N030psss(0) <='1';
          else
          cVar2S10S13N030psss(0) <='0';
          end if;
        if(cVar1S11S13P064P037P067P066(0)='1' AND  A( 9)='0' AND E( 9)='0' AND B(15)='0' )then
          cVar2S11S13P001P065P024nsss(0) <='1';
          else
          cVar2S11S13P001P065P024nsss(0) <='0';
          end if;
        if(cVar1S12S13P064P037P067P066(0)='1' AND  A( 9)='0' AND E( 9)='1' AND B(10)='1' )then
          cVar2S12S13P001P065P034nsss(0) <='1';
          else
          cVar2S12S13P001P065P034nsss(0) <='0';
          end if;
        if(cVar1S13S13P064P037P067N066(0)='1' AND  D(11)='1' )then
          cVar2S13S13P055nsss(0) <='1';
          else
          cVar2S13S13P055nsss(0) <='0';
          end if;
        if(cVar1S14S13P064P037P067N066(0)='1' AND  D(11)='0' AND A( 0)='1' AND D( 2)='0' )then
          cVar2S14S13N055P019P058nsss(0) <='1';
          else
          cVar2S14S13N055P019P058nsss(0) <='0';
          end if;
        if(cVar1S15S13P064P037P067N066(0)='1' AND  D(11)='0' AND A( 0)='0' AND E( 3)='1' )then
          cVar2S15S13N055N019P056nsss(0) <='1';
          else
          cVar2S15S13N055N019P056nsss(0) <='0';
          end if;
        if(cVar1S16S13P064P037N067P060(0)='1' AND  E(13)='0' AND A( 8)='0' )then
          cVar2S16S13P049P003nsss(0) <='1';
          else
          cVar2S16S13P049P003nsss(0) <='0';
          end if;
        if(cVar1S17S13P064P037N067P060(0)='1' AND  E(13)='0' AND A( 8)='1' AND E( 0)='1' )then
          cVar2S17S13P049P003P068nsss(0) <='1';
          else
          cVar2S17S13P049P003P068nsss(0) <='0';
          end if;
        if(cVar1S18S13P064P037N067N060(0)='1' AND  A( 5)='0' AND E( 9)='1' AND D( 0)='0' )then
          cVar2S18S13P009P065P066nsss(0) <='1';
          else
          cVar2S18S13P009P065P066nsss(0) <='0';
          end if;
        if(cVar1S19S13P064P037N067N060(0)='1' AND  A( 5)='1' AND B(14)='1' AND A(10)='1' )then
          cVar2S19S13P009P026P018nsss(0) <='1';
          else
          cVar2S19S13P009P026P018nsss(0) <='0';
          end if;
        if(cVar1S20S13P064P037N067N060(0)='1' AND  A( 5)='1' AND B(14)='0' AND B( 5)='1' )then
          cVar2S20S13P009N026P027nsss(0) <='1';
          else
          cVar2S20S13P009N026P027nsss(0) <='0';
          end if;
        if(cVar1S21S13P064P010P063P061(0)='1' AND  E( 8)='0' AND D( 1)='1' )then
          cVar2S21S13P069P062nsss(0) <='1';
          else
          cVar2S21S13P069P062nsss(0) <='0';
          end if;
        if(cVar1S22S13P064P010P063P061(0)='1' AND  E( 8)='0' AND D( 1)='0' AND B( 9)='1' )then
          cVar2S22S13P069N062P036nsss(0) <='1';
          else
          cVar2S22S13P069N062P036nsss(0) <='0';
          end if;
        if(cVar1S23S13P064P010P063P061(0)='1' AND  E( 8)='1' AND D( 2)='0' AND E(11)='1' )then
          cVar2S23S13P069P058P057nsss(0) <='1';
          else
          cVar2S23S13P069P058P057nsss(0) <='0';
          end if;
        if(cVar1S24S13P064P010P063P061(0)='1' AND  B(11)='1' AND D( 0)='0' )then
          cVar2S24S13P032P066nsss(0) <='1';
          else
          cVar2S24S13P032P066nsss(0) <='0';
          end if;
        if(cVar1S25S13P064P010P063P061(0)='1' AND  B(11)='0' AND A(12)='1' AND B( 0)='0' )then
          cVar2S25S13N032P014P037nsss(0) <='1';
          else
          cVar2S25S13N032P014P037nsss(0) <='0';
          end if;
        if(cVar1S26S13P064P010P063P018(0)='1' AND  E( 9)='1' AND A( 2)='1' AND A( 4)='0' )then
          cVar2S26S13P065P015P011nsss(0) <='1';
          else
          cVar2S26S13P065P015P011nsss(0) <='0';
          end if;
        if(cVar1S27S13P064P010P063P018(0)='1' AND  E( 9)='1' AND A( 2)='0' AND A(13)='0' )then
          cVar2S27S13P065N015P012nsss(0) <='1';
          else
          cVar2S27S13P065N015P012nsss(0) <='0';
          end if;
        if(cVar1S28S13P064P010P063P018(0)='1' AND  E( 9)='0' AND D( 8)='0' AND B( 9)='1' )then
          cVar2S28S13N065P067P036nsss(0) <='1';
          else
          cVar2S28S13N065P067P036nsss(0) <='0';
          end if;
        if(cVar1S29S13P064P010P063N018(0)='1' AND  E( 9)='0' AND B( 0)='1' AND B( 9)='0' )then
          cVar2S29S13P065P037P036nsss(0) <='1';
          else
          cVar2S29S13P065P037P036nsss(0) <='0';
          end if;
        if(cVar1S30S13P064P010P063N018(0)='1' AND  E( 9)='0' AND B( 0)='0' AND A( 2)='1' )then
          cVar2S30S13P065N037P015nsss(0) <='1';
          else
          cVar2S30S13P065N037P015nsss(0) <='0';
          end if;
        if(cVar1S31S13P064P010P063N018(0)='1' AND  E( 9)='1' AND A(12)='1' AND A(11)='0' )then
          cVar2S31S13P065P014P016nsss(0) <='1';
          else
          cVar2S31S13P065P014P016nsss(0) <='0';
          end if;
        if(cVar1S32S13P064P010P063N018(0)='1' AND  E( 9)='1' AND A(12)='0' AND E( 2)='1' )then
          cVar2S32S13P065N014P060nsss(0) <='1';
          else
          cVar2S32S13P065N014P060nsss(0) <='0';
          end if;
        if(cVar1S34S13P064P010N032P061(0)='1' AND  B(12)='1' AND A( 2)='1' )then
          cVar2S34S13P030P015nsss(0) <='1';
          else
          cVar2S34S13P030P015nsss(0) <='0';
          end if;
        if(cVar1S35S13P064P010N032P061(0)='1' AND  B(12)='1' AND A( 2)='0' AND B( 1)='0' )then
          cVar2S35S13P030N015P035nsss(0) <='1';
          else
          cVar2S35S13P030N015P035nsss(0) <='0';
          end if;
        if(cVar1S36S13P064P010N032P061(0)='1' AND  B(12)='0' AND D(11)='0' AND B( 4)='1' )then
          cVar2S36S13N030P055P029nsss(0) <='1';
          else
          cVar2S36S13N030P055P029nsss(0) <='0';
          end if;
        if(cVar1S1S14P030P057N063P013(0)='1' AND  A( 4)='1' AND A(10)='0' )then
          cVar2S1S14P011P018nsss(0) <='1';
          else
          cVar2S1S14P011P018nsss(0) <='0';
          end if;
        if(cVar1S2S14P030P057N063P013(0)='1' AND  A( 4)='1' AND A(10)='1' AND E( 0)='0' )then
          cVar2S2S14P011P018P068nsss(0) <='1';
          else
          cVar2S2S14P011P018P068nsss(0) <='0';
          end if;
        if(cVar1S3S14P030P057N063P013(0)='1' AND  A( 4)='0' AND E( 1)='0' )then
          cVar2S3S14N011P064nsss(0) <='1';
          else
          cVar2S3S14N011P064nsss(0) <='0';
          end if;
        if(cVar1S4S14P030P057N063P013(0)='1' AND  A( 4)='0' AND E( 1)='1' AND B( 0)='1' )then
          cVar2S4S14N011P064P037nsss(0) <='1';
          else
          cVar2S4S14N011P064P037nsss(0) <='0';
          end if;
        if(cVar1S5S14P030P057N063P013(0)='1' AND  A(10)='1' )then
          cVar2S5S14P018nsss(0) <='1';
          else
          cVar2S5S14P018nsss(0) <='0';
          end if;
        if(cVar1S6S14P030P057N063P013(0)='1' AND  A(10)='0' AND B( 0)='1' )then
          cVar2S6S14N018P037nsss(0) <='1';
          else
          cVar2S6S14N018P037nsss(0) <='0';
          end if;
        if(cVar1S7S14P030P057N063P013(0)='1' AND  A(10)='0' AND B( 0)='0' AND D(10)='1' )then
          cVar2S7S14N018N037P059nsss(0) <='1';
          else
          cVar2S7S14N018N037P059nsss(0) <='0';
          end if;
        if(cVar1S8S14P030N057P056P037(0)='1' AND  A(15)='0' AND A( 0)='0' )then
          cVar2S8S14P008P019nsss(0) <='1';
          else
          cVar2S8S14P008P019nsss(0) <='0';
          end if;
        if(cVar1S9S14P030N057P056P037(0)='1' AND  A(15)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar2S9S14P008P019P018nsss(0) <='1';
          else
          cVar2S9S14P008P019P018nsss(0) <='0';
          end if;
        if(cVar1S10S14P030N057P056P037(0)='1' AND  E( 8)='0' AND A(13)='1' )then
          cVar2S10S14P069P012nsss(0) <='1';
          else
          cVar2S10S14P069P012nsss(0) <='0';
          end if;
        if(cVar1S11S14P030N057N056P061(0)='1' AND  A( 3)='1' AND D( 1)='0' )then
          cVar2S11S14P013P062nsss(0) <='1';
          else
          cVar2S11S14P013P062nsss(0) <='0';
          end if;
        if(cVar1S12S14P030N057N056P061(0)='1' AND  A( 3)='0' AND B(10)='0' AND A( 4)='1' )then
          cVar2S12S14N013P034P011nsss(0) <='1';
          else
          cVar2S12S14N013P034P011nsss(0) <='0';
          end if;
        if(cVar1S13S14P030N057N056N061(0)='1' AND  B( 4)='0' AND D( 1)='0' AND D(12)='1' )then
          cVar2S13S14P029N062P051nsss(0) <='1';
          else
          cVar2S13S14P029N062P051nsss(0) <='0';
          end if;
        if(cVar1S14S14N030P029P010P012(0)='1' AND  E( 1)='0' )then
          cVar2S14S14P064nsss(0) <='1';
          else
          cVar2S14S14P064nsss(0) <='0';
          end if;
        if(cVar1S15S14N030P029P010P012(0)='1' AND  E( 1)='1' AND A( 1)='1' )then
          cVar2S15S14P064P017nsss(0) <='1';
          else
          cVar2S15S14P064P017nsss(0) <='0';
          end if;
        if(cVar1S16S14N030P029P010P012(0)='1' AND  D( 1)='0' AND E( 4)='1' )then
          cVar2S16S14P062P052nsss(0) <='1';
          else
          cVar2S16S14P062P052nsss(0) <='0';
          end if;
        if(cVar1S17S14N030P029P010P012(0)='1' AND  D( 1)='0' AND E( 4)='0' AND D( 3)='1' )then
          cVar2S17S14P062N052P054nsss(0) <='1';
          else
          cVar2S17S14P062N052P054nsss(0) <='0';
          end if;
        if(cVar1S18S14N030P029N010P053(0)='1' AND  D( 4)='0' )then
          cVar2S18S14P050nsss(0) <='1';
          else
          cVar2S18S14P050nsss(0) <='0';
          end if;
        if(cVar1S19S14N030P029N010P053(0)='1' AND  D( 4)='1' AND A(12)='1' )then
          cVar2S19S14P050P014nsss(0) <='1';
          else
          cVar2S19S14P050P014nsss(0) <='0';
          end if;
        if(cVar1S20S14N030P029N010P053(0)='1' AND  D( 4)='1' AND A(12)='0' AND A(10)='1' )then
          cVar2S20S14P050N014P018nsss(0) <='1';
          else
          cVar2S20S14P050N014P018nsss(0) <='0';
          end if;
        if(cVar1S21S14N030P029N010N053(0)='1' AND  E( 4)='1' AND A(15)='1' )then
          cVar2S21S14P052P008nsss(0) <='1';
          else
          cVar2S21S14P052P008nsss(0) <='0';
          end if;
        if(cVar1S22S14N030P029N010N053(0)='1' AND  E( 4)='1' AND A(15)='0' AND A(13)='1' )then
          cVar2S22S14P052N008P012nsss(0) <='1';
          else
          cVar2S22S14P052N008P012nsss(0) <='0';
          end if;
        if(cVar1S23S14N030N029P046P068(0)='1' AND  A(19)='0' AND B(10)='0' AND E( 7)='0' )then
          cVar2S23S14P000P034P040nsss(0) <='1';
          else
          cVar2S23S14P000P034P040nsss(0) <='0';
          end if;
        if(cVar1S24S14N030N029P046P068(0)='1' AND  A(19)='0' AND B(10)='1' AND A( 1)='1' )then
          cVar2S24S14P000P034P017nsss(0) <='1';
          else
          cVar2S24S14P000P034P017nsss(0) <='0';
          end if;
        if(cVar1S25S14N030N029P046P068(0)='1' AND  B( 6)='1' AND E( 5)='1' )then
          cVar2S25S14P025P048nsss(0) <='1';
          else
          cVar2S25S14P025P048nsss(0) <='0';
          end if;
        if(cVar1S26S14N030N029P046P068(0)='1' AND  B( 6)='0' AND B( 5)='1' )then
          cVar2S26S14N025P027nsss(0) <='1';
          else
          cVar2S26S14N025P027nsss(0) <='0';
          end if;
        if(cVar1S27S14N030N029P046P068(0)='1' AND  B( 6)='0' AND B( 5)='0' AND D( 1)='1' )then
          cVar2S27S14N025N027P062nsss(0) <='1';
          else
          cVar2S27S14N025N027P062nsss(0) <='0';
          end if;
        if(cVar1S28S14N030N029N046P037(0)='1' AND  A(13)='0' AND E( 4)='0' AND A( 5)='0' )then
          cVar2S28S14P012P052P009nsss(0) <='1';
          else
          cVar2S28S14P012P052P009nsss(0) <='0';
          end if;
        if(cVar1S29S14N030N029N046P037(0)='1' AND  A(13)='0' AND E( 4)='1' AND B( 5)='1' )then
          cVar2S29S14P012P052P027nsss(0) <='1';
          else
          cVar2S29S14P012P052P027nsss(0) <='0';
          end if;
        if(cVar1S30S14N030N029N046P037(0)='1' AND  A(13)='1' AND B( 3)='1' AND D( 1)='0' )then
          cVar2S30S14P012P031P062nsss(0) <='1';
          else
          cVar2S30S14P012P031P062nsss(0) <='0';
          end if;
        if(cVar1S31S14N030N029N046N037(0)='1' AND  E( 7)='1' AND B( 8)='1' )then
          cVar2S31S14P040P021nsss(0) <='1';
          else
          cVar2S31S14P040P021nsss(0) <='0';
          end if;
        if(cVar1S32S14N030N029N046N037(0)='1' AND  E( 7)='1' AND B( 8)='0' AND A( 3)='0' )then
          cVar2S32S14P040N021P013nsss(0) <='1';
          else
          cVar2S32S14P040N021P013nsss(0) <='0';
          end if;
        if(cVar1S33S14N030N029N046N037(0)='1' AND  E( 7)='0' AND B(11)='1' AND A( 3)='1' )then
          cVar2S33S14N040P032P013nsss(0) <='1';
          else
          cVar2S33S14N040P032P013nsss(0) <='0';
          end if;
        if(cVar1S2S15P037P039N020N022(0)='1' AND  B( 8)='1' AND D( 7)='0' )then
          cVar2S2S15P021P038nsss(0) <='1';
          else
          cVar2S2S15P021P038nsss(0) <='0';
          end if;
        if(cVar1S3S15P037P039N020N022(0)='1' AND  B( 8)='0' AND B( 1)='1' AND D( 1)='1' )then
          cVar2S3S15N021P035P062nsss(0) <='1';
          else
          cVar2S3S15N021P035P062nsss(0) <='0';
          end if;
        if(cVar1S4S15P037P039N020N022(0)='1' AND  B( 8)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar2S4S15N021N035P026nsss(0) <='1';
          else
          cVar2S4S15N021N035P026nsss(0) <='0';
          end if;
        if(cVar1S5S15P037N039P027P050(0)='1' AND  D( 5)='0' )then
          cVar2S5S15P046nsss(0) <='1';
          else
          cVar2S5S15P046nsss(0) <='0';
          end if;
        if(cVar1S6S15P037N039P027P050(0)='1' AND  D( 5)='1' AND A( 5)='1' )then
          cVar2S6S15P046P009nsss(0) <='1';
          else
          cVar2S6S15P046P009nsss(0) <='0';
          end if;
        if(cVar1S7S15P037N039P027N050(0)='1' AND  A(15)='1' AND D( 5)='1' )then
          cVar2S7S15P008P046nsss(0) <='1';
          else
          cVar2S7S15P008P046nsss(0) <='0';
          end if;
        if(cVar1S8S15P037N039P027N050(0)='1' AND  A(15)='0' AND E(13)='1' AND A(10)='1' )then
          cVar2S8S15N008P049P018nsss(0) <='1';
          else
          cVar2S8S15N008P049P018nsss(0) <='0';
          end if;
        if(cVar1S9S15P037N039N027P026(0)='1' AND  A( 5)='1' AND A( 3)='0' AND A( 6)='0' )then
          cVar2S9S15P009P013P007nsss(0) <='1';
          else
          cVar2S9S15P009P013P007nsss(0) <='0';
          end if;
        if(cVar1S10S15P037N039N027P026(0)='1' AND  A( 5)='1' AND A( 3)='1' AND A( 4)='0' )then
          cVar2S10S15P009P013P011nsss(0) <='1';
          else
          cVar2S10S15P009P013P011nsss(0) <='0';
          end if;
        if(cVar1S11S15P037N039N027P026(0)='1' AND  A( 5)='0' AND E( 0)='0' AND A(16)='0' )then
          cVar2S11S15N009P068P006nsss(0) <='1';
          else
          cVar2S11S15N009P068P006nsss(0) <='0';
          end if;
        if(cVar1S12S15P037N039N027N026(0)='1' AND  A(15)='0' AND D( 8)='1' AND D( 2)='0' )then
          cVar2S12S15P008P067P058nsss(0) <='1';
          else
          cVar2S12S15P008P067P058nsss(0) <='0';
          end if;
        if(cVar1S13S15P037N039N027N026(0)='1' AND  A(15)='0' AND D( 8)='0' AND D( 2)='1' )then
          cVar2S13S15P008N067P058nsss(0) <='1';
          else
          cVar2S13S15P008N067P058nsss(0) <='0';
          end if;
        if(cVar1S14S15P037N039N027N026(0)='1' AND  A(15)='1' AND E( 4)='1' AND B( 4)='1' )then
          cVar2S14S15P008P052P029nsss(0) <='1';
          else
          cVar2S14S15P008P052P029nsss(0) <='0';
          end if;
        if(cVar1S16S15P037P030P057N016(0)='1' AND  E( 8)='1' )then
          cVar2S16S15P069nsss(0) <='1';
          else
          cVar2S16S15P069nsss(0) <='0';
          end if;
        if(cVar1S17S15P037P030P057N016(0)='1' AND  E( 8)='0' AND A( 0)='1' AND E( 3)='0' )then
          cVar2S17S15N069P019P056nsss(0) <='1';
          else
          cVar2S17S15N069P019P056nsss(0) <='0';
          end if;
        if(cVar1S18S15P037P030P057N016(0)='1' AND  E( 8)='0' AND A( 0)='0' AND A( 3)='1' )then
          cVar2S18S15N069N019P013nsss(0) <='1';
          else
          cVar2S18S15N069N019P013nsss(0) <='0';
          end if;
        if(cVar1S19S15P037P030N057P065(0)='1' AND  A(10)='1' )then
          cVar2S19S15P018nsss(0) <='1';
          else
          cVar2S19S15P018nsss(0) <='0';
          end if;
        if(cVar1S20S15P037P030N057P065(0)='1' AND  A(10)='0' AND A( 1)='0' )then
          cVar2S20S15N018P017nsss(0) <='1';
          else
          cVar2S20S15N018P017nsss(0) <='0';
          end if;
        if(cVar1S21S15P037N030P055P009(0)='1' AND  D(13)='1' AND B(14)='1' )then
          cVar2S21S15P047P026nsss(0) <='1';
          else
          cVar2S21S15P047P026nsss(0) <='0';
          end if;
        if(cVar1S22S15P037N030P055P009(0)='1' AND  D(13)='1' AND B(14)='0' AND A(10)='1' )then
          cVar2S22S15P047N026P018nsss(0) <='1';
          else
          cVar2S22S15P047N026P018nsss(0) <='0';
          end if;
        if(cVar1S23S15P037N030P055P009(0)='1' AND  D(13)='0' AND D( 2)='1' AND A( 1)='1' )then
          cVar2S23S15N047P058P017nsss(0) <='1';
          else
          cVar2S23S15N047P058P017nsss(0) <='0';
          end if;
        if(cVar1S24S15P037N030P055N009(0)='1' AND  D(13)='0' AND B( 3)='1' AND E(10)='0' )then
          cVar2S24S15P047P031P061nsss(0) <='1';
          else
          cVar2S24S15P047P031P061nsss(0) <='0';
          end if;
        if(cVar1S25S15P037N030P055N009(0)='1' AND  D(13)='0' AND B( 3)='0' AND B( 4)='1' )then
          cVar2S25S15P047N031P029nsss(0) <='1';
          else
          cVar2S25S15P047N031P029nsss(0) <='0';
          end if;
        if(cVar1S26S15P037N030P055N009(0)='1' AND  D(13)='1' AND A( 6)='1' AND B(15)='1' )then
          cVar2S26S15P047P007P024nsss(0) <='1';
          else
          cVar2S26S15P047P007P024nsss(0) <='0';
          end if;
        if(cVar1S27S15P037N030P055P031(0)='1' AND  A(10)='1' )then
          cVar2S27S15P018nsss(0) <='1';
          else
          cVar2S27S15P018nsss(0) <='0';
          end if;
        if(cVar1S28S15P037N030P055P031(0)='1' AND  A(10)='0' AND E( 0)='1' )then
          cVar2S28S15N018P068nsss(0) <='1';
          else
          cVar2S28S15N018P068nsss(0) <='0';
          end if;
        if(cVar1S29S15P037N030P055N031(0)='1' AND  B(13)='1' AND A(10)='0' AND E(12)='0' )then
          cVar2S29S15P028P018P053nsss(0) <='1';
          else
          cVar2S29S15P028P018P053nsss(0) <='0';
          end if;
        if(cVar1S30S15P037N030P055N031(0)='1' AND  B(13)='0' AND E( 8)='1' AND A(10)='1' )then
          cVar2S30S15N028P069P018nsss(0) <='1';
          else
          cVar2S30S15N028P069P018nsss(0) <='0';
          end if;
        if(cVar1S1S16P043P022N007P019(0)='1' AND  E( 0)='0' )then
          cVar2S1S16P068nsss(0) <='1';
          else
          cVar2S1S16P068nsss(0) <='0';
          end if;
        if(cVar1S2S16P043P022N007P019(0)='1' AND  E( 0)='1' AND A(17)='0' )then
          cVar2S2S16P068P004nsss(0) <='1';
          else
          cVar2S2S16P068P004nsss(0) <='0';
          end if;
        if(cVar1S3S16P043P022N007N019(0)='1' AND  E( 8)='0' AND A( 7)='1' )then
          cVar2S3S16P069P005nsss(0) <='1';
          else
          cVar2S3S16P069P005nsss(0) <='0';
          end if;
        if(cVar1S4S16P043P022N007N019(0)='1' AND  E( 8)='0' AND A( 7)='0' AND D( 1)='0' )then
          cVar2S4S16P069N005P062nsss(0) <='1';
          else
          cVar2S4S16P069N005P062nsss(0) <='0';
          end if;
        if(cVar1S6S16P043N022P062N016(0)='1' AND  A( 0)='1' )then
          cVar2S6S16P019nsss(0) <='1';
          else
          cVar2S6S16P019nsss(0) <='0';
          end if;
        if(cVar1S7S16P043N022N062P006(0)='1' AND  E( 0)='0' AND B(15)='1' )then
          cVar2S7S16P068P024nsss(0) <='1';
          else
          cVar2S7S16P068P024nsss(0) <='0';
          end if;
        if(cVar1S8S16P043N022N062P006(0)='1' AND  E( 0)='1' )then
          cVar2S8S16P068psss(0) <='1';
          else
          cVar2S8S16P068psss(0) <='0';
          end if;
        if(cVar1S9S16P043N022N062N006(0)='1' AND  E(13)='0' AND E( 6)='0' AND E( 5)='0' )then
          cVar2S9S16P049P044P048nsss(0) <='1';
          else
          cVar2S9S16P049P044P048nsss(0) <='0';
          end if;
        if(cVar1S10S16N043P030P057P063(0)='1' AND  D(11)='1' )then
          cVar2S10S16P055nsss(0) <='1';
          else
          cVar2S10S16P055nsss(0) <='0';
          end if;
        if(cVar1S11S16N043P030P057N063(0)='1' AND  A( 4)='1' AND A( 3)='0' )then
          cVar2S11S16P011P013nsss(0) <='1';
          else
          cVar2S11S16P011P013nsss(0) <='0';
          end if;
        if(cVar1S12S16N043P030P057N063(0)='1' AND  A( 4)='1' AND A( 3)='1' AND D( 0)='1' )then
          cVar2S12S16P011P013P066nsss(0) <='1';
          else
          cVar2S12S16P011P013P066nsss(0) <='0';
          end if;
        if(cVar1S13S16N043P030P057N063(0)='1' AND  A( 4)='0' AND A(10)='1' )then
          cVar2S13S16N011P018nsss(0) <='1';
          else
          cVar2S13S16N011P018nsss(0) <='0';
          end if;
        if(cVar1S14S16N043P030P057N063(0)='1' AND  A( 4)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar2S14S16N011N018P013nsss(0) <='1';
          else
          cVar2S14S16N011N018P013nsss(0) <='0';
          end if;
        if(cVar1S15S16N043P030N057P029(0)='1' AND  A(12)='0' AND E(10)='1' )then
          cVar2S15S16P014P061nsss(0) <='1';
          else
          cVar2S15S16P014P061nsss(0) <='0';
          end if;
        if(cVar1S16S16N043P030N057P029(0)='1' AND  A(12)='0' AND E(10)='0' AND D( 3)='1' )then
          cVar2S16S16P014N061P054nsss(0) <='1';
          else
          cVar2S16S16P014N061P054nsss(0) <='0';
          end if;
        if(cVar1S17S16N043P030N057P029(0)='1' AND  A(12)='1' AND D( 2)='1' AND D( 0)='0' )then
          cVar2S17S16P014P058P066nsss(0) <='1';
          else
          cVar2S17S16P014P058P066nsss(0) <='0';
          end if;
        if(cVar1S18S16N043P030N057P029(0)='1' AND  A(12)='1' AND D( 2)='0' AND E(12)='1' )then
          cVar2S18S16P014N058P053nsss(0) <='1';
          else
          cVar2S18S16P014N058P053nsss(0) <='0';
          end if;
        if(cVar1S19S16N043P030N057P029(0)='1' AND  A( 3)='0' AND A(13)='1' )then
          cVar2S19S16P013P012nsss(0) <='1';
          else
          cVar2S19S16P013P012nsss(0) <='0';
          end if;
        if(cVar1S20S16N043N030P039P020(0)='1' AND  A( 7)='1' )then
          cVar2S20S16P005nsss(0) <='1';
          else
          cVar2S20S16P005nsss(0) <='0';
          end if;
        if(cVar1S21S16N043N030P039P020(0)='1' AND  A( 7)='0' AND E(15)='1' )then
          cVar2S21S16N005P041nsss(0) <='1';
          else
          cVar2S21S16N005P041nsss(0) <='0';
          end if;
        if(cVar1S22S16N043N030P039N020(0)='1' AND  A( 3)='0' AND B(16)='1' )then
          cVar2S22S16P013P022nsss(0) <='1';
          else
          cVar2S22S16P013P022nsss(0) <='0';
          end if;
        if(cVar1S23S16N043N030P039N020(0)='1' AND  A( 3)='0' AND B(16)='0' AND E(12)='0' )then
          cVar2S23S16P013N022P053nsss(0) <='1';
          else
          cVar2S23S16P013N022P053nsss(0) <='0';
          end if;
        if(cVar1S24S16N043N030N039P034(0)='1' AND  B( 2)='0' AND D( 3)='0' )then
          cVar2S24S16P033P054nsss(0) <='1';
          else
          cVar2S24S16P033P054nsss(0) <='0';
          end if;
        if(cVar1S25S16N043N030N039P034(0)='1' AND  B( 2)='0' AND D( 3)='1' AND D( 9)='1' )then
          cVar2S25S16P033P054P063nsss(0) <='1';
          else
          cVar2S25S16P033P054P063nsss(0) <='0';
          end if;
        if(cVar1S26S16N043N030N039P034(0)='1' AND  B( 2)='1' AND E( 8)='1' AND A( 2)='0' )then
          cVar2S26S16P033P069P015nsss(0) <='1';
          else
          cVar2S26S16P033P069P015nsss(0) <='0';
          end if;
        if(cVar1S27S16N043N030N039P034(0)='1' AND  B( 2)='1' AND E( 8)='0' AND B( 5)='1' )then
          cVar2S27S16P033N069P027nsss(0) <='1';
          else
          cVar2S27S16P033N069P027nsss(0) <='0';
          end if;
        if(cVar1S28S16N043N030N039N034(0)='1' AND  E( 6)='1' AND B( 7)='1' )then
          cVar2S28S16P044P023nsss(0) <='1';
          else
          cVar2S28S16P044P023nsss(0) <='0';
          end if;
        if(cVar1S29S16N043N030N039N034(0)='1' AND  E( 6)='1' AND B( 7)='0' AND B(16)='1' )then
          cVar2S29S16P044N023P022nsss(0) <='1';
          else
          cVar2S29S16P044N023P022nsss(0) <='0';
          end if;
        if(cVar1S30S16N043N030N039N034(0)='1' AND  E( 6)='0' AND B( 4)='1' )then
          cVar2S30S16N044P029nsss(0) <='1';
          else
          cVar2S30S16N044P029nsss(0) <='0';
          end if;
        if(cVar1S31S16N043N030N039N034(0)='1' AND  E( 6)='0' AND B( 4)='0' AND B( 5)='1' )then
          cVar2S31S16N044N029P027nsss(0) <='1';
          else
          cVar2S31S16N044N029P027nsss(0) <='0';
          end if;
        if(cVar1S0S17P001P032P068P031(0)='1' AND  D(10)='1' AND D( 9)='1' AND D( 8)='0' )then
          cVar2S0S17P059P063P067nsss(0) <='1';
          else
          cVar2S0S17P059P063P067nsss(0) <='0';
          end if;
        if(cVar1S1S17P001P032P068P031(0)='1' AND  D(10)='1' AND D( 9)='0' )then
          cVar2S1S17P059N063psss(0) <='1';
          else
          cVar2S1S17P059N063psss(0) <='0';
          end if;
        if(cVar1S2S17P001P032P068P031(0)='1' AND  D(10)='0' AND D( 2)='1' AND B(12)='0' )then
          cVar2S2S17N059P058P030nsss(0) <='1';
          else
          cVar2S2S17N059P058P030nsss(0) <='0';
          end if;
        if(cVar1S3S17P001P032P068P031(0)='1' AND  B( 2)='0' AND A(10)='1' )then
          cVar2S3S17P033P018nsss(0) <='1';
          else
          cVar2S3S17P033P018nsss(0) <='0';
          end if;
        if(cVar1S4S17P001P032P068P031(0)='1' AND  B( 2)='0' AND A(10)='0' AND A(12)='0' )then
          cVar2S4S17P033N018P014nsss(0) <='1';
          else
          cVar2S4S17P033N018P014nsss(0) <='0';
          end if;
        if(cVar1S5S17P001P032P068P066(0)='1' AND  B( 9)='1' AND A(10)='1' )then
          cVar2S5S17P036P018nsss(0) <='1';
          else
          cVar2S5S17P036P018nsss(0) <='0';
          end if;
        if(cVar1S6S17P001P032P068P066(0)='1' AND  B( 9)='1' AND A(10)='0' AND A(12)='1' )then
          cVar2S6S17P036N018P014nsss(0) <='1';
          else
          cVar2S6S17P036N018P014nsss(0) <='0';
          end if;
        if(cVar1S7S17P001P032P068P066(0)='1' AND  B( 9)='0' AND A( 3)='1' AND D(10)='1' )then
          cVar2S7S17N036P013P059nsss(0) <='1';
          else
          cVar2S7S17N036P013P059nsss(0) <='0';
          end if;
        if(cVar1S8S17P001P032P068N066(0)='1' AND  B( 9)='0' AND A(13)='0' AND E(10)='1' )then
          cVar2S8S17P036P012P061nsss(0) <='1';
          else
          cVar2S8S17P036P012P061nsss(0) <='0';
          end if;
        if(cVar1S9S17P001N032P000P019(0)='1' AND  A( 1)='0' AND D( 3)='0' )then
          cVar2S9S17P017P054nsss(0) <='1';
          else
          cVar2S9S17P017P054nsss(0) <='0';
          end if;
        if(cVar1S10S17P001N032P000P019(0)='1' AND  A( 1)='0' AND D( 3)='1' AND E( 8)='0' )then
          cVar2S10S17P017P054P069nsss(0) <='1';
          else
          cVar2S10S17P017P054P069nsss(0) <='0';
          end if;
        if(cVar1S11S17P001N032P000P019(0)='1' AND  A( 1)='1' AND A(10)='0' AND D( 1)='1' )then
          cVar2S11S17P017P018P062nsss(0) <='1';
          else
          cVar2S11S17P017P018P062nsss(0) <='0';
          end if;
        if(cVar1S12S17P001N032P000P019(0)='1' AND  A( 1)='1' AND A(10)='1' AND B( 9)='1' )then
          cVar2S12S17P017P018P036nsss(0) <='1';
          else
          cVar2S12S17P017P018P036nsss(0) <='0';
          end if;
        if(cVar1S13S17P001N032P000N019(0)='1' AND  A( 1)='1' AND E( 0)='0' )then
          cVar2S13S17P017P068nsss(0) <='1';
          else
          cVar2S13S17P017P068nsss(0) <='0';
          end if;
        if(cVar1S14S17P001N032P000N019(0)='1' AND  A( 1)='1' AND E( 0)='1' AND A( 2)='0' )then
          cVar2S14S17P017P068P015nsss(0) <='1';
          else
          cVar2S14S17P017P068P015nsss(0) <='0';
          end if;
        if(cVar1S15S17P001N032P000N019(0)='1' AND  A( 1)='0' AND B(14)='1' AND A(17)='0' )then
          cVar2S15S17N017P026P004nsss(0) <='1';
          else
          cVar2S15S17N017P026P004nsss(0) <='0';
          end if;
        if(cVar1S16S17P001N032P000N019(0)='1' AND  A( 1)='0' AND B(14)='0' AND A(10)='1' )then
          cVar2S16S17N017N026P018nsss(0) <='1';
          else
          cVar2S16S17N017N026P018nsss(0) <='0';
          end if;
        if(cVar1S17S17P001N032P000P069(0)='1' AND  A(12)='0' AND E( 1)='0' AND A(16)='0' )then
          cVar2S17S17P014P064P006nsss(0) <='1';
          else
          cVar2S17S17P014P064P006nsss(0) <='0';
          end if;
        if(cVar1S18S17P001N032P000P069(0)='1' AND  A(12)='1' AND E( 1)='1' )then
          cVar2S18S17P014P064nsss(0) <='1';
          else
          cVar2S18S17P014P064nsss(0) <='0';
          end if;
        if(cVar1S19S17P001N032P000P069(0)='1' AND  A(12)='1' AND E( 1)='0' AND E( 0)='1' )then
          cVar2S19S17P014N064P068nsss(0) <='1';
          else
          cVar2S19S17P014N064P068nsss(0) <='0';
          end if;
        if(cVar1S20S17P001N032P000N069(0)='1' AND  A(14)='1' AND B( 2)='1' )then
          cVar2S20S17P010P033nsss(0) <='1';
          else
          cVar2S20S17P010P033nsss(0) <='0';
          end if;
        if(cVar1S21S17P001N032P000N069(0)='1' AND  A(14)='1' AND B( 2)='0' AND A(15)='0' )then
          cVar2S21S17P010N033P008nsss(0) <='1';
          else
          cVar2S21S17P010N033P008nsss(0) <='0';
          end if;
        if(cVar1S22S17P001N032P000N069(0)='1' AND  A(14)='0' AND D(15)='1' )then
          cVar2S22S17N010P039nsss(0) <='1';
          else
          cVar2S22S17N010P039nsss(0) <='0';
          end if;
        if(cVar1S23S17P001N032P000N069(0)='1' AND  A(14)='0' AND D(15)='0' AND B( 3)='1' )then
          cVar2S23S17N010N039P031nsss(0) <='1';
          else
          cVar2S23S17N010N039P031nsss(0) <='0';
          end if;
        if(cVar1S25S17P001P015N041P059(0)='1' AND  E( 0)='1' AND D( 8)='1' AND B( 0)='0' )then
          cVar2S25S17P068P067P037nsss(0) <='1';
          else
          cVar2S25S17P068P067P037nsss(0) <='0';
          end if;
        if(cVar1S26S17P001P015N041P059(0)='1' AND  E( 0)='1' AND D( 8)='0' AND A( 0)='1' )then
          cVar2S26S17P068N067P019nsss(0) <='1';
          else
          cVar2S26S17P068N067P019nsss(0) <='0';
          end if;
        if(cVar1S27S17P001P015N041P059(0)='1' AND  E( 0)='0' AND A(12)='1' AND A( 3)='0' )then
          cVar2S27S17N068P014P013nsss(0) <='1';
          else
          cVar2S27S17N068P014P013nsss(0) <='0';
          end if;
        if(cVar1S28S17P001P015N041P059(0)='1' AND  E( 0)='0' AND A(12)='0' AND A(10)='1' )then
          cVar2S28S17N068N014P018nsss(0) <='1';
          else
          cVar2S28S17N068N014P018nsss(0) <='0';
          end if;
        if(cVar1S29S17P001P015P012P066(0)='1' AND  A( 1)='0' )then
          cVar2S29S17P017nsss(0) <='1';
          else
          cVar2S29S17P017nsss(0) <='0';
          end if;
        if(cVar1S30S17P001P015P012P066(0)='1' AND  A( 1)='1' AND A(11)='0' AND A(12)='0' )then
          cVar2S30S17P017P016P014nsss(0) <='1';
          else
          cVar2S30S17P017P016P014nsss(0) <='0';
          end if;
        if(cVar1S31S17P001P015P012P066(0)='1' AND  B( 0)='1' )then
          cVar2S31S17P037nsss(0) <='1';
          else
          cVar2S31S17P037nsss(0) <='0';
          end if;
        if(cVar1S32S17P001P015N012P063(0)='1' AND  A( 7)='0' AND E(12)='0' AND B(14)='1' )then
          cVar2S32S17P005P053P026nsss(0) <='1';
          else
          cVar2S32S17P005P053P026nsss(0) <='0';
          end if;
        if(cVar1S0S18P067P037P069P031(0)='1' AND  A(13)='1' AND A(12)='0' )then
          cVar2S0S18P012P014nsss(0) <='1';
          else
          cVar2S0S18P012P014nsss(0) <='0';
          end if;
        if(cVar1S1S18P067P037P069P031(0)='1' AND  A(13)='1' AND A(12)='1' AND E( 3)='1' )then
          cVar2S1S18P012P014P056nsss(0) <='1';
          else
          cVar2S1S18P012P014P056nsss(0) <='0';
          end if;
        if(cVar1S2S18P067P037P069P031(0)='1' AND  A(13)='0' AND E( 1)='1' AND E( 2)='0' )then
          cVar2S2S18N012P064P060nsss(0) <='1';
          else
          cVar2S2S18N012P064P060nsss(0) <='0';
          end if;
        if(cVar1S3S18P067P037P069P031(0)='1' AND  A(13)='0' AND E( 1)='0' AND B(13)='1' )then
          cVar2S3S18N012N064P028nsss(0) <='1';
          else
          cVar2S3S18N012N064P028nsss(0) <='0';
          end if;
        if(cVar1S4S18P067P037P069N031(0)='1' AND  E(12)='1' AND D( 4)='0' )then
          cVar2S4S18P053P050nsss(0) <='1';
          else
          cVar2S4S18P053P050nsss(0) <='0';
          end if;
        if(cVar1S5S18P067P037P069N031(0)='1' AND  E(12)='1' AND D( 4)='1' AND B(14)='1' )then
          cVar2S5S18P053P050P026nsss(0) <='1';
          else
          cVar2S5S18P053P050P026nsss(0) <='0';
          end if;
        if(cVar1S6S18P067P037P069N031(0)='1' AND  E(12)='0' AND B( 9)='1' AND B(10)='0' )then
          cVar2S6S18N053P036P034nsss(0) <='1';
          else
          cVar2S6S18N053P036P034nsss(0) <='0';
          end if;
        if(cVar1S7S18P067P037P069N031(0)='1' AND  E(12)='0' AND B( 9)='0' )then
          cVar2S7S18N053N036psss(0) <='1';
          else
          cVar2S7S18N053N036psss(0) <='0';
          end if;
        if(cVar1S8S18P067P037P069P017(0)='1' AND  B( 9)='1' AND D( 9)='1' )then
          cVar2S8S18P036P063nsss(0) <='1';
          else
          cVar2S8S18P036P063nsss(0) <='0';
          end if;
        if(cVar1S9S18P067P037P069P017(0)='1' AND  B( 9)='0' AND A( 0)='1' AND A(14)='0' )then
          cVar2S9S18N036P019P010nsss(0) <='1';
          else
          cVar2S9S18N036P019P010nsss(0) <='0';
          end if;
        if(cVar1S10S18P067P037P069N017(0)='1' AND  E( 1)='1' AND A(10)='0' )then
          cVar2S10S18P064P018nsss(0) <='1';
          else
          cVar2S10S18P064P018nsss(0) <='0';
          end if;
        if(cVar1S11S18P067P037P069N017(0)='1' AND  E( 1)='0' AND B(11)='1' AND A(12)='0' )then
          cVar2S11S18N064P032P014nsss(0) <='1';
          else
          cVar2S11S18N064P032P014nsss(0) <='0';
          end if;
        if(cVar1S12S18P067P037P016P018(0)='1' AND  E( 0)='1' AND B( 9)='0' AND A(14)='0' )then
          cVar2S12S18P068P036P010nsss(0) <='1';
          else
          cVar2S12S18P068P036P010nsss(0) <='0';
          end if;
        if(cVar1S13S18P067P037P016P018(0)='1' AND  E( 0)='1' AND B( 9)='1' AND A( 4)='1' )then
          cVar2S13S18P068P036P011nsss(0) <='1';
          else
          cVar2S13S18P068P036P011nsss(0) <='0';
          end if;
        if(cVar1S14S18P067P037P016P018(0)='1' AND  E( 0)='0' AND E(14)='1' )then
          cVar2S14S18N068P045nsss(0) <='1';
          else
          cVar2S14S18N068P045nsss(0) <='0';
          end if;
        if(cVar1S15S18P067P037P016P018(0)='1' AND  E( 0)='0' AND E(14)='0' AND D( 0)='0' )then
          cVar2S15S18N068N045P066nsss(0) <='1';
          else
          cVar2S15S18N068N045P066nsss(0) <='0';
          end if;
        if(cVar1S16S18P067P037P016P018(0)='1' AND  B( 2)='1' AND D( 0)='1' )then
          cVar2S16S18P033P066nsss(0) <='1';
          else
          cVar2S16S18P033P066nsss(0) <='0';
          end if;
        if(cVar1S17S18P067P037P016P018(0)='1' AND  B( 2)='0' AND A(18)='0' AND B(11)='1' )then
          cVar2S17S18N033P002P032nsss(0) <='1';
          else
          cVar2S17S18N033P002P032nsss(0) <='0';
          end if;
        if(cVar1S18S18P067P037N016P019(0)='1' AND  E( 8)='1' )then
          cVar2S18S18P069nsss(0) <='1';
          else
          cVar2S18S18P069nsss(0) <='0';
          end if;
        if(cVar1S19S18P067P037N016P019(0)='1' AND  E( 8)='0' AND D(13)='0' )then
          cVar2S19S18N069P047nsss(0) <='1';
          else
          cVar2S19S18N069P047nsss(0) <='0';
          end if;
        if(cVar1S20S18P067P037N016N019(0)='1' AND  A(10)='1' AND D(11)='0' AND E( 8)='0' )then
          cVar2S20S18P018P055P069nsss(0) <='1';
          else
          cVar2S20S18P018P055P069nsss(0) <='0';
          end if;
        if(cVar1S21S18P067P037N016N019(0)='1' AND  A(10)='1' AND D(11)='1' AND A( 3)='1' )then
          cVar2S21S18P018P055P013nsss(0) <='1';
          else
          cVar2S21S18P018P055P013nsss(0) <='0';
          end if;
        if(cVar1S22S18P067P037N016N019(0)='1' AND  A(10)='0' AND A( 1)='1' AND E( 8)='1' )then
          cVar2S22S18N018P017P069nsss(0) <='1';
          else
          cVar2S22S18N018P017P069nsss(0) <='0';
          end if;
        if(cVar1S23S18P067P007P069P036(0)='1' AND  A(10)='0' AND D(11)='0' AND D( 9)='0' )then
          cVar2S23S18P018P055P063nsss(0) <='1';
          else
          cVar2S23S18P018P055P063nsss(0) <='0';
          end if;
        if(cVar1S24S18P067P007P069P036(0)='1' AND  A(10)='1' AND D( 0)='0' AND D( 1)='0' )then
          cVar2S24S18P018P066P062nsss(0) <='1';
          else
          cVar2S24S18P018P066P062nsss(0) <='0';
          end if;
        if(cVar1S25S18P067P007P069P036(0)='1' AND  A(10)='1' AND D( 0)='1' AND A(13)='1' )then
          cVar2S25S18P018P066P012nsss(0) <='1';
          else
          cVar2S25S18P018P066P012nsss(0) <='0';
          end if;
        if(cVar1S26S18P067P007P069P036(0)='1' AND  D( 0)='1' AND A(14)='0' )then
          cVar2S26S18P066P010nsss(0) <='1';
          else
          cVar2S26S18P066P010nsss(0) <='0';
          end if;
        if(cVar1S27S18P067P007P069P036(0)='1' AND  D( 0)='1' AND A(14)='1' AND A(10)='1' )then
          cVar2S27S18P066P010P018nsss(0) <='1';
          else
          cVar2S27S18P066P010P018nsss(0) <='0';
          end if;
        if(cVar1S28S18P067P007P069P036(0)='1' AND  D( 0)='0' AND D(10)='0' AND B( 2)='1' )then
          cVar2S28S18N066P059P033nsss(0) <='1';
          else
          cVar2S28S18N066P059P033nsss(0) <='0';
          end if;
        if(cVar1S29S18P067P007N069P018(0)='1' AND  A(12)='0' AND B(13)='0' )then
          cVar2S29S18P014P028nsss(0) <='1';
          else
          cVar2S29S18P014P028nsss(0) <='0';
          end if;
        if(cVar1S30S18P067P007N069P018(0)='1' AND  A(12)='1' AND B(10)='0' AND A(13)='1' )then
          cVar2S30S18P014P034P012nsss(0) <='1';
          else
          cVar2S30S18P014P034P012nsss(0) <='0';
          end if;
        if(cVar1S31S18P067P007N069N018(0)='1' AND  A( 2)='1' AND A(11)='1' AND D( 9)='1' )then
          cVar2S31S18P015P016P063nsss(0) <='1';
          else
          cVar2S31S18P015P016P063nsss(0) <='0';
          end if;
        if(cVar1S32S18P067P007N069N018(0)='1' AND  A( 2)='1' AND A(11)='0' AND E( 0)='1' )then
          cVar2S32S18P015N016P068nsss(0) <='1';
          else
          cVar2S32S18P015N016P068nsss(0) <='0';
          end if;
        if(cVar1S34S18P067P007N049P044(0)='1' AND  A( 1)='0' AND E( 9)='0' AND B( 0)='1' )then
          cVar2S34S18P017P065P037nsss(0) <='1';
          else
          cVar2S34S18P017P065P037nsss(0) <='0';
          end if;
        if(cVar1S0S19P031P012P008P060(0)='1' AND  D( 3)='0' )then
          cVar2S0S19P054nsss(0) <='1';
          else
          cVar2S0S19P054nsss(0) <='0';
          end if;
        if(cVar1S1S19P031P012P008P060(0)='1' AND  D( 3)='1' AND A( 3)='1' )then
          cVar2S1S19P054P013nsss(0) <='1';
          else
          cVar2S1S19P054P013nsss(0) <='0';
          end if;
        if(cVar1S2S19P031P012P008N060(0)='1' AND  E( 3)='1' AND D( 1)='0' )then
          cVar2S2S19P056P062nsss(0) <='1';
          else
          cVar2S2S19P056P062nsss(0) <='0';
          end if;
        if(cVar1S3S19P031P012P008N060(0)='1' AND  E( 3)='1' AND D( 1)='1' AND B( 0)='0' )then
          cVar2S3S19P056P062P037nsss(0) <='1';
          else
          cVar2S3S19P056P062P037nsss(0) <='0';
          end if;
        if(cVar1S4S19P031P012P008N060(0)='1' AND  E( 3)='0' AND D(11)='1' AND A( 3)='1' )then
          cVar2S4S19N056P055P013nsss(0) <='1';
          else
          cVar2S4S19N056P055P013nsss(0) <='0';
          end if;
        if(cVar1S5S19P031P012P008P033(0)='1' AND  E( 3)='1' )then
          cVar2S5S19P056nsss(0) <='1';
          else
          cVar2S5S19P056nsss(0) <='0';
          end if;
        if(cVar1S6S19P031P012P008P033(0)='1' AND  E( 3)='0' AND A(11)='0' )then
          cVar2S6S19N056P016nsss(0) <='1';
          else
          cVar2S6S19N056P016nsss(0) <='0';
          end if;
        if(cVar1S7S19P031N012P013P059(0)='1' AND  E( 8)='0' AND D( 1)='1' AND E( 9)='0' )then
          cVar2S7S19P069P062P065nsss(0) <='1';
          else
          cVar2S7S19P069P062P065nsss(0) <='0';
          end if;
        if(cVar1S8S19P031N012P013P059(0)='1' AND  E( 8)='0' AND D( 1)='0' )then
          cVar2S8S19P069N062psss(0) <='1';
          else
          cVar2S8S19P069N062psss(0) <='0';
          end if;
        if(cVar1S9S19P031N012P013P059(0)='1' AND  E( 8)='1' AND D(11)='1' )then
          cVar2S9S19P069P055nsss(0) <='1';
          else
          cVar2S9S19P069P055nsss(0) <='0';
          end if;
        if(cVar1S10S19P031N012P013P059(0)='1' AND  B( 0)='0' AND A(10)='1' )then
          cVar2S10S19P037P018nsss(0) <='1';
          else
          cVar2S10S19P037P018nsss(0) <='0';
          end if;
        if(cVar1S11S19P031N012P013P059(0)='1' AND  B( 0)='0' AND A(10)='0' AND A(11)='0' )then
          cVar2S11S19P037N018P016nsss(0) <='1';
          else
          cVar2S11S19P037N018P016nsss(0) <='0';
          end if;
        if(cVar1S12S19P031N012N013P054(0)='1' AND  A(12)='1' )then
          cVar2S12S19P014nsss(0) <='1';
          else
          cVar2S12S19P014nsss(0) <='0';
          end if;
        if(cVar1S13S19P031N012N013P054(0)='1' AND  A(12)='0' AND A(14)='1' )then
          cVar2S13S19N014P010nsss(0) <='1';
          else
          cVar2S13S19N014P010nsss(0) <='0';
          end if;
        if(cVar1S14S19P031N012N013N054(0)='1' AND  A( 4)='1' AND E( 8)='0' AND B( 0)='0' )then
          cVar2S14S19P011P069P037nsss(0) <='1';
          else
          cVar2S14S19P011P069P037nsss(0) <='0';
          end if;
        if(cVar1S15S19P031N012N013N054(0)='1' AND  A( 4)='0' AND E( 3)='1' AND A( 2)='0' )then
          cVar2S15S19N011P056P015nsss(0) <='1';
          else
          cVar2S15S19N011P056P015nsss(0) <='0';
          end if;
        if(cVar1S16S19N031P036P007P037(0)='1' AND  A(14)='0' AND D( 3)='0' AND E( 2)='0' )then
          cVar2S16S19P010P054P060nsss(0) <='1';
          else
          cVar2S16S19P010P054P060nsss(0) <='0';
          end if;
        if(cVar1S17S19N031P036P007P037(0)='1' AND  A(14)='0' AND D( 3)='1' AND B( 2)='1' )then
          cVar2S17S19P010P054P033nsss(0) <='1';
          else
          cVar2S17S19P010P054P033nsss(0) <='0';
          end if;
        if(cVar1S18S19N031P036P007P037(0)='1' AND  A(14)='1' AND A(12)='0' AND A(16)='0' )then
          cVar2S18S19P010P014P006nsss(0) <='1';
          else
          cVar2S18S19P010P014P006nsss(0) <='0';
          end if;
        if(cVar1S19S19N031P036P007P037(0)='1' AND  A(14)='1' AND A(12)='1' AND E( 2)='1' )then
          cVar2S19S19P010P014P060nsss(0) <='1';
          else
          cVar2S19S19P010P014P060nsss(0) <='0';
          end if;
        if(cVar1S20S19N031P036P007P037(0)='1' AND  B( 1)='0' AND A( 5)='1' AND A(15)='0' )then
          cVar2S20S19P035P009P008nsss(0) <='1';
          else
          cVar2S20S19P035P009P008nsss(0) <='0';
          end if;
        if(cVar1S21S19N031P036P007P037(0)='1' AND  B( 1)='1' AND D(10)='1' )then
          cVar2S21S19P035P059nsss(0) <='1';
          else
          cVar2S21S19P035P059nsss(0) <='0';
          end if;
        if(cVar1S22S19N031P036P007P008(0)='1' AND  D(10)='0' AND A(14)='1' AND A( 5)='0' )then
          cVar2S22S19P059P010P009nsss(0) <='1';
          else
          cVar2S22S19P059P010P009nsss(0) <='0';
          end if;
        if(cVar1S23S19N031P036P007P008(0)='1' AND  B( 1)='1' AND A( 5)='0' )then
          cVar2S23S19P035P009nsss(0) <='1';
          else
          cVar2S23S19P035P009nsss(0) <='0';
          end if;
        if(cVar1S24S19N031P036P007P008(0)='1' AND  B( 1)='0' AND A(11)='1' AND A( 3)='0' )then
          cVar2S24S19N035P016P013nsss(0) <='1';
          else
          cVar2S24S19N035P016P013nsss(0) <='0';
          end if;
        if(cVar1S25S19N031N036P045P007(0)='1' AND  B(16)='1' )then
          cVar2S25S19P022nsss(0) <='1';
          else
          cVar2S25S19P022nsss(0) <='0';
          end if;
        if(cVar1S26S19N031N036P045P007(0)='1' AND  B(16)='0' AND B(15)='1' )then
          cVar2S26S19N022P024nsss(0) <='1';
          else
          cVar2S26S19N022P024nsss(0) <='0';
          end if;
        if(cVar1S27S19N031N036P045P007(0)='1' AND  B(16)='0' AND B(15)='0' AND A( 3)='0' )then
          cVar2S27S19N022N024P013nsss(0) <='1';
          else
          cVar2S27S19N022N024P013nsss(0) <='0';
          end if;
        if(cVar1S28S19N031N036P045N007(0)='1' AND  A(15)='1' AND A( 5)='1' )then
          cVar2S28S19P008P009nsss(0) <='1';
          else
          cVar2S28S19P008P009nsss(0) <='0';
          end if;
        if(cVar1S29S19N031N036P045N007(0)='1' AND  A(15)='1' AND A( 5)='0' AND D(14)='1' )then
          cVar2S29S19P008N009P043nsss(0) <='1';
          else
          cVar2S29S19P008N009P043nsss(0) <='0';
          end if;
        if(cVar1S30S19N031N036P045N007(0)='1' AND  A(15)='0' AND D( 0)='0' )then
          cVar2S30S19N008P066nsss(0) <='1';
          else
          cVar2S30S19N008P066nsss(0) <='0';
          end if;
        if(cVar1S31S19N031N036N045P053(0)='1' AND  D(12)='1' AND B(14)='1' AND A(13)='0' )then
          cVar2S31S19P051P026P012nsss(0) <='1';
          else
          cVar2S31S19P051P026P012nsss(0) <='0';
          end if;
        if(cVar1S32S19N031N036N045P053(0)='1' AND  D(12)='1' AND B(14)='0' AND D( 0)='0' )then
          cVar2S32S19P051N026P066nsss(0) <='1';
          else
          cVar2S32S19P051N026P066nsss(0) <='0';
          end if;
        if(cVar1S33S19N031N036N045P053(0)='1' AND  D(12)='0' AND B(13)='1' AND A( 0)='0' )then
          cVar2S33S19N051P028P019nsss(0) <='1';
          else
          cVar2S33S19N051P028P019nsss(0) <='0';
          end if;
        if(cVar1S34S19N031N036N045N053(0)='1' AND  D(15)='1' AND B(17)='1' )then
          cVar2S34S19P039P020nsss(0) <='1';
          else
          cVar2S34S19P039P020nsss(0) <='0';
          end if;
        if(cVar1S35S19N031N036N045N053(0)='1' AND  D(15)='1' AND B(17)='0' AND B(16)='1' )then
          cVar2S35S19P039N020P022nsss(0) <='1';
          else
          cVar2S35S19P039N020P022nsss(0) <='0';
          end if;
        if(cVar1S36S19N031N036N045N053(0)='1' AND  D(15)='0' AND B(12)='1' AND A( 4)='1' )then
          cVar2S36S19N039P030P011nsss(0) <='1';
          else
          cVar2S36S19N039P030P011nsss(0) <='0';
          end if;
        if(cVar1S0S20P032P031P016P013(0)='1' AND  A(16)='0' AND A( 0)='0' )then
          cVar2S0S20P006P019nsss(0) <='1';
          else
          cVar2S0S20P006P019nsss(0) <='0';
          end if;
        if(cVar1S1S20P032P031P016P013(0)='1' AND  A(16)='0' AND A( 0)='1' AND D(11)='0' )then
          cVar2S1S20P006P019P055nsss(0) <='1';
          else
          cVar2S1S20P006P019P055nsss(0) <='0';
          end if;
        if(cVar1S2S20P032P031P016P013(0)='1' AND  A(16)='1' AND A(10)='0' )then
          cVar2S2S20P006P018nsss(0) <='1';
          else
          cVar2S2S20P006P018nsss(0) <='0';
          end if;
        if(cVar1S3S20P032P031P016P013(0)='1' AND  A( 7)='0' AND A( 2)='0' )then
          cVar2S3S20P005P015nsss(0) <='1';
          else
          cVar2S3S20P005P015nsss(0) <='0';
          end if;
        if(cVar1S4S20P032P031P016P013(0)='1' AND  A( 7)='0' AND A( 2)='1' AND B( 0)='1' )then
          cVar2S4S20P005P015P037nsss(0) <='1';
          else
          cVar2S4S20P005P015P037nsss(0) <='0';
          end if;
        if(cVar1S5S20P032P031N016P018(0)='1' AND  A( 8)='0' AND E( 0)='0' AND A( 0)='0' )then
          cVar2S5S20P003P068P019nsss(0) <='1';
          else
          cVar2S5S20P003P068P019nsss(0) <='0';
          end if;
        if(cVar1S6S20P032P031N016P018(0)='1' AND  A( 8)='0' AND E( 0)='1' )then
          cVar2S6S20P003P068psss(0) <='1';
          else
          cVar2S6S20P003P068psss(0) <='0';
          end if;
        if(cVar1S7S20P032P031N016P018(0)='1' AND  A( 8)='1' AND D(10)='1' )then
          cVar2S7S20P003P059nsss(0) <='1';
          else
          cVar2S7S20P003P059nsss(0) <='0';
          end if;
        if(cVar1S8S20P032P031N016N018(0)='1' AND  A(12)='1' )then
          cVar2S8S20P014nsss(0) <='1';
          else
          cVar2S8S20P014nsss(0) <='0';
          end if;
        if(cVar1S9S20P032P031N016N018(0)='1' AND  A(12)='0' AND A( 0)='1' AND B( 1)='0' )then
          cVar2S9S20N014P019P035nsss(0) <='1';
          else
          cVar2S9S20N014P019P035nsss(0) <='0';
          end if;
        if(cVar1S10S20P032P031N016N018(0)='1' AND  A(12)='0' AND A( 0)='0' AND D( 3)='1' )then
          cVar2S10S20N014N019P054nsss(0) <='1';
          else
          cVar2S10S20N014N019P054nsss(0) <='0';
          end if;
        if(cVar1S11S20P032P031P003P018(0)='1' AND  A(12)='1' )then
          cVar2S11S20P014nsss(0) <='1';
          else
          cVar2S11S20P014nsss(0) <='0';
          end if;
        if(cVar1S12S20P032P031P003N018(0)='1' AND  D( 0)='0' AND A(14)='1' )then
          cVar2S12S20P066P010nsss(0) <='1';
          else
          cVar2S12S20P066P010nsss(0) <='0';
          end if;
        if(cVar1S13S20N032P036P024P047(0)='1' AND  A( 6)='1' )then
          cVar2S13S20P007nsss(0) <='1';
          else
          cVar2S13S20P007nsss(0) <='0';
          end if;
        if(cVar1S14S20N032P036P024P047(0)='1' AND  A( 6)='0' AND A( 5)='1' )then
          cVar2S14S20N007P009nsss(0) <='1';
          else
          cVar2S14S20N007P009nsss(0) <='0';
          end if;
        if(cVar1S15S20N032P036P024P047(0)='1' AND  A( 6)='0' AND A( 5)='0' AND E( 8)='1' )then
          cVar2S15S20N007N009P069nsss(0) <='1';
          else
          cVar2S15S20N007N009P069nsss(0) <='0';
          end if;
        if(cVar1S16S20N032P036P024N047(0)='1' AND  A(14)='0' AND D( 5)='1' )then
          cVar2S16S20P010P046nsss(0) <='1';
          else
          cVar2S16S20P010P046nsss(0) <='0';
          end if;
        if(cVar1S17S20N032P036P024N047(0)='1' AND  A(14)='0' AND D( 5)='0' AND E( 1)='1' )then
          cVar2S17S20P010N046P064nsss(0) <='1';
          else
          cVar2S17S20P010N046P064nsss(0) <='0';
          end if;
        if(cVar1S18S20N032P036P024N047(0)='1' AND  A(14)='1' AND B( 6)='1' )then
          cVar2S18S20P010P025nsss(0) <='1';
          else
          cVar2S18S20P010P025nsss(0) <='0';
          end if;
        if(cVar1S19S20N032P036N024P019(0)='1' AND  A( 2)='0' AND D(10)='0' )then
          cVar2S19S20P015P059nsss(0) <='1';
          else
          cVar2S19S20P015P059nsss(0) <='0';
          end if;
        if(cVar1S20S20N032P036N024P019(0)='1' AND  A( 2)='0' AND D(10)='1' AND B(10)='1' )then
          cVar2S20S20P015P059P034nsss(0) <='1';
          else
          cVar2S20S20P015P059P034nsss(0) <='0';
          end if;
        if(cVar1S21S20N032P036N024P019(0)='1' AND  A( 2)='1' AND E(10)='1' AND D( 0)='1' )then
          cVar2S21S20P015P061P066nsss(0) <='1';
          else
          cVar2S21S20P015P061P066nsss(0) <='0';
          end if;
        if(cVar1S22S20N032P036N024P019(0)='1' AND  A( 2)='1' AND E(10)='0' AND E( 2)='1' )then
          cVar2S22S20P015N061P060nsss(0) <='1';
          else
          cVar2S22S20P015N061P060nsss(0) <='0';
          end if;
        if(cVar1S23S20N032P036N024N019(0)='1' AND  A( 2)='1' AND E(10)='1' )then
          cVar2S23S20P015P061nsss(0) <='1';
          else
          cVar2S23S20P015P061nsss(0) <='0';
          end if;
        if(cVar1S24S20N032P036N024N019(0)='1' AND  A( 2)='1' AND E(10)='0' AND A(10)='0' )then
          cVar2S24S20P015N061P018nsss(0) <='1';
          else
          cVar2S24S20P015N061P018nsss(0) <='0';
          end if;
        if(cVar1S25S20N032P036N024N019(0)='1' AND  A( 2)='0' AND A(11)='1' AND E(10)='0' )then
          cVar2S25S20N015P016P061nsss(0) <='1';
          else
          cVar2S25S20N015P016P061nsss(0) <='0';
          end if;
        if(cVar1S26S20N032P036N024N019(0)='1' AND  A( 2)='0' AND A(11)='0' AND A(14)='1' )then
          cVar2S26S20N015N016P010nsss(0) <='1';
          else
          cVar2S26S20N015N016P010nsss(0) <='0';
          end if;
        if(cVar1S27S20N032P036P010P029(0)='1' AND  D( 4)='0' AND D( 6)='1' AND A( 3)='0' )then
          cVar2S27S20P050P042P013nsss(0) <='1';
          else
          cVar2S27S20P050P042P013nsss(0) <='0';
          end if;
        if(cVar1S28S20N032P036P010P029(0)='1' AND  D( 4)='0' AND D( 6)='0' AND B( 0)='1' )then
          cVar2S28S20P050N042P037nsss(0) <='1';
          else
          cVar2S28S20P050N042P037nsss(0) <='0';
          end if;
        if(cVar1S29S20N032P036P010P029(0)='1' AND  D( 4)='1' AND A(15)='1' AND D( 8)='0' )then
          cVar2S29S20P050P008P067nsss(0) <='1';
          else
          cVar2S29S20P050P008P067nsss(0) <='0';
          end if;
        if(cVar1S30S20N032P036P010P029(0)='1' AND  E( 1)='0' AND D( 8)='0' AND B(10)='0' )then
          cVar2S30S20P064P067P034nsss(0) <='1';
          else
          cVar2S30S20P064P067P034nsss(0) <='0';
          end if;
        if(cVar1S31S20N032P036P010P029(0)='1' AND  E( 1)='0' AND D( 8)='1' AND A( 4)='1' )then
          cVar2S31S20P064P067P011nsss(0) <='1';
          else
          cVar2S31S20P064P067P011nsss(0) <='0';
          end if;
        if(cVar1S32S20N032P036P010P055(0)='1' AND  B(12)='1' )then
          cVar2S32S20P030nsss(0) <='1';
          else
          cVar2S32S20P030nsss(0) <='0';
          end if;
        if(cVar1S33S20N032P036P010P055(0)='1' AND  B(12)='0' AND D( 8)='0' )then
          cVar2S33S20N030P067nsss(0) <='1';
          else
          cVar2S33S20N030P067nsss(0) <='0';
          end if;
        if(cVar1S34S20N032P036P010N055(0)='1' AND  D( 4)='1' AND A( 3)='0' )then
          cVar2S34S20P050P013nsss(0) <='1';
          else
          cVar2S34S20P050P013nsss(0) <='0';
          end if;
        if(cVar1S0S21P024P047P066P063(0)='1' AND  B( 1)='0' AND D( 5)='0' )then
          cVar2S0S21P035P046nsss(0) <='1';
          else
          cVar2S0S21P035P046nsss(0) <='0';
          end if;
        if(cVar1S1S21P024P047P066P063(0)='1' AND  B( 1)='0' AND D( 5)='1' AND E(13)='1' )then
          cVar2S1S21P035P046P049nsss(0) <='1';
          else
          cVar2S1S21P035P046P049nsss(0) <='0';
          end if;
        if(cVar1S2S21P024P047P066P063(0)='1' AND  B( 1)='1' )then
          cVar2S2S21P035psss(0) <='1';
          else
          cVar2S2S21P035psss(0) <='0';
          end if;
        if(cVar1S4S21P024P047P066N007(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S4S21P016P018nsss(0) <='1';
          else
          cVar2S4S21P016P018nsss(0) <='0';
          end if;
        if(cVar1S5S21P024N047P010P043(0)='1' AND  A(11)='1' )then
          cVar2S5S21P016nsss(0) <='1';
          else
          cVar2S5S21P016nsss(0) <='0';
          end if;
        if(cVar1S6S21P024N047P010P043(0)='1' AND  A(11)='0' AND E( 6)='0' )then
          cVar2S6S21N016P044nsss(0) <='1';
          else
          cVar2S6S21N016P044nsss(0) <='0';
          end if;
        if(cVar1S7S21P024N047P010N043(0)='1' AND  D( 5)='1' AND B( 9)='0' )then
          cVar2S7S21P046P036nsss(0) <='1';
          else
          cVar2S7S21P046P036nsss(0) <='0';
          end if;
        if(cVar1S8S21P024N047P010N043(0)='1' AND  D( 5)='0' AND E(10)='1' AND B( 2)='1' )then
          cVar2S8S21N046P061P033nsss(0) <='1';
          else
          cVar2S8S21N046P061P033nsss(0) <='0';
          end if;
        if(cVar1S9S21P024N047P010N043(0)='1' AND  D( 5)='0' AND E(10)='0' AND E( 6)='1' )then
          cVar2S9S21N046N061P044nsss(0) <='1';
          else
          cVar2S9S21N046N061P044nsss(0) <='0';
          end if;
        if(cVar1S11S21P024N047P010N032(0)='1' AND  B( 0)='1' AND A( 1)='1' )then
          cVar2S11S21P037P017nsss(0) <='1';
          else
          cVar2S11S21P037P017nsss(0) <='0';
          end if;
        if(cVar1S12S21N024P030P057P063(0)='1' AND  A( 4)='0' )then
          cVar2S12S21P011nsss(0) <='1';
          else
          cVar2S12S21P011nsss(0) <='0';
          end if;
        if(cVar1S13S21N024P030P057N063(0)='1' AND  A( 4)='1' AND A( 3)='0' )then
          cVar2S13S21P011P013nsss(0) <='1';
          else
          cVar2S13S21P011P013nsss(0) <='0';
          end if;
        if(cVar1S14S21N024P030P057N063(0)='1' AND  A( 4)='1' AND A( 3)='1' AND A(10)='1' )then
          cVar2S14S21P011P013P018nsss(0) <='1';
          else
          cVar2S14S21P011P013P018nsss(0) <='0';
          end if;
        if(cVar1S15S21N024P030P057N063(0)='1' AND  A( 4)='0' AND D(11)='0' AND A( 3)='1' )then
          cVar2S15S21N011P055P013nsss(0) <='1';
          else
          cVar2S15S21N011P055P013nsss(0) <='0';
          end if;
        if(cVar1S16S21N024P030P057N063(0)='1' AND  A( 4)='0' AND D(11)='1' )then
          cVar2S16S21N011P055psss(0) <='1';
          else
          cVar2S16S21N011P055psss(0) <='0';
          end if;
        if(cVar1S17S21N024P030N057P029(0)='1' AND  A(12)='0' AND E( 7)='1' )then
          cVar2S17S21P014P040nsss(0) <='1';
          else
          cVar2S17S21P014P040nsss(0) <='0';
          end if;
        if(cVar1S18S21N024P030N057P029(0)='1' AND  A(12)='0' AND E( 7)='0' AND E( 3)='1' )then
          cVar2S18S21P014N040P056nsss(0) <='1';
          else
          cVar2S18S21P014N040P056nsss(0) <='0';
          end if;
        if(cVar1S19S21N024P030N057P029(0)='1' AND  A(12)='1' AND A(13)='1' AND A( 4)='0' )then
          cVar2S19S21P014P012P011nsss(0) <='1';
          else
          cVar2S19S21P014P012P011nsss(0) <='0';
          end if;
        if(cVar1S20S21N024P030N057P029(0)='1' AND  A(12)='1' AND A(13)='0' AND E( 2)='1' )then
          cVar2S20S21P014N012P060nsss(0) <='1';
          else
          cVar2S20S21P014N012P060nsss(0) <='0';
          end if;
        if(cVar1S21S21N024N030P031P019(0)='1' AND  B(10)='0' AND A(13)='1' AND A(15)='0' )then
          cVar2S21S21P034P012P008nsss(0) <='1';
          else
          cVar2S21S21P034P012P008nsss(0) <='0';
          end if;
        if(cVar1S22S21N024N030P031P019(0)='1' AND  B(10)='0' AND A(13)='0' AND D(10)='0' )then
          cVar2S22S21P034N012P059nsss(0) <='1';
          else
          cVar2S22S21P034N012P059nsss(0) <='0';
          end if;
        if(cVar1S23S21N024N030P031P019(0)='1' AND  B(10)='1' AND A( 6)='0' AND B( 2)='1' )then
          cVar2S23S21P034P007P033nsss(0) <='1';
          else
          cVar2S23S21P034P007P033nsss(0) <='0';
          end if;
        if(cVar1S24S21N024N030P031P019(0)='1' AND  D( 8)='0' AND E( 3)='1' )then
          cVar2S24S21P067P056nsss(0) <='1';
          else
          cVar2S24S21P067P056nsss(0) <='0';
          end if;
        if(cVar1S25S21N024N030P031P019(0)='1' AND  D( 8)='0' AND E( 3)='0' AND E(11)='1' )then
          cVar2S25S21P067N056P057nsss(0) <='1';
          else
          cVar2S25S21P067N056P057nsss(0) <='0';
          end if;
        if(cVar1S26S21N024N030P031P019(0)='1' AND  D( 8)='1' AND E( 0)='1' AND A(13)='0' )then
          cVar2S26S21P067P068P012nsss(0) <='1';
          else
          cVar2S26S21P067P068P012nsss(0) <='0';
          end if;
        if(cVar1S27S21N024N030N031P055(0)='1' AND  A( 1)='1' AND A(12)='1' AND A(15)='0' )then
          cVar2S27S21P017P014P008nsss(0) <='1';
          else
          cVar2S27S21P017P014P008nsss(0) <='0';
          end if;
        if(cVar1S28S21N024N030N031P055(0)='1' AND  A( 1)='1' AND A(12)='0' )then
          cVar2S28S21P017N014psss(0) <='1';
          else
          cVar2S28S21P017N014psss(0) <='0';
          end if;
        if(cVar1S29S21N024N030N031P055(0)='1' AND  A( 1)='0' AND A( 2)='1' AND E(10)='1' )then
          cVar2S29S21N017P015P061nsss(0) <='1';
          else
          cVar2S29S21N017P015P061nsss(0) <='0';
          end if;
        if(cVar1S30S21N024N030N031P055(0)='1' AND  A( 1)='0' AND A( 2)='0' AND D( 8)='1' )then
          cVar2S30S21N017N015P067nsss(0) <='1';
          else
          cVar2S30S21N017N015P067nsss(0) <='0';
          end if;
        if(cVar1S31S21N024N030N031P055(0)='1' AND  B(13)='1' AND D( 1)='0' AND A(15)='0' )then
          cVar2S31S21P028P062P008nsss(0) <='1';
          else
          cVar2S31S21P028P062P008nsss(0) <='0';
          end if;
        if(cVar1S32S21N024N030N031P055(0)='1' AND  B(13)='1' AND D( 1)='1' AND A( 4)='1' )then
          cVar2S32S21P028P062P011nsss(0) <='1';
          else
          cVar2S32S21P028P062P011nsss(0) <='0';
          end if;
        if(cVar1S33S21N024N030N031P055(0)='1' AND  B(13)='0' AND B( 4)='1' AND A( 0)='0' )then
          cVar2S33S21N028P029P019nsss(0) <='1';
          else
          cVar2S33S21N028P029P019nsss(0) <='0';
          end if;
        if(cVar1S1S22P024P047P066P068(0)='1' AND  E(14)='0' AND A( 0)='0' )then
          cVar2S1S22P045P019nsss(0) <='1';
          else
          cVar2S1S22P045P019nsss(0) <='0';
          end if;
        if(cVar1S2S22P024P047P066P068(0)='1' AND  E(14)='0' AND A( 0)='1' AND B( 0)='1' )then
          cVar2S2S22P045P019P037nsss(0) <='1';
          else
          cVar2S2S22P045P019P037nsss(0) <='0';
          end if;
        if(cVar1S3S22P024N047P010P001(0)='1' AND  D(14)='1' )then
          cVar2S3S22P043nsss(0) <='1';
          else
          cVar2S3S22P043nsss(0) <='0';
          end if;
        if(cVar1S4S22P024N047P010P001(0)='1' AND  D(14)='0' AND D( 5)='1' AND B( 9)='0' )then
          cVar2S4S22N043P046P036nsss(0) <='1';
          else
          cVar2S4S22N043P046P036nsss(0) <='0';
          end if;
        if(cVar1S5S22P024N047P010P001(0)='1' AND  D(14)='0' AND D( 5)='0' AND A( 1)='1' )then
          cVar2S5S22N043N046P017nsss(0) <='1';
          else
          cVar2S5S22N043N046P017nsss(0) <='0';
          end if;
        if(cVar1S7S22P024N047P010N032(0)='1' AND  B( 0)='1' AND A( 2)='1' )then
          cVar2S7S22P037P015nsss(0) <='1';
          else
          cVar2S7S22P037P015nsss(0) <='0';
          end if;
        if(cVar1S8S22N024P067P017P022(0)='1' AND  A( 6)='1' )then
          cVar2S8S22P007nsss(0) <='1';
          else
          cVar2S8S22P007nsss(0) <='0';
          end if;
        if(cVar1S9S22N024P067P017P022(0)='1' AND  A( 6)='0' AND A( 7)='1' )then
          cVar2S9S22N007P005nsss(0) <='1';
          else
          cVar2S9S22N007P005nsss(0) <='0';
          end if;
        if(cVar1S10S22N024P067P017P022(0)='1' AND  A( 6)='0' AND A( 7)='0' AND D( 6)='1' )then
          cVar2S10S22N007N005P042nsss(0) <='1';
          else
          cVar2S10S22N007N005P042nsss(0) <='0';
          end if;
        if(cVar1S11S22N024P067P017N022(0)='1' AND  B( 9)='1' AND E( 8)='0' )then
          cVar2S11S22P036P069nsss(0) <='1';
          else
          cVar2S11S22P036P069nsss(0) <='0';
          end if;
        if(cVar1S12S22N024P067P017N022(0)='1' AND  B( 9)='0' )then
          cVar2S12S22N036psss(0) <='1';
          else
          cVar2S12S22N036psss(0) <='0';
          end if;
        if(cVar1S13S22N024P067P017P014(0)='1' AND  D( 0)='0' AND A(14)='0' )then
          cVar2S13S22P066P010nsss(0) <='1';
          else
          cVar2S13S22P066P010nsss(0) <='0';
          end if;
        if(cVar1S14S22N024P067P017P014(0)='1' AND  D( 0)='1' AND B( 0)='1' AND D(11)='0' )then
          cVar2S14S22P066P037P055nsss(0) <='1';
          else
          cVar2S14S22P066P037P055nsss(0) <='0';
          end if;
        if(cVar1S15S22N024P067P017N014(0)='1' AND  B( 3)='1' AND A(13)='1' AND D( 1)='0' )then
          cVar2S15S22P031P012P062nsss(0) <='1';
          else
          cVar2S15S22P031P012P062nsss(0) <='0';
          end if;
        if(cVar1S16S22N024P067P017N014(0)='1' AND  B( 3)='1' AND A(13)='0' AND D( 9)='1' )then
          cVar2S16S22P031N012P063nsss(0) <='1';
          else
          cVar2S16S22P031N012P063nsss(0) <='0';
          end if;
        if(cVar1S17S22N024P067P017N014(0)='1' AND  B( 3)='0' AND E( 8)='1' AND D( 9)='1' )then
          cVar2S17S22N031P069P063nsss(0) <='1';
          else
          cVar2S17S22N031P069P063nsss(0) <='0';
          end if;
        if(cVar1S18S22N024P067P017N014(0)='1' AND  B( 3)='0' AND E( 8)='0' AND B(12)='1' )then
          cVar2S18S22N031N069P030nsss(0) <='1';
          else
          cVar2S18S22N031N069P030nsss(0) <='0';
          end if;
        if(cVar1S19S22N024P067P060P064(0)='1' AND  B( 9)='1' AND B( 0)='0' )then
          cVar2S19S22P036P037nsss(0) <='1';
          else
          cVar2S19S22P036P037nsss(0) <='0';
          end if;
        if(cVar1S20S22N024P067P060P064(0)='1' AND  B( 9)='1' AND B( 0)='1' AND D( 2)='1' )then
          cVar2S20S22P036P037P058nsss(0) <='1';
          else
          cVar2S20S22P036P037P058nsss(0) <='0';
          end if;
        if(cVar1S21S22N024P067P060P064(0)='1' AND  B( 9)='0' AND A( 0)='0' AND D( 1)='0' )then
          cVar2S21S22N036P019P062nsss(0) <='1';
          else
          cVar2S21S22N036P019P062nsss(0) <='0';
          end if;
        if(cVar1S22S22N024P067P060P064(0)='1' AND  B( 9)='0' AND A( 0)='1' AND D( 2)='0' )then
          cVar2S22S22N036P019P058nsss(0) <='1';
          else
          cVar2S22S22N036P019P058nsss(0) <='0';
          end if;
        if(cVar1S23S22N024P067P060P064(0)='1' AND  A( 8)='1' )then
          cVar2S23S22P003nsss(0) <='1';
          else
          cVar2S23S22P003nsss(0) <='0';
          end if;
        if(cVar1S24S22N024P067P060P064(0)='1' AND  A( 8)='0' AND B( 2)='0' AND A(12)='1' )then
          cVar2S24S22N003P033P014nsss(0) <='1';
          else
          cVar2S24S22N003P033P014nsss(0) <='0';
          end if;
        if(cVar1S25S22N024P067N060P064(0)='1' AND  A( 1)='0' AND D( 5)='0' AND E( 0)='0' )then
          cVar2S25S22P017P046P068nsss(0) <='1';
          else
          cVar2S25S22P017P046P068nsss(0) <='0';
          end if;
        if(cVar1S26S22N024P067N060P064(0)='1' AND  A( 1)='1' AND B( 9)='0' AND A(10)='0' )then
          cVar2S26S22P017P036P018nsss(0) <='1';
          else
          cVar2S26S22P017P036P018nsss(0) <='0';
          end if;
        if(cVar1S27S22N024P067N060P064(0)='1' AND  A( 1)='1' AND B( 9)='1' AND A(12)='1' )then
          cVar2S27S22P017P036P014nsss(0) <='1';
          else
          cVar2S27S22P017P036P014nsss(0) <='0';
          end if;
        if(cVar1S28S22N024P067N060N064(0)='1' AND  D( 1)='0' AND A(10)='1' AND D(11)='1' )then
          cVar2S28S22P062P018P055nsss(0) <='1';
          else
          cVar2S28S22P062P018P055nsss(0) <='0';
          end if;
        if(cVar1S29S22N024P067N060N064(0)='1' AND  D( 1)='0' AND A(10)='0' AND B( 7)='1' )then
          cVar2S29S22P062N018P023nsss(0) <='1';
          else
          cVar2S29S22P062N018P023nsss(0) <='0';
          end if;
        if(cVar1S30S22N024P067N060N064(0)='1' AND  D( 1)='1' AND A( 0)='1' AND A(11)='1' )then
          cVar2S30S22P062P019P016nsss(0) <='1';
          else
          cVar2S30S22P062P019P016nsss(0) <='0';
          end if;
        if(cVar1S2S23P024P047P066N007(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S2S23P016P018nsss(0) <='1';
          else
          cVar2S2S23P016P018nsss(0) <='0';
          end if;
        if(cVar1S3S23P024P047P066N007(0)='1' AND  A(11)='0' AND A(10)='0' AND A(16)='1' )then
          cVar2S3S23P016N018P006nsss(0) <='1';
          else
          cVar2S3S23P016N018P006nsss(0) <='0';
          end if;
        if(cVar1S4S23P024N047P010P049(0)='1' AND  A(18)='0' AND E(10)='1' )then
          cVar2S4S23P002P061nsss(0) <='1';
          else
          cVar2S4S23P002P061nsss(0) <='0';
          end if;
        if(cVar1S5S23P024N047P010P049(0)='1' AND  A(18)='0' AND E(10)='0' AND D(10)='0' )then
          cVar2S5S23P002N061P059nsss(0) <='1';
          else
          cVar2S5S23P002N061P059nsss(0) <='0';
          end if;
        if(cVar1S6S23P024N047P010P049(0)='1' AND  A(18)='1' AND A(13)='0' AND A(10)='0' )then
          cVar2S6S23P002P012P018nsss(0) <='1';
          else
          cVar2S6S23P002P012P018nsss(0) <='0';
          end if;
        if(cVar1S7S23P024N047P010P018(0)='1' AND  A( 4)='1' )then
          cVar2S7S23P011nsss(0) <='1';
          else
          cVar2S7S23P011nsss(0) <='0';
          end if;
        if(cVar1S8S23N024P069P047P007(0)='1' AND  B(17)='0' AND E( 7)='1' AND B( 8)='1' )then
          cVar2S8S23P020P040P021nsss(0) <='1';
          else
          cVar2S8S23P020P040P021nsss(0) <='0';
          end if;
        if(cVar1S9S23N024P069P047P007(0)='1' AND  B(17)='0' AND E( 7)='0' )then
          cVar2S9S23P020N040psss(0) <='1';
          else
          cVar2S9S23P020N040psss(0) <='0';
          end if;
        if(cVar1S10S23N024P069P047P007(0)='1' AND  B(17)='1' AND A(11)='0' AND E( 0)='1' )then
          cVar2S10S23P020P016P068nsss(0) <='1';
          else
          cVar2S10S23P020P016P068nsss(0) <='0';
          end if;
        if(cVar1S11S23N024P069P047P007(0)='1' AND  E( 6)='0' AND E( 4)='1' )then
          cVar2S11S23P044P052nsss(0) <='1';
          else
          cVar2S11S23P044P052nsss(0) <='0';
          end if;
        if(cVar1S12S23N024P069P047P063(0)='1' AND  B(14)='1' )then
          cVar2S12S23P026nsss(0) <='1';
          else
          cVar2S12S23P026nsss(0) <='0';
          end if;
        if(cVar1S13S23N024P069P047P063(0)='1' AND  B(14)='0' AND A(12)='1' )then
          cVar2S13S23N026P014nsss(0) <='1';
          else
          cVar2S13S23N026P014nsss(0) <='0';
          end if;
        if(cVar1S14S23N024P069P047P063(0)='1' AND  B(14)='0' AND A(12)='0' AND A( 0)='0' )then
          cVar2S14S23N026N014P019nsss(0) <='1';
          else
          cVar2S14S23N026N014P019nsss(0) <='0';
          end if;
        if(cVar1S16S23N024N069P022N043(0)='1' AND  A(17)='1' )then
          cVar2S16S23P004nsss(0) <='1';
          else
          cVar2S16S23P004nsss(0) <='0';
          end if;
        if(cVar1S17S23N024N069P022N043(0)='1' AND  A(17)='0' AND A( 8)='0' AND D(15)='1' )then
          cVar2S17S23N004P003P039nsss(0) <='1';
          else
          cVar2S17S23N004P003P039nsss(0) <='0';
          end if;
        if(cVar1S18S23N024N069N022P036(0)='1' AND  A( 5)='0' AND D(13)='0' AND B( 0)='0' )then
          cVar2S18S23P009P047P037nsss(0) <='1';
          else
          cVar2S18S23P009P047P037nsss(0) <='0';
          end if;
        if(cVar1S19S23N024N069N022P036(0)='1' AND  A( 5)='0' AND D(13)='1' AND A( 0)='0' )then
          cVar2S19S23P009P047P019nsss(0) <='1';
          else
          cVar2S19S23P009P047P019nsss(0) <='0';
          end if;
        if(cVar1S20S23N024N069N022N036(0)='1' AND  B( 5)='1' AND A(19)='0' AND B( 6)='0' )then
          cVar2S20S23P027P000P025nsss(0) <='1';
          else
          cVar2S20S23P027P000P025nsss(0) <='0';
          end if;
        if(cVar1S21S23N024N069N022N036(0)='1' AND  B( 5)='0' AND A( 1)='1' AND D(11)='0' )then
          cVar2S21S23N027P017P055nsss(0) <='1';
          else
          cVar2S21S23N027P017P055nsss(0) <='0';
          end if;
        if(cVar1S22S23N024N069N022N036(0)='1' AND  B( 5)='0' AND A( 1)='0' AND B( 6)='1' )then
          cVar2S22S23N027N017P025nsss(0) <='1';
          else
          cVar2S22S23N027N017P025nsss(0) <='0';
          end if;
        if(cVar1S0S24P024P047P066P060(0)='1' AND  D( 5)='0' )then
          cVar2S0S24P046nsss(0) <='1';
          else
          cVar2S0S24P046nsss(0) <='0';
          end if;
        if(cVar1S1S24P024P047P066P060(0)='1' AND  D( 5)='1' AND E(13)='1' )then
          cVar2S1S24P046P049nsss(0) <='1';
          else
          cVar2S1S24P046P049nsss(0) <='0';
          end if;
        if(cVar1S4S24P024P047P066N069(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S4S24P016P018nsss(0) <='1';
          else
          cVar2S4S24P016P018nsss(0) <='0';
          end if;
        if(cVar1S5S24P024P047P066N069(0)='1' AND  A(11)='0' AND A(10)='0' AND A( 0)='1' )then
          cVar2S5S24P016N018P019nsss(0) <='1';
          else
          cVar2S5S24P016N018P019nsss(0) <='0';
          end if;
        if(cVar1S6S24P024N047P010P064(0)='1' AND  E(14)='1' )then
          cVar2S6S24P045nsss(0) <='1';
          else
          cVar2S6S24P045nsss(0) <='0';
          end if;
        if(cVar1S7S24P024N047P010P064(0)='1' AND  E(14)='0' AND B( 0)='1' AND E( 0)='0' )then
          cVar2S7S24N045P037P068nsss(0) <='1';
          else
          cVar2S7S24N045P037P068nsss(0) <='0';
          end if;
        if(cVar1S8S24P024N047P010P064(0)='1' AND  E(14)='0' AND B( 0)='0' AND A( 0)='1' )then
          cVar2S8S24N045N037P019nsss(0) <='1';
          else
          cVar2S8S24N045N037P019nsss(0) <='0';
          end if;
        if(cVar1S9S24P024N047P010N064(0)='1' AND  D(10)='1' AND A( 2)='1' )then
          cVar2S9S24P059P015nsss(0) <='1';
          else
          cVar2S9S24P059P015nsss(0) <='0';
          end if;
        if(cVar1S10S24P024N047P010N064(0)='1' AND  D(10)='1' AND A( 2)='0' AND B(11)='1' )then
          cVar2S10S24P059N015P032nsss(0) <='1';
          else
          cVar2S10S24P059N015P032nsss(0) <='0';
          end if;
        if(cVar1S11S24P024N047P010N064(0)='1' AND  D(10)='0' AND A(16)='1' AND E( 0)='0' )then
          cVar2S11S24N059P006P068nsss(0) <='1';
          else
          cVar2S11S24N059P006P068nsss(0) <='0';
          end if;
        if(cVar1S13S24P024N047P010N025(0)='1' AND  A(10)='0' AND A( 4)='1' )then
          cVar2S13S24P018P011nsss(0) <='1';
          else
          cVar2S13S24P018P011nsss(0) <='0';
          end if;
        if(cVar1S15S24N024P040N021P037(0)='1' AND  D( 1)='1' )then
          cVar2S15S24P062nsss(0) <='1';
          else
          cVar2S15S24P062nsss(0) <='0';
          end if;
        if(cVar1S16S24N024P040N021P037(0)='1' AND  D( 1)='0' AND A(13)='1' )then
          cVar2S16S24N062P012nsss(0) <='1';
          else
          cVar2S16S24N062P012nsss(0) <='0';
          end if;
        if(cVar1S17S24N024P040N021P037(0)='1' AND  D( 1)='0' AND A(13)='0' AND A( 0)='1' )then
          cVar2S17S24N062N012P019nsss(0) <='1';
          else
          cVar2S17S24N062N012P019nsss(0) <='0';
          end if;
        if(cVar1S18S24N024P040N021N037(0)='1' AND  B( 7)='1' AND A(10)='1' )then
          cVar2S18S24P023P018nsss(0) <='1';
          else
          cVar2S18S24P023P018nsss(0) <='0';
          end if;
        if(cVar1S19S24N024P040N021N037(0)='1' AND  B( 7)='1' AND A(10)='0' AND A(17)='1' )then
          cVar2S19S24P023N018P004nsss(0) <='1';
          else
          cVar2S19S24P023N018P004nsss(0) <='0';
          end if;
        if(cVar1S20S24N024P040N021N037(0)='1' AND  B( 7)='0' AND A(18)='1' AND D( 7)='1' )then
          cVar2S20S24N023P002P038nsss(0) <='1';
          else
          cVar2S20S24N023P002P038nsss(0) <='0';
          end if;
        if(cVar1S21S24N024N040P002P039(0)='1' AND  B(17)='1' AND A( 7)='1' )then
          cVar2S21S24P020P005nsss(0) <='1';
          else
          cVar2S21S24P020P005nsss(0) <='0';
          end if;
        if(cVar1S22S24N024N040P002P039(0)='1' AND  B(17)='1' AND A( 7)='0' AND E(15)='1' )then
          cVar2S22S24P020N005P041nsss(0) <='1';
          else
          cVar2S22S24P020N005P041nsss(0) <='0';
          end if;
        if(cVar1S23S24N024N040P002P039(0)='1' AND  B(17)='0' AND E(15)='1' )then
          cVar2S23S24N020P041nsss(0) <='1';
          else
          cVar2S23S24N020P041nsss(0) <='0';
          end if;
        if(cVar1S24S24N024N040P002N039(0)='1' AND  B( 8)='0' AND B(14)='1' AND E(13)='1' )then
          cVar2S24S24P021P026P049nsss(0) <='1';
          else
          cVar2S24S24P021P026P049nsss(0) <='0';
          end if;
        if(cVar1S25S24N024N040P002N039(0)='1' AND  B( 8)='1' AND A( 0)='1' AND B( 9)='1' )then
          cVar2S25S24P021P019P036nsss(0) <='1';
          else
          cVar2S25S24P021P019P036nsss(0) <='0';
          end if;
        if(cVar1S26S24N024N040P002P053(0)='1' AND  A( 0)='0' )then
          cVar2S26S24P019nsss(0) <='1';
          else
          cVar2S26S24P019nsss(0) <='0';
          end if;
        if(cVar1S27S24N024N040P002N053(0)='1' AND  E( 5)='1' AND A( 3)='0' AND D( 5)='1' )then
          cVar2S27S24P048P013P046nsss(0) <='1';
          else
          cVar2S27S24P048P013P046nsss(0) <='0';
          end if;
        if(cVar1S28S24N024N040P002N053(0)='1' AND  E( 5)='0' AND E( 8)='0' AND B(17)='1' )then
          cVar2S28S24N048N069P020nsss(0) <='1';
          else
          cVar2S28S24N048N069P020nsss(0) <='0';
          end if;
        if(cVar1S0S25P001P031P012P062(0)='1' AND  A( 1)='1' AND E( 3)='1' )then
          cVar2S0S25P017P056nsss(0) <='1';
          else
          cVar2S0S25P017P056nsss(0) <='0';
          end if;
        if(cVar1S1S25P001P031P012P062(0)='1' AND  A( 1)='1' AND E( 3)='0' AND E( 2)='1' )then
          cVar2S1S25P017N056P060nsss(0) <='1';
          else
          cVar2S1S25P017N056P060nsss(0) <='0';
          end if;
        if(cVar1S2S25P001P031P012P062(0)='1' AND  A( 1)='0' AND A(10)='1' )then
          cVar2S2S25N017P018nsss(0) <='1';
          else
          cVar2S2S25N017P018nsss(0) <='0';
          end if;
        if(cVar1S3S25P001P031P012P062(0)='1' AND  A( 1)='0' AND A(10)='0' AND A(15)='0' )then
          cVar2S3S25N017N018P008nsss(0) <='1';
          else
          cVar2S3S25N017N018P008nsss(0) <='0';
          end if;
        if(cVar1S4S25P001P031P012P062(0)='1' AND  A(10)='0' AND E( 1)='1' AND D( 9)='0' )then
          cVar2S4S25P018P064P063nsss(0) <='1';
          else
          cVar2S4S25P018P064P063nsss(0) <='0';
          end if;
        if(cVar1S5S25P001P031N012P013(0)='1' AND  D( 1)='1' AND D(10)='0' )then
          cVar2S5S25P062P059nsss(0) <='1';
          else
          cVar2S5S25P062P059nsss(0) <='0';
          end if;
        if(cVar1S6S25P001P031N012P013(0)='1' AND  D( 1)='0' AND A( 7)='0' AND B(12)='0' )then
          cVar2S6S25N062P005P030nsss(0) <='1';
          else
          cVar2S6S25N062P005P030nsss(0) <='0';
          end if;
        if(cVar1S7S25P001P031N012N013(0)='1' AND  D( 3)='1' AND A(12)='1' )then
          cVar2S7S25P054P014nsss(0) <='1';
          else
          cVar2S7S25P054P014nsss(0) <='0';
          end if;
        if(cVar1S8S25P001P031N012N013(0)='1' AND  D( 3)='1' AND A(12)='0' AND B(10)='0' )then
          cVar2S8S25P054N014P034nsss(0) <='1';
          else
          cVar2S8S25P054N014P034nsss(0) <='0';
          end if;
        if(cVar1S9S25P001N031P030P063(0)='1' AND  D(11)='1' )then
          cVar2S9S25P055nsss(0) <='1';
          else
          cVar2S9S25P055nsss(0) <='0';
          end if;
        if(cVar1S10S25P001N031P030P063(0)='1' AND  D(11)='0' AND A(12)='0' )then
          cVar2S10S25N055P014nsss(0) <='1';
          else
          cVar2S10S25N055P014nsss(0) <='0';
          end if;
        if(cVar1S11S25P001N031P030N063(0)='1' AND  D(10)='1' AND A( 3)='1' )then
          cVar2S11S25P059P013nsss(0) <='1';
          else
          cVar2S11S25P059P013nsss(0) <='0';
          end if;
        if(cVar1S12S25P001N031P030N063(0)='1' AND  D(10)='1' AND A( 3)='0' AND E( 1)='0' )then
          cVar2S12S25P059N013P064nsss(0) <='1';
          else
          cVar2S12S25P059N013P064nsss(0) <='0';
          end if;
        if(cVar1S13S25P001N031P030N063(0)='1' AND  D(10)='0' AND A( 3)='0' )then
          cVar2S13S25N059P013nsss(0) <='1';
          else
          cVar2S13S25N059P013nsss(0) <='0';
          end if;
        if(cVar1S14S25P001N031P030N063(0)='1' AND  D(10)='0' AND A( 3)='1' AND E( 8)='1' )then
          cVar2S14S25N059P013P069nsss(0) <='1';
          else
          cVar2S14S25N059P013P069nsss(0) <='0';
          end if;
        if(cVar1S15S25P001N031N030P055(0)='1' AND  A( 2)='1' AND E( 0)='1' )then
          cVar2S15S25P015P068nsss(0) <='1';
          else
          cVar2S15S25P015P068nsss(0) <='0';
          end if;
        if(cVar1S16S25P001N031N030P055(0)='1' AND  A( 2)='1' AND E( 0)='0' AND B( 1)='1' )then
          cVar2S16S25P015N068P035nsss(0) <='1';
          else
          cVar2S16S25P015N068P035nsss(0) <='0';
          end if;
        if(cVar1S17S25P001N031N030P055(0)='1' AND  A( 2)='0' AND E(13)='1' AND D( 9)='0' )then
          cVar2S17S25N015P049P063nsss(0) <='1';
          else
          cVar2S17S25N015P049P063nsss(0) <='0';
          end if;
        if(cVar1S18S25P001N031N030P055(0)='1' AND  A( 2)='0' AND E(13)='0' AND D(13)='0' )then
          cVar2S18S25N015N049P047nsss(0) <='1';
          else
          cVar2S18S25N015N049P047nsss(0) <='0';
          end if;
        if(cVar1S19S25P001N031N030P055(0)='1' AND  B(13)='1' AND D(12)='0' )then
          cVar2S19S25P028P051nsss(0) <='1';
          else
          cVar2S19S25P028P051nsss(0) <='0';
          end if;
        if(cVar1S20S25P001N031N030P055(0)='1' AND  B(13)='1' AND D(12)='1' AND A(14)='1' )then
          cVar2S20S25P028P051P010nsss(0) <='1';
          else
          cVar2S20S25P028P051P010nsss(0) <='0';
          end if;
        if(cVar1S21S25P001N031N030P055(0)='1' AND  B(13)='0' AND B(11)='1' AND E(10)='0' )then
          cVar2S21S25N028P032P061nsss(0) <='1';
          else
          cVar2S21S25N028P032P061nsss(0) <='0';
          end if;
        if(cVar1S22S25P001N031N030P055(0)='1' AND  B(13)='0' AND B(11)='0' AND B( 4)='1' )then
          cVar2S22S25N028N032P029nsss(0) <='1';
          else
          cVar2S22S25N028N032P029nsss(0) <='0';
          end if;
        if(cVar1S23S25P001P023P067P012(0)='1' AND  B( 9)='0' )then
          cVar2S23S25P036nsss(0) <='1';
          else
          cVar2S23S25P036nsss(0) <='0';
          end if;
        if(cVar1S24S25P001P023P067N012(0)='1' AND  A(11)='0' AND A( 0)='1' AND A( 1)='0' )then
          cVar2S24S25P016P019P017nsss(0) <='1';
          else
          cVar2S24S25P016P019P017nsss(0) <='0';
          end if;
        if(cVar1S25S25P001P023P067N012(0)='1' AND  A(11)='0' AND A( 0)='0' AND E( 0)='1' )then
          cVar2S25S25P016N019P068nsss(0) <='1';
          else
          cVar2S25S25P016N019P068nsss(0) <='0';
          end if;
        if(cVar1S27S25P001P023N067N041(0)='1' AND  B( 4)='1' AND A( 0)='0' )then
          cVar2S27S25P029P019nsss(0) <='1';
          else
          cVar2S27S25P029P019nsss(0) <='0';
          end if;
        if(cVar1S28S25P001P023N067N041(0)='1' AND  B( 4)='0' AND B( 0)='1' AND A( 3)='0' )then
          cVar2S28S25N029P037P013nsss(0) <='1';
          else
          cVar2S28S25N029P037P013nsss(0) <='0';
          end if;
        if(cVar1S29S25P001P023N067N041(0)='1' AND  B( 4)='0' AND B( 0)='0' AND B(12)='1' )then
          cVar2S29S25N029N037P030nsss(0) <='1';
          else
          cVar2S29S25N029N037P030nsss(0) <='0';
          end if;
        if(cVar1S0S26P015P017P034P058(0)='1' AND  B(13)='0' AND D(12)='0' AND A(19)='0' )then
          cVar2S0S26P028P051P000nsss(0) <='1';
          else
          cVar2S0S26P028P051P000nsss(0) <='0';
          end if;
        if(cVar1S1S26P015P017P034P058(0)='1' AND  E( 8)='1' )then
          cVar2S1S26P069nsss(0) <='1';
          else
          cVar2S1S26P069nsss(0) <='0';
          end if;
        if(cVar1S2S26P015P017P034P058(0)='1' AND  E( 8)='0' AND D( 9)='0' AND A( 3)='0' )then
          cVar2S2S26N069P063P013nsss(0) <='1';
          else
          cVar2S2S26N069P063P013nsss(0) <='0';
          end if;
        if(cVar1S3S26P015P017N034P033(0)='1' AND  D(13)='0' AND E(14)='0' )then
          cVar2S3S26P047P045nsss(0) <='1';
          else
          cVar2S3S26P047P045nsss(0) <='0';
          end if;
        if(cVar1S4S26P015P017N034N033(0)='1' AND  E( 9)='1' AND B( 1)='1' AND A( 3)='0' )then
          cVar2S4S26P065P035P013nsss(0) <='1';
          else
          cVar2S4S26P065P035P013nsss(0) <='0';
          end if;
        if(cVar1S5S26P015P017N034N033(0)='1' AND  E( 9)='1' AND B( 1)='0' AND B( 9)='1' )then
          cVar2S5S26P065N035P036nsss(0) <='1';
          else
          cVar2S5S26P065N035P036nsss(0) <='0';
          end if;
        if(cVar1S6S26P015P017N034N033(0)='1' AND  E( 9)='0' AND D( 8)='1' AND A( 0)='1' )then
          cVar2S6S26N065P067P019nsss(0) <='1';
          else
          cVar2S6S26N065P067P019nsss(0) <='0';
          end if;
        if(cVar1S7S26P015P017N034N033(0)='1' AND  E( 9)='0' AND D( 8)='0' AND E(11)='1' )then
          cVar2S7S26N065N067P057nsss(0) <='1';
          else
          cVar2S7S26N065N067P057nsss(0) <='0';
          end if;
        if(cVar1S8S26P015P017P006P001(0)='1' AND  A(18)='0' AND E( 9)='1' AND A(11)='1' )then
          cVar2S8S26P002P065P016nsss(0) <='1';
          else
          cVar2S8S26P002P065P016nsss(0) <='0';
          end if;
        if(cVar1S9S26P015P017P006P001(0)='1' AND  A(18)='0' AND E( 9)='0' AND B( 2)='1' )then
          cVar2S9S26P002N065P033nsss(0) <='1';
          else
          cVar2S9S26P002N065P033nsss(0) <='0';
          end if;
        if(cVar1S10S26P015P017P006P001(0)='1' AND  A(18)='1' AND A(13)='1' AND A( 4)='1' )then
          cVar2S10S26P002P012P011nsss(0) <='1';
          else
          cVar2S10S26P002P012P011nsss(0) <='0';
          end if;
        if(cVar1S11S26P015P017P006P001(0)='1' AND  B(10)='0' AND B( 9)='0' AND A(10)='1' )then
          cVar2S11S26P034P036P018nsss(0) <='1';
          else
          cVar2S11S26P034P036P018nsss(0) <='0';
          end if;
        if(cVar1S12S26P015P017P006P062(0)='1' AND  B( 0)='1' )then
          cVar2S12S26P037nsss(0) <='1';
          else
          cVar2S12S26P037nsss(0) <='0';
          end if;
        if(cVar1S13S26P015P017P006P062(0)='1' AND  B( 0)='0' AND B( 1)='0' )then
          cVar2S13S26N037P035nsss(0) <='1';
          else
          cVar2S13S26N037P035nsss(0) <='0';
          end if;
        if(cVar1S14S26P015P017P006N062(0)='1' AND  B(15)='1' )then
          cVar2S14S26P024nsss(0) <='1';
          else
          cVar2S14S26P024nsss(0) <='0';
          end if;
        if(cVar1S15S26P015P017P006N062(0)='1' AND  B(15)='0' AND B( 6)='1' )then
          cVar2S15S26N024P025nsss(0) <='1';
          else
          cVar2S15S26N024P025nsss(0) <='0';
          end if;
        if(cVar1S16S26P015P017P006N062(0)='1' AND  B(15)='0' AND B( 6)='0' AND B( 3)='1' )then
          cVar2S16S26N024N025P031nsss(0) <='1';
          else
          cVar2S16S26N024N025P031nsss(0) <='0';
          end if;
        if(cVar1S17S26N015P031P012P017(0)='1' AND  A(11)='0' )then
          cVar2S17S26P016nsss(0) <='1';
          else
          cVar2S17S26P016nsss(0) <='0';
          end if;
        if(cVar1S18S26N015P031P012P017(0)='1' AND  A(11)='1' AND A(12)='0' AND A( 0)='0' )then
          cVar2S18S26P016P014P019nsss(0) <='1';
          else
          cVar2S18S26P016P014P019nsss(0) <='0';
          end if;
        if(cVar1S19S26N015P031P012N017(0)='1' AND  A(10)='1' AND E( 8)='1' )then
          cVar2S19S26P018P069nsss(0) <='1';
          else
          cVar2S19S26P018P069nsss(0) <='0';
          end if;
        if(cVar1S20S26N015P031P012N017(0)='1' AND  A(10)='1' AND E( 8)='0' AND E( 3)='1' )then
          cVar2S20S26P018N069P056nsss(0) <='1';
          else
          cVar2S20S26P018N069P056nsss(0) <='0';
          end if;
        if(cVar1S21S26N015P031P012N017(0)='1' AND  A(10)='0' AND A(14)='0' )then
          cVar2S21S26N018P010nsss(0) <='1';
          else
          cVar2S21S26N018P010nsss(0) <='0';
          end if;
        if(cVar1S22S26N015P031N012P014(0)='1' AND  E(11)='1' )then
          cVar2S22S26P057nsss(0) <='1';
          else
          cVar2S22S26P057nsss(0) <='0';
          end if;
        if(cVar1S23S26N015P031N012P014(0)='1' AND  E(11)='0' AND E( 3)='1' AND A(10)='0' )then
          cVar2S23S26N057P056P018nsss(0) <='1';
          else
          cVar2S23S26N057P056P018nsss(0) <='0';
          end if;
        if(cVar1S24S26N015P031N012P014(0)='1' AND  E(11)='0' AND E( 3)='0' AND D( 2)='1' )then
          cVar2S24S26N057N056P058nsss(0) <='1';
          else
          cVar2S24S26N057N056P058nsss(0) <='0';
          end if;
        if(cVar1S25S26N015P031N012N014(0)='1' AND  E( 1)='1' AND D( 3)='0' AND E(11)='1' )then
          cVar2S25S26P064P054P057nsss(0) <='1';
          else
          cVar2S25S26P064P054P057nsss(0) <='0';
          end if;
        if(cVar1S26S26N015P031N012N014(0)='1' AND  E( 1)='1' AND D( 3)='1' AND B( 0)='0' )then
          cVar2S26S26P064P054P037nsss(0) <='1';
          else
          cVar2S26S26P064P054P037nsss(0) <='0';
          end if;
        if(cVar1S27S26N015P031N012N014(0)='1' AND  E( 1)='0' AND A(14)='1' AND D( 8)='0' )then
          cVar2S27S26N064P010P067nsss(0) <='1';
          else
          cVar2S27S26N064P010P067nsss(0) <='0';
          end if;
        if(cVar1S28S26N015P031N012N014(0)='1' AND  E( 1)='0' AND A(14)='0' AND B( 5)='1' )then
          cVar2S28S26N064N010P027nsss(0) <='1';
          else
          cVar2S28S26N064N010P027nsss(0) <='0';
          end if;
        if(cVar1S29S26N015N031P030P059(0)='1' AND  A( 3)='1' )then
          cVar2S29S26P013nsss(0) <='1';
          else
          cVar2S29S26P013nsss(0) <='0';
          end if;
        if(cVar1S30S26N015N031P030P059(0)='1' AND  A( 3)='0' AND A(12)='1' AND A(13)='1' )then
          cVar2S30S26N013P014P012nsss(0) <='1';
          else
          cVar2S30S26N013P014P012nsss(0) <='0';
          end if;
        if(cVar1S31S26N015N031P030P059(0)='1' AND  A( 3)='0' AND A(12)='0' AND A( 4)='1' )then
          cVar2S31S26N013N014P011nsss(0) <='1';
          else
          cVar2S31S26N013N014P011nsss(0) <='0';
          end if;
        if(cVar1S32S26N015N031P030N059(0)='1' AND  D( 9)='1' AND D(11)='1' )then
          cVar2S32S26P063P055nsss(0) <='1';
          else
          cVar2S32S26P063P055nsss(0) <='0';
          end if;
        if(cVar1S33S26N015N031P030N059(0)='1' AND  D( 9)='1' AND D(11)='0' AND B( 9)='1' )then
          cVar2S33S26P063N055P036nsss(0) <='1';
          else
          cVar2S33S26P063N055P036nsss(0) <='0';
          end if;
        if(cVar1S34S26N015N031P030N059(0)='1' AND  D( 9)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar2S34S26N063P060P017nsss(0) <='1';
          else
          cVar2S34S26N063P060P017nsss(0) <='0';
          end if;
        if(cVar1S35S26N015N031N030P007(0)='1' AND  D(13)='1' AND B( 5)='0' )then
          cVar2S35S26P047P027nsss(0) <='1';
          else
          cVar2S35S26P047P027nsss(0) <='0';
          end if;
        if(cVar1S36S26N015N031N030P007(0)='1' AND  D(13)='0' AND D( 5)='1' AND B( 6)='1' )then
          cVar2S36S26N047P046P025nsss(0) <='1';
          else
          cVar2S36S26N047P046P025nsss(0) <='0';
          end if;
        if(cVar1S37S26N015N031N030P007(0)='1' AND  D(13)='0' AND D( 5)='0' AND B(16)='1' )then
          cVar2S37S26N047N046P022nsss(0) <='1';
          else
          cVar2S37S26N047N046P022nsss(0) <='0';
          end if;
        if(cVar1S38S26N015N031N030N007(0)='1' AND  B( 7)='1' AND D( 6)='1' AND D( 0)='0' )then
          cVar2S38S26P023P042P066nsss(0) <='1';
          else
          cVar2S38S26P023P042P066nsss(0) <='0';
          end if;
        if(cVar1S39S26N015N031N030N007(0)='1' AND  B( 7)='1' AND D( 6)='0' AND E( 1)='1' )then
          cVar2S39S26P023N042P064nsss(0) <='1';
          else
          cVar2S39S26P023N042P064nsss(0) <='0';
          end if;
        if(cVar1S40S26N015N031N030N007(0)='1' AND  B( 7)='0' AND E(12)='1' AND E( 0)='1' )then
          cVar2S40S26N023P053P068nsss(0) <='1';
          else
          cVar2S40S26N023P053P068nsss(0) <='0';
          end if;
        if(cVar1S1S27P002P022P043N007(0)='1' AND  A( 8)='1' )then
          cVar2S1S27P003nsss(0) <='1';
          else
          cVar2S1S27P003nsss(0) <='0';
          end if;
        if(cVar1S2S27P002P022P043N007(0)='1' AND  A( 8)='0' AND A( 7)='1' )then
          cVar2S2S27N003P005nsss(0) <='1';
          else
          cVar2S2S27N003P005nsss(0) <='0';
          end if;
        if(cVar1S3S27P002P022P043N007(0)='1' AND  A( 8)='0' AND A( 7)='0' AND A(17)='1' )then
          cVar2S3S27N003N005P004nsss(0) <='1';
          else
          cVar2S3S27N003N005P004nsss(0) <='0';
          end if;
        if(cVar1S4S27P002P022N043P042(0)='1' AND  A(10)='0' AND A(17)='1' )then
          cVar2S4S27P018P004nsss(0) <='1';
          else
          cVar2S4S27P018P004nsss(0) <='0';
          end if;
        if(cVar1S5S27P002P022N043P042(0)='1' AND  A(10)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S5S27P018N004P006nsss(0) <='1';
          else
          cVar2S5S27P018N004P006nsss(0) <='0';
          end if;
        if(cVar1S6S27P002P022N043N042(0)='1' AND  A( 8)='0' AND D(15)='1' )then
          cVar2S6S27P003P039nsss(0) <='1';
          else
          cVar2S6S27P003P039nsss(0) <='0';
          end if;
        if(cVar1S7S27P002P022N043N042(0)='1' AND  A( 8)='0' AND D(15)='0' AND E(11)='1' )then
          cVar2S7S27P003N039P057nsss(0) <='1';
          else
          cVar2S7S27P003N039P057nsss(0) <='0';
          end if;
        if(cVar1S8S27P002N022P027P026(0)='1' AND  A( 1)='1' AND A(16)='0' )then
          cVar2S8S27P017P006nsss(0) <='1';
          else
          cVar2S8S27P017P006nsss(0) <='0';
          end if;
        if(cVar1S9S27P002N022P027P026(0)='1' AND  A( 1)='0' AND A(15)='1' )then
          cVar2S9S27N017P008nsss(0) <='1';
          else
          cVar2S9S27N017P008nsss(0) <='0';
          end if;
        if(cVar1S10S27P002N022P027P026(0)='1' AND  A( 1)='0' AND A(15)='0' AND A(16)='1' )then
          cVar2S10S27N017N008P006nsss(0) <='1';
          else
          cVar2S10S27N017N008P006nsss(0) <='0';
          end if;
        if(cVar1S11S27P002N022P027P026(0)='1' AND  A(14)='0' AND E( 8)='0' AND A( 2)='0' )then
          cVar2S11S27P010P069P015nsss(0) <='1';
          else
          cVar2S11S27P010P069P015nsss(0) <='0';
          end if;
        if(cVar1S12S27P002N022N027P032(0)='1' AND  B( 1)='0' AND E( 2)='0' AND B( 2)='0' )then
          cVar2S12S27P035P060P033nsss(0) <='1';
          else
          cVar2S12S27P035P060P033nsss(0) <='0';
          end if;
        if(cVar1S13S27P002N022N027P032(0)='1' AND  B( 1)='0' AND E( 2)='1' AND B( 2)='1' )then
          cVar2S13S27P035P060P033nsss(0) <='1';
          else
          cVar2S13S27P035P060P033nsss(0) <='0';
          end if;
        if(cVar1S14S27P002N022N027P032(0)='1' AND  B( 1)='1' AND A(11)='1' AND E( 2)='1' )then
          cVar2S14S27P035P016P060nsss(0) <='1';
          else
          cVar2S14S27P035P016P060nsss(0) <='0';
          end if;
        if(cVar1S15S27P002N022N027N032(0)='1' AND  D(10)='0' AND E(10)='0' )then
          cVar2S15S27P059P061nsss(0) <='1';
          else
          cVar2S15S27P059P061nsss(0) <='0';
          end if;
        if(cVar1S16S27P002N022N027N032(0)='1' AND  D(10)='0' AND E(10)='1' AND A( 3)='1' )then
          cVar2S16S27P059P061P013nsss(0) <='1';
          else
          cVar2S16S27P059P061P013nsss(0) <='0';
          end if;
        if(cVar1S17S27P002N022N027N032(0)='1' AND  D(10)='1' AND E(10)='1' AND E( 1)='0' )then
          cVar2S17S27P059P061P064nsss(0) <='1';
          else
          cVar2S17S27P059P061P064nsss(0) <='0';
          end if;
        if(cVar1S18S27P002N022N027N032(0)='1' AND  D(10)='1' AND E(10)='0' AND A( 3)='1' )then
          cVar2S18S27P059N061P013nsss(0) <='1';
          else
          cVar2S18S27P059N061P013nsss(0) <='0';
          end if;
        if(cVar1S21S27P002N040P050P048(0)='1' AND  A( 0)='1' )then
          cVar2S21S27P019nsss(0) <='1';
          else
          cVar2S21S27P019nsss(0) <='0';
          end if;
        if(cVar1S22S27P002N040P050N048(0)='1' AND  E(12)='1' AND A( 0)='0' )then
          cVar2S22S27P053P019nsss(0) <='1';
          else
          cVar2S22S27P053P019nsss(0) <='0';
          end if;
        if(cVar1S23S27P002N040P050N048(0)='1' AND  E(12)='0' AND E( 8)='1' AND A(14)='0' )then
          cVar2S23S27N053P069P010nsss(0) <='1';
          else
          cVar2S23S27N053P069P010nsss(0) <='0';
          end if;
        if(cVar1S0S28P032P002P016P049(0)='1' AND  B( 9)='0' )then
          cVar2S0S28P036nsss(0) <='1';
          else
          cVar2S0S28P036nsss(0) <='0';
          end if;
        if(cVar1S1S28P032P002P016P049(0)='1' AND  B( 9)='1' AND E( 8)='0' AND D( 9)='1' )then
          cVar2S1S28P036P069P063nsss(0) <='1';
          else
          cVar2S1S28P036P069P063nsss(0) <='0';
          end if;
        if(cVar1S2S28P032P002N016P063(0)='1' AND  D(10)='1' AND D( 2)='0' AND E( 8)='0' )then
          cVar2S2S28P059P058P069nsss(0) <='1';
          else
          cVar2S2S28P059P058P069nsss(0) <='0';
          end if;
        if(cVar1S3S28P032P002N016P063(0)='1' AND  D(10)='1' AND D( 2)='1' AND A(13)='1' )then
          cVar2S3S28P059P058P012nsss(0) <='1';
          else
          cVar2S3S28P059P058P012nsss(0) <='0';
          end if;
        if(cVar1S4S28P032P002N016P063(0)='1' AND  D(10)='0' AND D( 2)='1' )then
          cVar2S4S28N059P058nsss(0) <='1';
          else
          cVar2S4S28N059P058nsss(0) <='0';
          end if;
        if(cVar1S5S28P032P002N016N063(0)='1' AND  B(10)='0' AND A(14)='1' AND D(10)='1' )then
          cVar2S5S28P034P010P059nsss(0) <='1';
          else
          cVar2S5S28P034P010P059nsss(0) <='0';
          end if;
        if(cVar1S6S28P032P002N016N063(0)='1' AND  B(10)='0' AND A(14)='0' )then
          cVar2S6S28P034N010psss(0) <='1';
          else
          cVar2S6S28P034N010psss(0) <='0';
          end if;
        if(cVar1S7S28P032P002N016N063(0)='1' AND  B(10)='1' AND E( 1)='1' )then
          cVar2S7S28P034P064nsss(0) <='1';
          else
          cVar2S7S28P034P064nsss(0) <='0';
          end if;
        if(cVar1S8S28P032P002N016N063(0)='1' AND  B(10)='1' AND E( 1)='0' AND A( 1)='1' )then
          cVar2S8S28P034N064P017nsss(0) <='1';
          else
          cVar2S8S28P034N064P017nsss(0) <='0';
          end if;
        if(cVar1S10S28N032P027P026P000(0)='1' AND  A( 8)='0' )then
          cVar2S10S28P003nsss(0) <='1';
          else
          cVar2S10S28P003nsss(0) <='0';
          end if;
        if(cVar1S11S28N032P027P026P000(0)='1' AND  A( 8)='1' AND A(10)='0' AND A(11)='1' )then
          cVar2S11S28P003P018P016nsss(0) <='1';
          else
          cVar2S11S28P003P018P016nsss(0) <='0';
          end if;
        if(cVar1S12S28N032P027P026P000(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S12S28P016P018nsss(0) <='1';
          else
          cVar2S12S28P016P018nsss(0) <='0';
          end if;
        if(cVar1S13S28N032P027P026P036(0)='1' AND  A(14)='0' AND D( 0)='1' )then
          cVar2S13S28P010P066nsss(0) <='1';
          else
          cVar2S13S28P010P066nsss(0) <='0';
          end if;
        if(cVar1S14S28N032P027P026P036(0)='1' AND  A(14)='0' AND D( 0)='0' AND A(15)='1' )then
          cVar2S14S28P010N066P008nsss(0) <='1';
          else
          cVar2S14S28P010N066P008nsss(0) <='0';
          end if;
        if(cVar1S15S28N032N027P022P069(0)='1' AND  A(18)='0' AND A( 6)='1' AND A(13)='0' )then
          cVar2S15S28P002P007P012nsss(0) <='1';
          else
          cVar2S15S28P002P007P012nsss(0) <='0';
          end if;
        if(cVar1S16S28N032N027P022P069(0)='1' AND  A(18)='0' AND A( 6)='0' )then
          cVar2S16S28P002N007psss(0) <='1';
          else
          cVar2S16S28P002N007psss(0) <='0';
          end if;
        if(cVar1S17S28N032N027P022P069(0)='1' AND  A(18)='1' AND D(14)='1' )then
          cVar2S17S28P002P043nsss(0) <='1';
          else
          cVar2S17S28P002P043nsss(0) <='0';
          end if;
        if(cVar1S18S28N032N027P022P069(0)='1' AND  B( 1)='0' AND E( 0)='0' AND A( 2)='0' )then
          cVar2S18S28P035P068P015nsss(0) <='1';
          else
          cVar2S18S28P035P068P015nsss(0) <='0';
          end if;
        if(cVar1S19S28N032N027N022P030(0)='1' AND  B( 3)='0' AND E(11)='1' AND E( 3)='0' )then
          cVar2S19S28P031P057P056nsss(0) <='1';
          else
          cVar2S19S28P031P057P056nsss(0) <='0';
          end if;
        if(cVar1S20S28N032N027N022P030(0)='1' AND  B( 3)='1' AND A( 0)='1' AND B( 0)='0' )then
          cVar2S20S28P031P019P037nsss(0) <='1';
          else
          cVar2S20S28P031P019P037nsss(0) <='0';
          end if;
        if(cVar1S21S28N032N027N022P030(0)='1' AND  B( 3)='1' AND A( 0)='0' AND E( 9)='1' )then
          cVar2S21S28P031N019P065nsss(0) <='1';
          else
          cVar2S21S28P031N019P065nsss(0) <='0';
          end if;
        if(cVar1S22S28N032N027N022N030(0)='1' AND  D(15)='1' AND B(17)='1' )then
          cVar2S22S28P039P020nsss(0) <='1';
          else
          cVar2S22S28P039P020nsss(0) <='0';
          end if;
        if(cVar1S23S28N032N027N022N030(0)='1' AND  D(15)='1' AND B(17)='0' AND A( 7)='1' )then
          cVar2S23S28P039N020P005nsss(0) <='1';
          else
          cVar2S23S28P039N020P005nsss(0) <='0';
          end if;
        if(cVar1S24S28N032N027N022N030(0)='1' AND  D(15)='0' AND B( 6)='1' AND D( 5)='1' )then
          cVar2S24S28N039P025P046nsss(0) <='1';
          else
          cVar2S24S28N039P025P046nsss(0) <='0';
          end if;
        if(cVar1S1S29P040P021P035N002(0)='1' AND  A(17)='1' )then
          cVar2S1S29P004nsss(0) <='1';
          else
          cVar2S1S29P004nsss(0) <='0';
          end if;
        if(cVar1S2S29P040P021P035N002(0)='1' AND  A(17)='0' AND A( 0)='1' )then
          cVar2S2S29N004P019nsss(0) <='1';
          else
          cVar2S2S29N004P019nsss(0) <='0';
          end if;
        if(cVar1S3S29P040P021P035N002(0)='1' AND  A(17)='0' AND A( 0)='0' AND D( 7)='1' )then
          cVar2S3S29N004N019P038nsss(0) <='1';
          else
          cVar2S3S29N004N019P038nsss(0) <='0';
          end if;
        if(cVar1S4S29P040N021P037P005(0)='1' AND  D( 1)='1' )then
          cVar2S4S29P062nsss(0) <='1';
          else
          cVar2S4S29P062nsss(0) <='0';
          end if;
        if(cVar1S5S29P040N021P037P005(0)='1' AND  D( 1)='0' AND A(13)='1' )then
          cVar2S5S29N062P012nsss(0) <='1';
          else
          cVar2S5S29N062P012nsss(0) <='0';
          end if;
        if(cVar1S6S29P040N021P037P005(0)='1' AND  D( 1)='0' AND A(13)='0' AND E( 0)='1' )then
          cVar2S6S29N062N012P068nsss(0) <='1';
          else
          cVar2S6S29N062N012P068nsss(0) <='0';
          end if;
        if(cVar1S7S29P040N021N037P017(0)='1' AND  B( 9)='1' )then
          cVar2S7S29P036nsss(0) <='1';
          else
          cVar2S7S29P036nsss(0) <='0';
          end if;
        if(cVar1S8S29P040N021N037P017(0)='1' AND  B( 9)='0' AND A( 2)='1' )then
          cVar2S8S29N036P015nsss(0) <='1';
          else
          cVar2S8S29N036P015nsss(0) <='0';
          end if;
        if(cVar1S9S29P040N021N037N017(0)='1' AND  D( 5)='0' AND B( 1)='0' AND A(19)='1' )then
          cVar2S9S29P046P035P000nsss(0) <='1';
          else
          cVar2S9S29P046P035P000nsss(0) <='0';
          end if;
        if(cVar1S10S29N040P038P021P002(0)='1' AND  D( 9)='1' AND D( 1)='0' )then
          cVar2S10S29P063P062nsss(0) <='1';
          else
          cVar2S10S29P063P062nsss(0) <='0';
          end if;
        if(cVar1S11S29N040P038P021P002(0)='1' AND  D( 9)='1' AND D( 1)='1' AND A( 2)='1' )then
          cVar2S11S29P063P062P015nsss(0) <='1';
          else
          cVar2S11S29P063P062P015nsss(0) <='0';
          end if;
        if(cVar1S12S29N040P038P021P002(0)='1' AND  D( 9)='0' AND E( 1)='1' AND A( 0)='0' )then
          cVar2S12S29N063P064P019nsss(0) <='1';
          else
          cVar2S12S29N063P064P019nsss(0) <='0';
          end if;
        if(cVar1S13S29N040P038P021P002(0)='1' AND  D( 9)='0' AND E( 1)='0' AND E( 0)='1' )then
          cVar2S13S29N063N064P068nsss(0) <='1';
          else
          cVar2S13S29N063N064P068nsss(0) <='0';
          end if;
        if(cVar1S14S29N040P038P021P002(0)='1' AND  D( 4)='0' AND A(11)='0' AND A(19)='0' )then
          cVar2S14S29P050P016P000nsss(0) <='1';
          else
          cVar2S14S29P050P016P000nsss(0) <='0';
          end if;
        if(cVar1S15S29N040P038P021P002(0)='1' AND  D( 4)='0' AND A(11)='1' AND A( 8)='1' )then
          cVar2S15S29P050P016P003nsss(0) <='1';
          else
          cVar2S15S29P050P016P003nsss(0) <='0';
          end if;
        if(cVar1S16S29N040P038P021P002(0)='1' AND  D( 4)='1' AND A( 3)='1' )then
          cVar2S16S29P050P013nsss(0) <='1';
          else
          cVar2S16S29P050P013nsss(0) <='0';
          end if;
        if(cVar1S17S29N040P038P021P010(0)='1' AND  D(12)='0' AND A(13)='1' AND A( 4)='0' )then
          cVar2S17S29P051P012P011nsss(0) <='1';
          else
          cVar2S17S29P051P012P011nsss(0) <='0';
          end if;
        if(cVar1S18S29N040P038P021P010(0)='1' AND  A(12)='0' AND A( 8)='1' )then
          cVar2S18S29P014P003nsss(0) <='1';
          else
          cVar2S18S29P014P003nsss(0) <='0';
          end if;
        if(cVar1S20S29N040P038N026N059(0)='1' AND  A( 2)='0' AND B( 9)='0' AND D( 1)='1' )then
          cVar2S20S29P015P036P062nsss(0) <='1';
          else
          cVar2S20S29P015P036P062nsss(0) <='0';
          end if;
        if(cVar1S0S30P068P047P049P065(0)='1' AND  A( 5)='1' AND E( 5)='0' )then
          cVar2S0S30P009P048nsss(0) <='1';
          else
          cVar2S0S30P009P048nsss(0) <='0';
          end if;
        if(cVar1S1S30P068P047P049P065(0)='1' AND  A( 5)='0' AND D( 1)='0' )then
          cVar2S1S30N009P062nsss(0) <='1';
          else
          cVar2S1S30N009P062nsss(0) <='0';
          end if;
        if(cVar1S2S30P068P047P049P065(0)='1' AND  A( 5)='0' AND D( 1)='1' AND A( 6)='1' )then
          cVar2S2S30N009P062P007nsss(0) <='1';
          else
          cVar2S2S30N009P062P007nsss(0) <='0';
          end if;
        if(cVar1S3S30P068P047P049P065(0)='1' AND  A(16)='0' AND B(14)='1' )then
          cVar2S3S30P006P026nsss(0) <='1';
          else
          cVar2S3S30P006P026nsss(0) <='0';
          end if;
        if(cVar1S4S30P068P047P049P065(0)='1' AND  A(16)='0' AND B(14)='0' AND A(11)='0' )then
          cVar2S4S30P006N026P016nsss(0) <='1';
          else
          cVar2S4S30P006N026P016nsss(0) <='0';
          end if;
        if(cVar1S5S30P068P047N049P024(0)='1' AND  E(14)='1' )then
          cVar2S5S30P045nsss(0) <='1';
          else
          cVar2S5S30P045nsss(0) <='0';
          end if;
        if(cVar1S6S30P068P047N049N024(0)='1' AND  A( 5)='1' AND A(10)='1' )then
          cVar2S6S30P009P018nsss(0) <='1';
          else
          cVar2S6S30P009P018nsss(0) <='0';
          end if;
        if(cVar1S7S30P068P047N049N024(0)='1' AND  A( 5)='0' AND E( 5)='1' )then
          cVar2S7S30N009P048nsss(0) <='1';
          else
          cVar2S7S30N009P048nsss(0) <='0';
          end if;
        if(cVar1S8S30P068N047P052P066(0)='1' AND  B( 4)='1' AND D(12)='0' )then
          cVar2S8S30P029P051nsss(0) <='1';
          else
          cVar2S8S30P029P051nsss(0) <='0';
          end if;
        if(cVar1S9S30P068N047P052P066(0)='1' AND  B( 4)='1' AND D(12)='1' AND A( 4)='0' )then
          cVar2S9S30P029P051P011nsss(0) <='1';
          else
          cVar2S9S30P029P051P011nsss(0) <='0';
          end if;
        if(cVar1S10S30P068N047P052P066(0)='1' AND  B( 4)='0' AND B(13)='1' )then
          cVar2S10S30N029P028nsss(0) <='1';
          else
          cVar2S10S30N029P028nsss(0) <='0';
          end if;
        if(cVar1S11S30P068N047P052P066(0)='1' AND  B( 4)='0' AND B(13)='0' AND B(14)='1' )then
          cVar2S11S30N029N028P026nsss(0) <='1';
          else
          cVar2S11S30N029N028P026nsss(0) <='0';
          end if;
        if(cVar1S12S30P068N047P052P066(0)='1' AND  B( 9)='0' AND A( 2)='1' )then
          cVar2S12S30P036P015nsss(0) <='1';
          else
          cVar2S12S30P036P015nsss(0) <='0';
          end if;
        if(cVar1S13S30P068N047N052P036(0)='1' AND  B( 1)='0' AND A( 1)='1' )then
          cVar2S13S30P035P017nsss(0) <='1';
          else
          cVar2S13S30P035P017nsss(0) <='0';
          end if;
        if(cVar1S14S30P068N047N052P036(0)='1' AND  B( 1)='0' AND A( 1)='0' AND D( 9)='0' )then
          cVar2S14S30P035N017P063nsss(0) <='1';
          else
          cVar2S14S30P035N017P063nsss(0) <='0';
          end if;
        if(cVar1S15S30P068N047N052P036(0)='1' AND  B( 1)='1' AND E( 9)='1' AND A( 1)='0' )then
          cVar2S15S30P035P065P017nsss(0) <='1';
          else
          cVar2S15S30P035P065P017nsss(0) <='0';
          end if;
        if(cVar1S16S30P068N047N052N036(0)='1' AND  E(12)='1' AND E(13)='0' AND D( 0)='0' )then
          cVar2S16S30P053P049P066nsss(0) <='1';
          else
          cVar2S16S30P053P049P066nsss(0) <='0';
          end if;
        if(cVar1S17S30P068N047N052N036(0)='1' AND  E(12)='0' AND E(11)='1' )then
          cVar2S17S30N053P057nsss(0) <='1';
          else
          cVar2S17S30N053P057nsss(0) <='0';
          end if;
        if(cVar1S18S30P068N047N052N036(0)='1' AND  E(12)='0' AND E(11)='0' AND A( 4)='0' )then
          cVar2S18S30N053N057P011nsss(0) <='1';
          else
          cVar2S18S30N053N057P011nsss(0) <='0';
          end if;
        if(cVar1S19S30P068P055P019P047(0)='1' AND  E( 9)='0' AND D( 8)='0' AND D( 0)='1' )then
          cVar2S19S30P065P067P066nsss(0) <='1';
          else
          cVar2S19S30P065P067P066nsss(0) <='0';
          end if;
        if(cVar1S20S30P068P055P019P047(0)='1' AND  E( 9)='0' AND D( 8)='1' AND B( 0)='0' )then
          cVar2S20S30P065P067P037nsss(0) <='1';
          else
          cVar2S20S30P065P067P037nsss(0) <='0';
          end if;
        if(cVar1S21S30P068P055P019P047(0)='1' AND  E( 9)='1' AND B( 9)='1' )then
          cVar2S21S30P065P036nsss(0) <='1';
          else
          cVar2S21S30P065P036nsss(0) <='0';
          end if;
        if(cVar1S22S30P068P055P019P047(0)='1' AND  E( 9)='1' AND B( 9)='0' AND D( 1)='1' )then
          cVar2S22S30P065N036P062nsss(0) <='1';
          else
          cVar2S22S30P065N036P062nsss(0) <='0';
          end if;
        if(cVar1S23S30P068P055P019P047(0)='1' AND  B(15)='1' AND E(13)='0' )then
          cVar2S23S30P024P049nsss(0) <='1';
          else
          cVar2S23S30P024P049nsss(0) <='0';
          end if;
        if(cVar1S24S30P068P055P019P047(0)='1' AND  B(15)='1' AND E(13)='1' AND A(16)='0' )then
          cVar2S24S30P024P049P006nsss(0) <='1';
          else
          cVar2S24S30P024P049P006nsss(0) <='0';
          end if;
        if(cVar1S25S30P068P055P019P047(0)='1' AND  B(15)='0' AND A( 5)='1' )then
          cVar2S25S30N024P009nsss(0) <='1';
          else
          cVar2S25S30N024P009nsss(0) <='0';
          end if;
        if(cVar1S26S30P068P055N019P051(0)='1' AND  E( 1)='0' AND B(13)='0' AND A( 3)='0' )then
          cVar2S26S30P064P028P013nsss(0) <='1';
          else
          cVar2S26S30P064P028P013nsss(0) <='0';
          end if;
        if(cVar1S27S30P068P055N019P051(0)='1' AND  E( 1)='0' AND B(13)='1' AND A( 4)='1' )then
          cVar2S27S30P064P028P011nsss(0) <='1';
          else
          cVar2S27S30P064P028P011nsss(0) <='0';
          end if;
        if(cVar1S28S30P068P055N019N051(0)='1' AND  B( 0)='1' AND B( 4)='0' AND A( 1)='1' )then
          cVar2S28S30P037P029P017nsss(0) <='1';
          else
          cVar2S28S30P037P029P017nsss(0) <='0';
          end if;
        if(cVar1S29S30P068P055N019N051(0)='1' AND  B( 0)='0' AND E(10)='1' AND B( 1)='1' )then
          cVar2S29S30N037P061P035nsss(0) <='1';
          else
          cVar2S29S30N037P061P035nsss(0) <='0';
          end if;
        if(cVar1S30S30P068P055N019N051(0)='1' AND  B( 0)='0' AND E(10)='0' AND E(15)='1' )then
          cVar2S30S30N037N061P041nsss(0) <='1';
          else
          cVar2S30S30N037N061P041nsss(0) <='0';
          end if;
        if(cVar1S31S30P068P055P016P018(0)='1' AND  E(12)='0' )then
          cVar2S31S30P053nsss(0) <='1';
          else
          cVar2S31S30P053nsss(0) <='0';
          end if;
        if(cVar1S32S30P068P055P016P018(0)='1' AND  E( 8)='1' )then
          cVar2S32S30P069nsss(0) <='1';
          else
          cVar2S32S30P069nsss(0) <='0';
          end if;
        if(cVar1S33S30P068P055P016P018(0)='1' AND  E( 8)='0' AND A( 4)='1' )then
          cVar2S33S30N069P011nsss(0) <='1';
          else
          cVar2S33S30N069P011nsss(0) <='0';
          end if;
        if(cVar1S34S30P068P055N016P049(0)='1' AND  A(14)='1' AND A( 0)='0' )then
          cVar2S34S30P010P019nsss(0) <='1';
          else
          cVar2S34S30P010P019nsss(0) <='0';
          end if;
        if(cVar1S35S30P068P055N016P049(0)='1' AND  A(14)='1' AND A( 0)='1' AND E( 3)='1' )then
          cVar2S35S30P010P019P056nsss(0) <='1';
          else
          cVar2S35S30P010P019P056nsss(0) <='0';
          end if;
        if(cVar1S36S30P068P055N016P049(0)='1' AND  A(14)='0' AND A( 1)='1' AND A( 4)='1' )then
          cVar2S36S30N010P017P011nsss(0) <='1';
          else
          cVar2S36S30N010P017P011nsss(0) <='0';
          end if;
        if(cVar1S37S30P068P055N016P049(0)='1' AND  A(14)='0' AND A( 1)='0' AND A( 8)='1' )then
          cVar2S37S30N010N017P003nsss(0) <='1';
          else
          cVar2S37S30N010N017P003nsss(0) <='0';
          end if;
        if(cVar1S0S31P036P063P005P048(0)='1' AND  A( 0)='0' AND A( 1)='1' AND B(10)='0' )then
          cVar2S0S31P019P017P034nsss(0) <='1';
          else
          cVar2S0S31P019P017P034nsss(0) <='0';
          end if;
        if(cVar1S1S31P036P063P005P048(0)='1' AND  A( 0)='0' AND A( 1)='0' AND B(10)='1' )then
          cVar2S1S31P019N017P034nsss(0) <='1';
          else
          cVar2S1S31P019N017P034nsss(0) <='0';
          end if;
        if(cVar1S2S31P036P063P005P048(0)='1' AND  A( 0)='1' AND D(10)='0' AND D( 0)='0' )then
          cVar2S2S31P019P059P066nsss(0) <='1';
          else
          cVar2S2S31P019P059P066nsss(0) <='0';
          end if;
        if(cVar1S3S31P036P063P005P048(0)='1' AND  A( 0)='1' AND D(10)='1' AND E( 8)='0' )then
          cVar2S3S31P019P059P069nsss(0) <='1';
          else
          cVar2S3S31P019P059P069nsss(0) <='0';
          end if;
        if(cVar1S4S31P036P063P005P048(0)='1' AND  D( 0)='0' AND A( 0)='1' )then
          cVar2S4S31P066P019nsss(0) <='1';
          else
          cVar2S4S31P066P019nsss(0) <='0';
          end if;
        if(cVar1S5S31P036P063P005P048(0)='1' AND  D( 0)='0' AND A( 0)='0' AND A( 1)='1' )then
          cVar2S5S31P066N019P017nsss(0) <='1';
          else
          cVar2S5S31P066N019P017nsss(0) <='0';
          end if;
        if(cVar1S7S31P036P063P005N035(0)='1' AND  D( 8)='0' AND A( 1)='0' AND A( 2)='0' )then
          cVar2S7S31P067P017P015nsss(0) <='1';
          else
          cVar2S7S31P067P017P015nsss(0) <='0';
          end if;
        if(cVar1S8S31P036N063P016P064(0)='1' AND  A( 1)='0' AND A(10)='0' )then
          cVar2S8S31P017P018nsss(0) <='1';
          else
          cVar2S8S31P017P018nsss(0) <='0';
          end if;
        if(cVar1S9S31P036N063P016P064(0)='1' AND  A( 1)='0' AND A(10)='1' AND A(12)='1' )then
          cVar2S9S31P017P018P014nsss(0) <='1';
          else
          cVar2S9S31P017P018P014nsss(0) <='0';
          end if;
        if(cVar1S10S31P036N063P016P064(0)='1' AND  A( 1)='1' AND A( 2)='1' AND A(15)='0' )then
          cVar2S10S31P017P015P008nsss(0) <='1';
          else
          cVar2S10S31P017P015P008nsss(0) <='0';
          end if;
        if(cVar1S11S31P036N063P016P064(0)='1' AND  A( 1)='1' AND A( 2)='0' AND A(12)='1' )then
          cVar2S11S31P017N015P014nsss(0) <='1';
          else
          cVar2S11S31P017N015P014nsss(0) <='0';
          end if;
        if(cVar1S12S31P036N063P016N064(0)='1' AND  D( 1)='1' AND B( 1)='1' AND E( 8)='1' )then
          cVar2S12S31P062P035P069nsss(0) <='1';
          else
          cVar2S12S31P062P035P069nsss(0) <='0';
          end if;
        if(cVar1S13S31P036N063P016N064(0)='1' AND  D( 1)='1' AND B( 1)='0' AND A( 3)='0' )then
          cVar2S13S31P062N035P013nsss(0) <='1';
          else
          cVar2S13S31P062N035P013nsss(0) <='0';
          end if;
        if(cVar1S14S31P036N063P016N064(0)='1' AND  D( 1)='0' AND D(11)='1' AND D( 8)='1' )then
          cVar2S14S31N062P055P067nsss(0) <='1';
          else
          cVar2S14S31N062P055P067nsss(0) <='0';
          end if;
        if(cVar1S15S31P036N063P016N064(0)='1' AND  D( 1)='0' AND D(11)='0' AND E( 3)='1' )then
          cVar2S15S31N062N055P056nsss(0) <='1';
          else
          cVar2S15S31N062N055P056nsss(0) <='0';
          end if;
        if(cVar1S16S31P036N063N016P018(0)='1' AND  B(10)='0' AND A( 2)='0' AND D( 0)='0' )then
          cVar2S16S31P034P015P066nsss(0) <='1';
          else
          cVar2S16S31P034P015P066nsss(0) <='0';
          end if;
        if(cVar1S17S31P036N063N016P018(0)='1' AND  B(10)='0' AND A( 2)='1' AND B( 8)='1' )then
          cVar2S17S31P034P015P021nsss(0) <='1';
          else
          cVar2S17S31P034P015P021nsss(0) <='0';
          end if;
        if(cVar1S18S31P036N063N016P018(0)='1' AND  B(10)='1' AND E( 0)='1' AND B( 0)='0' )then
          cVar2S18S31P034P068P037nsss(0) <='1';
          else
          cVar2S18S31P034P068P037nsss(0) <='0';
          end if;
        if(cVar1S19S31P036N063N016P018(0)='1' AND  B(10)='1' AND E( 0)='0' AND A(13)='1' )then
          cVar2S19S31P034N068P012nsss(0) <='1';
          else
          cVar2S19S31P034N068P012nsss(0) <='0';
          end if;
        if(cVar1S20S31P036N063N016N018(0)='1' AND  D( 8)='1' AND E( 2)='1' AND B( 2)='1' )then
          cVar2S20S31P067P060P033nsss(0) <='1';
          else
          cVar2S20S31P067P060P033nsss(0) <='0';
          end if;
        if(cVar1S21S31P036N063N016N018(0)='1' AND  D( 8)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar2S21S31N067P058P033nsss(0) <='1';
          else
          cVar2S21S31N067P058P033nsss(0) <='0';
          end if;
        if(cVar1S22S31N036P052P068P048(0)='1' AND  D(12)='0' AND D( 0)='0' )then
          cVar2S22S31P051P066nsss(0) <='1';
          else
          cVar2S22S31P051P066nsss(0) <='0';
          end if;
        if(cVar1S23S31N036P052P068P048(0)='1' AND  D(12)='0' AND D( 0)='1' AND A( 0)='1' )then
          cVar2S23S31P051P066P019nsss(0) <='1';
          else
          cVar2S23S31P051P066P019nsss(0) <='0';
          end if;
        if(cVar1S24S31N036P052P068P048(0)='1' AND  D(12)='1' AND A( 0)='1' )then
          cVar2S24S31P051P019nsss(0) <='1';
          else
          cVar2S24S31P051P019nsss(0) <='0';
          end if;
        if(cVar1S25S31N036P052P068P048(0)='1' AND  D(12)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar2S25S31P051N019P064nsss(0) <='1';
          else
          cVar2S25S31P051N019P064nsss(0) <='0';
          end if;
        if(cVar1S26S31N036P052P068P048(0)='1' AND  D( 5)='1' )then
          cVar2S26S31P046nsss(0) <='1';
          else
          cVar2S26S31P046nsss(0) <='0';
          end if;
        if(cVar1S27S31N036P052P068P055(0)='1' AND  E( 3)='0' AND E( 8)='1' )then
          cVar2S27S31P056P069nsss(0) <='1';
          else
          cVar2S27S31P056P069nsss(0) <='0';
          end if;
        if(cVar1S28S31N036P052P068P055(0)='1' AND  E( 3)='0' AND E( 8)='0' AND B( 4)='1' )then
          cVar2S28S31P056N069P029nsss(0) <='1';
          else
          cVar2S28S31P056N069P029nsss(0) <='0';
          end if;
        if(cVar1S29S31N036N052P018P016(0)='1' AND  D( 8)='1' AND E(13)='1' )then
          cVar2S29S31P067P049nsss(0) <='1';
          else
          cVar2S29S31P067P049nsss(0) <='0';
          end if;
        if(cVar1S30S31N036N052P018P016(0)='1' AND  D( 8)='1' AND E(13)='0' AND D( 2)='0' )then
          cVar2S30S31P067N049P058nsss(0) <='1';
          else
          cVar2S30S31P067N049P058nsss(0) <='0';
          end if;
        if(cVar1S31S31N036N052P018P016(0)='1' AND  D( 8)='0' AND D( 0)='1' AND D(11)='0' )then
          cVar2S31S31N067P066P055nsss(0) <='1';
          else
          cVar2S31S31N067P066P055nsss(0) <='0';
          end if;
        if(cVar1S32S31N036N052P018P016(0)='1' AND  D( 8)='0' AND D( 0)='0' AND E( 1)='1' )then
          cVar2S32S31N067N066P064nsss(0) <='1';
          else
          cVar2S32S31N067N066P064nsss(0) <='0';
          end if;
        if(cVar1S33S31N036N052P018P016(0)='1' AND  B( 0)='1' AND A( 7)='0' AND D( 0)='1' )then
          cVar2S33S31P037P005P066nsss(0) <='1';
          else
          cVar2S33S31P037P005P066nsss(0) <='0';
          end if;
        if(cVar1S34S31N036N052P018P016(0)='1' AND  B( 0)='0' AND D(10)='1' AND B(11)='1' )then
          cVar2S34S31N037P059P032nsss(0) <='1';
          else
          cVar2S34S31N037P059P032nsss(0) <='0';
          end if;
        if(cVar1S35S31N036N052P018P016(0)='1' AND  B( 0)='0' AND D(10)='0' AND E(14)='1' )then
          cVar2S35S31N037N059P045nsss(0) <='1';
          else
          cVar2S35S31N037N059P045nsss(0) <='0';
          end if;
        if(cVar1S36S31N036N052N018P014(0)='1' AND  A( 2)='0' AND D(13)='1' )then
          cVar2S36S31P015P047nsss(0) <='1';
          else
          cVar2S36S31P015P047nsss(0) <='0';
          end if;
        if(cVar1S37S31N036N052N018P014(0)='1' AND  A( 2)='0' AND D(13)='0' AND A( 3)='1' )then
          cVar2S37S31P015N047P013nsss(0) <='1';
          else
          cVar2S37S31P015N047P013nsss(0) <='0';
          end if;
        if(cVar1S38S31N036N052N018P014(0)='1' AND  A( 2)='1' AND A(11)='0' AND E( 1)='1' )then
          cVar2S38S31P015P016P064nsss(0) <='1';
          else
          cVar2S38S31P015P016P064nsss(0) <='0';
          end if;
        if(cVar1S39S31N036N052N018P014(0)='1' AND  A( 2)='1' AND A(11)='1' AND A( 4)='1' )then
          cVar2S39S31P015P016P011nsss(0) <='1';
          else
          cVar2S39S31P015P016P011nsss(0) <='0';
          end if;
        if(cVar1S40S31N036N052N018N014(0)='1' AND  A(11)='1' AND E( 0)='1' AND B( 0)='1' )then
          cVar2S40S31P016P068P037nsss(0) <='1';
          else
          cVar2S40S31P016P068P037nsss(0) <='0';
          end if;
        if(cVar1S41S31N036N052N018N014(0)='1' AND  A(11)='1' AND E( 0)='0' AND B( 1)='1' )then
          cVar2S41S31P016N068P035nsss(0) <='1';
          else
          cVar2S41S31P016N068P035nsss(0) <='0';
          end if;
        if(cVar1S42S31N036N052N018N014(0)='1' AND  A(11)='0' AND E( 5)='1' AND D( 6)='0' )then
          cVar2S42S31N016P048P042nsss(0) <='1';
          else
          cVar2S42S31N016P048P042nsss(0) <='0';
          end if;
        if(cVar1S43S31N036N052N018N014(0)='1' AND  A(11)='0' AND E( 5)='0' AND D( 6)='1' )then
          cVar2S43S31N016N048P042nsss(0) <='1';
          else
          cVar2S43S31N016N048P042nsss(0) <='0';
          end if;
        if(cVar1S0S32P036P066P006P027(0)='1' AND  B( 7)='0' AND A( 0)='0' AND E( 5)='0' )then
          cVar2S0S32P023P019P048nsss(0) <='1';
          else
          cVar2S0S32P023P019P048nsss(0) <='0';
          end if;
        if(cVar1S1S32P036P066P006P027(0)='1' AND  B( 7)='0' AND A( 0)='1' AND E( 1)='0' )then
          cVar2S1S32P023P019P064nsss(0) <='1';
          else
          cVar2S1S32P023P019P064nsss(0) <='0';
          end if;
        if(cVar1S2S32P036P066P006P027(0)='1' AND  A( 5)='1' )then
          cVar2S2S32P009nsss(0) <='1';
          else
          cVar2S2S32P009nsss(0) <='0';
          end if;
        if(cVar1S3S32P036P066P006P059(0)='1' AND  A(10)='1' AND A(13)='0' )then
          cVar2S3S32P018P012nsss(0) <='1';
          else
          cVar2S3S32P018P012nsss(0) <='0';
          end if;
        if(cVar1S4S32P036N066P016P018(0)='1' AND  B(10)='0' AND D(13)='0' )then
          cVar2S4S32P034P047nsss(0) <='1';
          else
          cVar2S4S32P034P047nsss(0) <='0';
          end if;
        if(cVar1S5S32P036N066P016P018(0)='1' AND  B(10)='1' AND D(10)='1' )then
          cVar2S5S32P034P059nsss(0) <='1';
          else
          cVar2S5S32P034P059nsss(0) <='0';
          end if;
        if(cVar1S6S32P036N066P016P018(0)='1' AND  B(10)='1' AND D(10)='0' AND A( 0)='0' )then
          cVar2S6S32P034N059P019nsss(0) <='1';
          else
          cVar2S6S32P034N059P019nsss(0) <='0';
          end if;
        if(cVar1S7S32P036N066P016P018(0)='1' AND  A( 8)='1' AND A( 3)='0' )then
          cVar2S7S32P003P013nsss(0) <='1';
          else
          cVar2S7S32P003P013nsss(0) <='0';
          end if;
        if(cVar1S8S32P036N066P016P018(0)='1' AND  A( 8)='0' AND A(15)='1' AND A(13)='0' )then
          cVar2S8S32N003P008P012nsss(0) <='1';
          else
          cVar2S8S32N003P008P012nsss(0) <='0';
          end if;
        if(cVar1S9S32P036N066N016P068(0)='1' AND  A( 1)='1' AND D( 1)='0' AND B( 0)='0' )then
          cVar2S9S32P017P062P037nsss(0) <='1';
          else
          cVar2S9S32P017P062P037nsss(0) <='0';
          end if;
        if(cVar1S10S32P036N066N016P068(0)='1' AND  A( 1)='1' AND D( 1)='1' AND A(12)='1' )then
          cVar2S10S32P017P062P014nsss(0) <='1';
          else
          cVar2S10S32P017P062P014nsss(0) <='0';
          end if;
        if(cVar1S11S32P036N066N016P068(0)='1' AND  A( 1)='0' AND A(10)='1' AND D( 4)='0' )then
          cVar2S11S32N017P018P050nsss(0) <='1';
          else
          cVar2S11S32N017P018P050nsss(0) <='0';
          end if;
        if(cVar1S12S32P036N066N016P068(0)='1' AND  A( 0)='1' AND E( 8)='1' )then
          cVar2S12S32P019P069nsss(0) <='1';
          else
          cVar2S12S32P019P069nsss(0) <='0';
          end if;
        if(cVar1S13S32N036P060P048P063(0)='1' AND  B( 2)='1' AND E( 1)='0' AND A(17)='0' )then
          cVar2S13S32P033P064P004nsss(0) <='1';
          else
          cVar2S13S32P033P064P004nsss(0) <='0';
          end if;
        if(cVar1S14S32N036P060P048P063(0)='1' AND  B( 2)='1' AND E( 1)='1' AND D(10)='0' )then
          cVar2S14S32P033P064P059nsss(0) <='1';
          else
          cVar2S14S32P033P064P059nsss(0) <='0';
          end if;
        if(cVar1S15S32N036P060P048P063(0)='1' AND  B( 2)='0' AND D( 3)='0' AND A(13)='1' )then
          cVar2S15S32N033P054P012nsss(0) <='1';
          else
          cVar2S15S32N033P054P012nsss(0) <='0';
          end if;
        if(cVar1S16S32N036P060P048P063(0)='1' AND  B( 1)='1' AND B(11)='1' )then
          cVar2S16S32P035P032nsss(0) <='1';
          else
          cVar2S16S32P035P032nsss(0) <='0';
          end if;
        if(cVar1S17S32N036P060P048P063(0)='1' AND  B( 1)='1' AND B(11)='0' AND E( 9)='1' )then
          cVar2S17S32P035N032P065nsss(0) <='1';
          else
          cVar2S17S32P035N032P065nsss(0) <='0';
          end if;
        if(cVar1S18S32N036P060P048P063(0)='1' AND  B( 1)='0' AND A( 1)='1' AND B( 0)='1' )then
          cVar2S18S32N035P017P037nsss(0) <='1';
          else
          cVar2S18S32N035P017P037nsss(0) <='0';
          end if;
        if(cVar1S19S32N036P060P048P063(0)='1' AND  B( 1)='0' AND A( 1)='0' AND E( 0)='1' )then
          cVar2S19S32N035N017P068nsss(0) <='1';
          else
          cVar2S19S32N035N017P068nsss(0) <='0';
          end if;
        if(cVar1S21S32N036P060P048N006(0)='1' AND  A( 5)='1' )then
          cVar2S21S32P009nsss(0) <='1';
          else
          cVar2S21S32P009nsss(0) <='0';
          end if;
        if(cVar1S22S32N036N060P058P054(0)='1' AND  A( 0)='0' AND D( 8)='1' AND E(11)='0' )then
          cVar2S22S32P019P067P057nsss(0) <='1';
          else
          cVar2S22S32P019P067P057nsss(0) <='0';
          end if;
        if(cVar1S23S32N036N060P058P054(0)='1' AND  A( 0)='0' AND D( 8)='0' )then
          cVar2S23S32P019N067psss(0) <='1';
          else
          cVar2S23S32P019N067psss(0) <='0';
          end if;
        if(cVar1S24S32N036N060P058P054(0)='1' AND  A( 0)='1' AND D( 8)='0' AND A(10)='0' )then
          cVar2S24S32P019P067P018nsss(0) <='1';
          else
          cVar2S24S32P019P067P018nsss(0) <='0';
          end if;
        if(cVar1S25S32N036N060P058P054(0)='1' AND  A( 0)='1' AND D( 8)='1' AND D( 0)='1' )then
          cVar2S25S32P019P067P066nsss(0) <='1';
          else
          cVar2S25S32P019P067P066nsss(0) <='0';
          end if;
        if(cVar1S26S32N036N060P058N054(0)='1' AND  E( 3)='0' AND D( 7)='1' AND E( 7)='1' )then
          cVar2S26S32P056P038P040nsss(0) <='1';
          else
          cVar2S26S32P056P038P040nsss(0) <='0';
          end if;
        if(cVar1S27S32N036N060P058N054(0)='1' AND  E( 3)='0' AND D( 7)='0' AND B(10)='1' )then
          cVar2S27S32P056N038P034nsss(0) <='1';
          else
          cVar2S27S32P056N038P034nsss(0) <='0';
          end if;
        if(cVar1S28S32N036N060P058N054(0)='1' AND  E( 3)='1' AND E( 8)='1' AND A( 0)='1' )then
          cVar2S28S32P056P069P019nsss(0) <='1';
          else
          cVar2S28S32P056P069P019nsss(0) <='0';
          end if;
        if(cVar1S29S32N036N060P058P056(0)='1' AND  A(12)='1' AND E(11)='0' )then
          cVar2S29S32P014P057nsss(0) <='1';
          else
          cVar2S29S32P014P057nsss(0) <='0';
          end if;
        if(cVar1S30S32N036N060P058P056(0)='1' AND  A(12)='0' AND A( 2)='1' AND A(13)='1' )then
          cVar2S30S32N014P015P012nsss(0) <='1';
          else
          cVar2S30S32N014P015P012nsss(0) <='0';
          end if;
        if(cVar1S31S32N036N060P058P056(0)='1' AND  A(12)='0' AND A( 2)='0' AND B( 0)='1' )then
          cVar2S31S32N014N015P037nsss(0) <='1';
          else
          cVar2S31S32N014N015P037nsss(0) <='0';
          end if;
        if(cVar1S32S32N036N060P058N056(0)='1' AND  A(10)='0' AND E(10)='1' AND A( 0)='1' )then
          cVar2S32S32P018P061P019nsss(0) <='1';
          else
          cVar2S32S32P018P061P019nsss(0) <='0';
          end if;
        if(cVar1S1S33P034P049P026N018(0)='1' AND  E(12)='0' AND A(15)='0' AND E( 5)='0' )then
          cVar2S1S33P053P008P048nsss(0) <='1';
          else
          cVar2S1S33P053P008P048nsss(0) <='0';
          end if;
        if(cVar1S2S33P034P049P026N018(0)='1' AND  E(12)='0' AND A(15)='1' AND D( 1)='0' )then
          cVar2S2S33P053P008P062nsss(0) <='1';
          else
          cVar2S2S33P053P008P062nsss(0) <='0';
          end if;
        if(cVar1S3S33P034P049N026P024(0)='1' AND  B( 1)='0' AND E(14)='0' AND E( 5)='0' )then
          cVar2S3S33P035P045P048nsss(0) <='1';
          else
          cVar2S3S33P035P045P048nsss(0) <='0';
          end if;
        if(cVar1S4S33P034P049N026P024(0)='1' AND  B( 1)='1' AND E( 1)='0' )then
          cVar2S4S33P035P064nsss(0) <='1';
          else
          cVar2S4S33P035P064nsss(0) <='0';
          end if;
        if(cVar1S5S33P034P049N026N024(0)='1' AND  B( 5)='1' AND E( 5)='0' )then
          cVar2S5S33P027P048nsss(0) <='1';
          else
          cVar2S5S33P027P048nsss(0) <='0';
          end if;
        if(cVar1S6S33P034P049N026N024(0)='1' AND  B( 5)='0' AND B( 6)='1' AND E( 5)='0' )then
          cVar2S6S33N027P025P048nsss(0) <='1';
          else
          cVar2S6S33N027P025P048nsss(0) <='0';
          end if;
        if(cVar1S7S33P034P049N026N024(0)='1' AND  B( 5)='0' AND B( 6)='0' AND E( 2)='1' )then
          cVar2S7S33N027N025P060nsss(0) <='1';
          else
          cVar2S7S33N027N025P060nsss(0) <='0';
          end if;
        if(cVar1S8S33P034N049P028P011(0)='1' AND  D( 0)='0' )then
          cVar2S8S33P066nsss(0) <='1';
          else
          cVar2S8S33P066nsss(0) <='0';
          end if;
        if(cVar1S9S33P034N049P028P011(0)='1' AND  D( 0)='1' AND D( 1)='0' AND A(13)='0' )then
          cVar2S9S33P066P062P012nsss(0) <='1';
          else
          cVar2S9S33P066P062P012nsss(0) <='0';
          end if;
        if(cVar1S10S33P034N049P028N011(0)='1' AND  A(14)='1' AND A( 2)='1' )then
          cVar2S10S33P010P015nsss(0) <='1';
          else
          cVar2S10S33P010P015nsss(0) <='0';
          end if;
        if(cVar1S11S33P034N049P028N011(0)='1' AND  A(14)='1' AND A( 2)='0' AND D( 1)='0' )then
          cVar2S11S33P010N015P062nsss(0) <='1';
          else
          cVar2S11S33P010N015P062nsss(0) <='0';
          end if;
        if(cVar1S12S33P034N049P028N011(0)='1' AND  A(14)='0' AND E(12)='1' AND D( 0)='0' )then
          cVar2S12S33N010P053P066nsss(0) <='1';
          else
          cVar2S12S33N010P053P066nsss(0) <='0';
          end if;
        if(cVar1S13S33P034N049P028N011(0)='1' AND  A(14)='0' AND E(12)='0' AND E( 4)='1' )then
          cVar2S13S33N010N053P052nsss(0) <='1';
          else
          cVar2S13S33N010N053P052nsss(0) <='0';
          end if;
        if(cVar1S14S33P034N049N028P066(0)='1' AND  A(14)='0' AND A(11)='1' AND A( 1)='0' )then
          cVar2S14S33P010P016P017nsss(0) <='1';
          else
          cVar2S14S33P010P016P017nsss(0) <='0';
          end if;
        if(cVar1S15S33P034N049N028P066(0)='1' AND  A(14)='0' AND A(11)='0' AND A( 0)='1' )then
          cVar2S15S33P010N016P019nsss(0) <='1';
          else
          cVar2S15S33P010N016P019nsss(0) <='0';
          end if;
        if(cVar1S16S33P034N049N028P066(0)='1' AND  A(14)='1' AND B( 4)='1' )then
          cVar2S16S33P010P029nsss(0) <='1';
          else
          cVar2S16S33P010P029nsss(0) <='0';
          end if;
        if(cVar1S17S33P034N049N028N066(0)='1' AND  B( 7)='1' AND E( 6)='1' )then
          cVar2S17S33P023P044nsss(0) <='1';
          else
          cVar2S17S33P023P044nsss(0) <='0';
          end if;
        if(cVar1S18S33P034N049N028N066(0)='1' AND  B( 7)='1' AND E( 6)='0' AND D(14)='1' )then
          cVar2S18S33P023N044P043nsss(0) <='1';
          else
          cVar2S18S33P023N044P043nsss(0) <='0';
          end if;
        if(cVar1S19S33P034N049N028N066(0)='1' AND  B( 7)='0' AND D( 4)='1' )then
          cVar2S19S33N023P050nsss(0) <='1';
          else
          cVar2S19S33N023P050nsss(0) <='0';
          end if;
        if(cVar1S20S33P034N049N028N066(0)='1' AND  B( 7)='0' AND D( 4)='0' AND D( 7)='1' )then
          cVar2S20S33N023N050P038nsss(0) <='1';
          else
          cVar2S20S33N023N050P038nsss(0) <='0';
          end if;
        if(cVar1S21S33P034P014P044P069(0)='1' AND  A( 0)='1' AND A( 3)='0' )then
          cVar2S21S33P019P013nsss(0) <='1';
          else
          cVar2S21S33P019P013nsss(0) <='0';
          end if;
        if(cVar1S22S33P034P014P044P069(0)='1' AND  A( 0)='1' AND A( 3)='1' AND A( 1)='0' )then
          cVar2S22S33P019P013P017nsss(0) <='1';
          else
          cVar2S22S33P019P013P017nsss(0) <='0';
          end if;
        if(cVar1S23S33P034P014P044P069(0)='1' AND  A( 0)='0' AND A( 6)='0' AND D(10)='0' )then
          cVar2S23S33N019P007P059nsss(0) <='1';
          else
          cVar2S23S33N019P007P059nsss(0) <='0';
          end if;
        if(cVar1S24S33P034P014P044N069(0)='1' AND  B( 1)='0' AND D( 1)='1' AND A(14)='0' )then
          cVar2S24S33P035P062P010nsss(0) <='1';
          else
          cVar2S24S33P035P062P010nsss(0) <='0';
          end if;
        if(cVar1S25S33P034P014P044N069(0)='1' AND  B( 1)='0' AND D( 1)='0' AND E(10)='1' )then
          cVar2S25S33P035N062P061nsss(0) <='1';
          else
          cVar2S25S33P035N062P061nsss(0) <='0';
          end if;
        if(cVar1S26S33P034P014P044N069(0)='1' AND  B( 1)='1' AND A(11)='0' AND D(10)='1' )then
          cVar2S26S33P035P016P059nsss(0) <='1';
          else
          cVar2S26S33P035P016P059nsss(0) <='0';
          end if;
        if(cVar1S28S33P034N014P045N062(0)='1' AND  A(10)='0' AND D( 9)='1' )then
          cVar2S28S33P018P063nsss(0) <='1';
          else
          cVar2S28S33P018P063nsss(0) <='0';
          end if;
        if(cVar1S29S33P034N014N045P046(0)='1' AND  A( 2)='1' AND A( 8)='0' AND D( 1)='0' )then
          cVar2S29S33P015P003P062nsss(0) <='1';
          else
          cVar2S29S33P015P003P062nsss(0) <='0';
          end if;
        if(cVar1S30S33P034N014N045P046(0)='1' AND  A( 2)='0' AND A( 0)='1' AND B( 4)='1' )then
          cVar2S30S33N015P019P029nsss(0) <='1';
          else
          cVar2S30S33N015P019P029nsss(0) <='0';
          end if;
        if(cVar1S31S33P034N014N045P046(0)='1' AND  A(11)='1' AND E( 5)='1' )then
          cVar2S31S33P016P048nsss(0) <='1';
          else
          cVar2S31S33P016P048nsss(0) <='0';
          end if;
        if(cVar1S0S34P034P068P032P054(0)='1' AND  E(15)='1' AND A(12)='1' )then
          cVar2S0S34P041P014nsss(0) <='1';
          else
          cVar2S0S34P041P014nsss(0) <='0';
          end if;
        if(cVar1S1S34P034P068P032P054(0)='1' AND  E(15)='0' AND D( 9)='1' AND D( 8)='0' )then
          cVar2S1S34N041P063P067nsss(0) <='1';
          else
          cVar2S1S34N041P063P067nsss(0) <='0';
          end if;
        if(cVar1S2S34P034P068P032P054(0)='1' AND  E(15)='0' AND D( 9)='0' )then
          cVar2S2S34N041N063psss(0) <='1';
          else
          cVar2S2S34N041N063psss(0) <='0';
          end if;
        if(cVar1S3S34P034P068P032P054(0)='1' AND  A(14)='1' )then
          cVar2S3S34P010nsss(0) <='1';
          else
          cVar2S3S34P010nsss(0) <='0';
          end if;
        if(cVar1S4S34P034P068P032P054(0)='1' AND  A(14)='0' AND D( 2)='1' )then
          cVar2S4S34N010P058nsss(0) <='1';
          else
          cVar2S4S34N010P058nsss(0) <='0';
          end if;
        if(cVar1S5S34P034P068N032P059(0)='1' AND  E(10)='0' )then
          cVar2S5S34P061nsss(0) <='1';
          else
          cVar2S5S34P061nsss(0) <='0';
          end if;
        if(cVar1S6S34P034P068N032P059(0)='1' AND  E(10)='1' AND A( 3)='1' AND E( 9)='0' )then
          cVar2S6S34P061P013P065nsss(0) <='1';
          else
          cVar2S6S34P061P013P065nsss(0) <='0';
          end if;
        if(cVar1S7S34P034P068N032P059(0)='1' AND  A( 3)='1' AND B( 1)='0' AND A( 4)='0' )then
          cVar2S7S34P013P035P011nsss(0) <='1';
          else
          cVar2S7S34P013P035P011nsss(0) <='0';
          end if;
        if(cVar1S8S34P034P068N032P059(0)='1' AND  A( 3)='1' AND B( 1)='1' AND B( 2)='1' )then
          cVar2S8S34P013P035P033nsss(0) <='1';
          else
          cVar2S8S34P013P035P033nsss(0) <='0';
          end if;
        if(cVar1S9S34P034P068N032P059(0)='1' AND  A( 3)='0' AND A( 2)='1' AND E( 4)='1' )then
          cVar2S9S34N013P015P052nsss(0) <='1';
          else
          cVar2S9S34N013P015P052nsss(0) <='0';
          end if;
        if(cVar1S10S34P034P068N032P059(0)='1' AND  A( 3)='0' AND A( 2)='0' AND B(12)='1' )then
          cVar2S10S34N013N015P030nsss(0) <='1';
          else
          cVar2S10S34N013N015P030nsss(0) <='0';
          end if;
        if(cVar1S11S34P034P068P019P064(0)='1' AND  D( 0)='1' )then
          cVar2S11S34P066nsss(0) <='1';
          else
          cVar2S11S34P066nsss(0) <='0';
          end if;
        if(cVar1S12S34P034P068P019P064(0)='1' AND  D( 0)='0' AND A( 2)='0' AND A(16)='0' )then
          cVar2S12S34N066P015P006nsss(0) <='1';
          else
          cVar2S12S34N066P015P006nsss(0) <='0';
          end if;
        if(cVar1S13S34P034P068P019P064(0)='1' AND  D( 0)='0' AND A( 2)='1' AND A( 6)='1' )then
          cVar2S13S34N066P015P007nsss(0) <='1';
          else
          cVar2S13S34N066P015P007nsss(0) <='0';
          end if;
        if(cVar1S14S34P034P068P019P064(0)='1' AND  A( 1)='1' AND D( 2)='0' AND B( 1)='1' )then
          cVar2S14S34P017P058P035nsss(0) <='1';
          else
          cVar2S14S34P017P058P035nsss(0) <='0';
          end if;
        if(cVar1S15S34P034P068P019P064(0)='1' AND  A( 1)='1' AND D( 2)='1' AND E( 2)='1' )then
          cVar2S15S34P017P058P060nsss(0) <='1';
          else
          cVar2S15S34P017P058P060nsss(0) <='0';
          end if;
        if(cVar1S16S34P034P068P019P064(0)='1' AND  A( 1)='0' AND A( 2)='1' AND A(12)='0' )then
          cVar2S16S34N017P015P014nsss(0) <='1';
          else
          cVar2S16S34N017P015P014nsss(0) <='0';
          end if;
        if(cVar1S17S34P034P068P019P036(0)='1' AND  A(11)='1' AND E( 2)='0' AND A( 4)='0' )then
          cVar2S17S34P016P060P011nsss(0) <='1';
          else
          cVar2S17S34P016P060P011nsss(0) <='0';
          end if;
        if(cVar1S18S34P034P068P019P036(0)='1' AND  A(11)='0' AND A(13)='0' AND D( 9)='0' )then
          cVar2S18S34N016P012P063nsss(0) <='1';
          else
          cVar2S18S34N016P012P063nsss(0) <='0';
          end if;
        if(cVar1S19S34P034P068P019P036(0)='1' AND  A(11)='0' AND A(13)='1' AND A(14)='1' )then
          cVar2S19S34N016P012P010nsss(0) <='1';
          else
          cVar2S19S34N016P012P010nsss(0) <='0';
          end if;
        if(cVar1S20S34P034P068P019P036(0)='1' AND  D( 0)='0' AND E( 8)='1' )then
          cVar2S20S34P066P069nsss(0) <='1';
          else
          cVar2S20S34P066P069nsss(0) <='0';
          end if;
        if(cVar1S21S34P034P068P019P036(0)='1' AND  D( 0)='0' AND E( 8)='0' AND A(11)='1' )then
          cVar2S21S34P066N069P016nsss(0) <='1';
          else
          cVar2S21S34P066N069P016nsss(0) <='0';
          end if;
        if(cVar1S22S34P034P068P019P036(0)='1' AND  D( 0)='1' AND A( 4)='1' AND A( 3)='0' )then
          cVar2S22S34P066P011P013nsss(0) <='1';
          else
          cVar2S22S34P066P011P013nsss(0) <='0';
          end if;
        if(cVar1S23S34P034P068P019P036(0)='1' AND  D( 0)='1' AND A( 4)='0' AND D(11)='1' )then
          cVar2S23S34P066N011P055nsss(0) <='1';
          else
          cVar2S23S34P066N011P055nsss(0) <='0';
          end if;
        if(cVar1S24S34P034P062P065P018(0)='1' AND  B( 1)='0' AND A(13)='0' )then
          cVar2S24S34P035P012nsss(0) <='1';
          else
          cVar2S24S34P035P012nsss(0) <='0';
          end if;
        if(cVar1S25S34P034P062P065P018(0)='1' AND  B( 1)='0' AND A(13)='1' AND A( 0)='1' )then
          cVar2S25S34P035P012P019nsss(0) <='1';
          else
          cVar2S25S34P035P012P019nsss(0) <='0';
          end if;
        if(cVar1S26S34P034P062P065P018(0)='1' AND  B( 1)='1' AND A( 0)='0' AND A(11)='0' )then
          cVar2S26S34P035P019P016nsss(0) <='1';
          else
          cVar2S26S34P035P019P016nsss(0) <='0';
          end if;
        if(cVar1S27S34P034P062P065P018(0)='1' AND  A(12)='1' AND B( 0)='0' )then
          cVar2S27S34P014P037nsss(0) <='1';
          else
          cVar2S27S34P014P037nsss(0) <='0';
          end if;
        if(cVar1S28S34P034P062P065P018(0)='1' AND  A(12)='0' AND E( 8)='0' AND E(10)='0' )then
          cVar2S28S34N014P069P061nsss(0) <='1';
          else
          cVar2S28S34N014P069P061nsss(0) <='0';
          end if;
        if(cVar1S29S34P034P062P065P017(0)='1' AND  D(10)='1' )then
          cVar2S29S34P059nsss(0) <='1';
          else
          cVar2S29S34P059nsss(0) <='0';
          end if;
        if(cVar1S30S34P034P062P065P017(0)='1' AND  D(10)='0' AND B( 0)='1' )then
          cVar2S30S34N059P037nsss(0) <='1';
          else
          cVar2S30S34N059P037nsss(0) <='0';
          end if;
        if(cVar1S31S34P034P062P065P017(0)='1' AND  D(10)='0' AND B( 0)='0' AND D( 2)='0' )then
          cVar2S31S34N059N037P058nsss(0) <='1';
          else
          cVar2S31S34N059N037P058nsss(0) <='0';
          end if;
        if(cVar1S32S34P034P062P065N017(0)='1' AND  B( 9)='1' AND A( 2)='1' )then
          cVar2S32S34P036P015nsss(0) <='1';
          else
          cVar2S32S34P036P015nsss(0) <='0';
          end if;
        if(cVar1S33S34P034P062P065N017(0)='1' AND  B( 9)='1' AND A( 2)='0' AND A( 0)='0' )then
          cVar2S33S34P036N015P019nsss(0) <='1';
          else
          cVar2S33S34P036N015P019nsss(0) <='0';
          end if;
        if(cVar1S34S34P034P062P065N017(0)='1' AND  B( 9)='0' AND A( 0)='1' AND B( 1)='1' )then
          cVar2S34S34N036P019P035nsss(0) <='1';
          else
          cVar2S34S34N036P019P035nsss(0) <='0';
          end if;
        if(cVar1S35S34P034P062P065N017(0)='1' AND  B( 9)='0' AND A( 0)='0' AND A(11)='0' )then
          cVar2S35S34N036N019P016nsss(0) <='1';
          else
          cVar2S35S34N036N019P016nsss(0) <='0';
          end if;
        if(cVar1S36S34P034N062P008P063(0)='1' AND  D( 0)='0' AND E( 2)='0' AND A( 1)='1' )then
          cVar2S36S34P066P060P017nsss(0) <='1';
          else
          cVar2S36S34P066P060P017nsss(0) <='0';
          end if;
        if(cVar1S37S34P034N062P008P063(0)='1' AND  D( 0)='0' AND E( 2)='1' AND A( 4)='1' )then
          cVar2S37S34P066P060P011nsss(0) <='1';
          else
          cVar2S37S34P066P060P011nsss(0) <='0';
          end if;
        if(cVar1S38S34P034N062P008P063(0)='1' AND  D( 0)='1' AND A( 1)='0' AND A(10)='0' )then
          cVar2S38S34P066P017P018nsss(0) <='1';
          else
          cVar2S38S34P066P017P018nsss(0) <='0';
          end if;
        if(cVar1S39S34P034N062P008N063(0)='1' AND  E(10)='1' AND E( 0)='1' AND A( 2)='1' )then
          cVar2S39S34P061P068P015nsss(0) <='1';
          else
          cVar2S39S34P061P068P015nsss(0) <='0';
          end if;
        if(cVar1S40S34P034N062P008N063(0)='1' AND  E(10)='1' AND E( 0)='0' AND A(11)='1' )then
          cVar2S40S34P061N068P016nsss(0) <='1';
          else
          cVar2S40S34P061N068P016nsss(0) <='0';
          end if;
        if(cVar1S41S34P034N062P008N063(0)='1' AND  E(10)='0' AND E( 2)='1' AND D( 2)='1' )then
          cVar2S41S34N061P060P058nsss(0) <='1';
          else
          cVar2S41S34N061P060P058nsss(0) <='0';
          end if;
        if(cVar1S42S34P034N062P008P026(0)='1' AND  A(11)='0' )then
          cVar2S42S34P016nsss(0) <='1';
          else
          cVar2S42S34P016nsss(0) <='0';
          end if;
        if(cVar1S43S34P034N062P008N026(0)='1' AND  D( 4)='1' AND E( 9)='1' )then
          cVar2S43S34P050P065nsss(0) <='1';
          else
          cVar2S43S34P050P065nsss(0) <='0';
          end if;
        if(cVar1S44S34P034N062P008N026(0)='1' AND  D( 4)='0' AND E( 3)='1' )then
          cVar2S44S34N050P056nsss(0) <='1';
          else
          cVar2S44S34N050P056nsss(0) <='0';
          end if;
        if(cVar1S1S35P061P064P030N013(0)='1' AND  A(11)='0' AND E(11)='1' )then
          cVar2S1S35P016P057nsss(0) <='1';
          else
          cVar2S1S35P016P057nsss(0) <='0';
          end if;
        if(cVar1S2S35P061P064P030N013(0)='1' AND  A(11)='0' AND E(11)='0' AND A( 2)='1' )then
          cVar2S2S35P016N057P015nsss(0) <='1';
          else
          cVar2S2S35P016N057P015nsss(0) <='0';
          end if;
        if(cVar1S3S35P061P064N030P057(0)='1' AND  B( 2)='1' AND D( 2)='0' AND B(11)='0' )then
          cVar2S3S35P033P058P032nsss(0) <='1';
          else
          cVar2S3S35P033P058P032nsss(0) <='0';
          end if;
        if(cVar1S4S35P061P064N030P057(0)='1' AND  B( 2)='1' AND D( 2)='1' AND D( 9)='0' )then
          cVar2S4S35P033P058P063nsss(0) <='1';
          else
          cVar2S4S35P033P058P063nsss(0) <='0';
          end if;
        if(cVar1S5S35P061P064N030P057(0)='1' AND  B( 2)='0' AND E( 3)='0' )then
          cVar2S5S35N033P056nsss(0) <='1';
          else
          cVar2S5S35N033P056nsss(0) <='0';
          end if;
        if(cVar1S6S35P061P064N030P057(0)='1' AND  B( 2)='0' AND E( 3)='1' AND A(13)='1' )then
          cVar2S6S35N033P056P012nsss(0) <='1';
          else
          cVar2S6S35N033P056P012nsss(0) <='0';
          end if;
        if(cVar1S7S35P061P064N030P057(0)='1' AND  B( 0)='1' )then
          cVar2S7S35P037nsss(0) <='1';
          else
          cVar2S7S35P037nsss(0) <='0';
          end if;
        if(cVar1S9S35P061P064P058N008(0)='1' AND  A(10)='1' AND B(10)='0' )then
          cVar2S9S35P018P034nsss(0) <='1';
          else
          cVar2S9S35P018P034nsss(0) <='0';
          end if;
        if(cVar1S10S35P061P064P058N008(0)='1' AND  A(10)='1' AND B(10)='1' AND A(12)='1' )then
          cVar2S10S35P018P034P014nsss(0) <='1';
          else
          cVar2S10S35P018P034P014nsss(0) <='0';
          end if;
        if(cVar1S11S35P061P064P058N008(0)='1' AND  A(10)='0' AND E( 0)='0' AND B( 2)='1' )then
          cVar2S11S35N018P068P033nsss(0) <='1';
          else
          cVar2S11S35N018P068P033nsss(0) <='0';
          end if;
        if(cVar1S12S35P061P064P058P063(0)='1' AND  B( 1)='1' )then
          cVar2S12S35P035nsss(0) <='1';
          else
          cVar2S12S35P035nsss(0) <='0';
          end if;
        if(cVar1S13S35N061P057P026P007(0)='1' AND  E( 3)='0' AND E( 4)='0' )then
          cVar2S13S35P056P052nsss(0) <='1';
          else
          cVar2S13S35P056P052nsss(0) <='0';
          end if;
        if(cVar1S14S35N061P057P026P007(0)='1' AND  E( 3)='0' AND E( 4)='1' AND A(13)='1' )then
          cVar2S14S35P056P052P012nsss(0) <='1';
          else
          cVar2S14S35P056P052P012nsss(0) <='0';
          end if;
        if(cVar1S15S35N061P057P026P007(0)='1' AND  E( 3)='1' AND D( 3)='1' AND E( 8)='0' )then
          cVar2S15S35P056P054P069nsss(0) <='1';
          else
          cVar2S15S35P056P054P069nsss(0) <='0';
          end if;
        if(cVar1S16S35N061P057P026P007(0)='1' AND  E( 1)='0' AND A(11)='0' AND A(10)='1' )then
          cVar2S16S35P064P016P018nsss(0) <='1';
          else
          cVar2S16S35P064P016P018nsss(0) <='0';
          end if;
        if(cVar1S17S35N061P057P026N030(0)='1' AND  A( 1)='1' AND A( 0)='0' )then
          cVar2S17S35P017P019nsss(0) <='1';
          else
          cVar2S17S35P017P019nsss(0) <='0';
          end if;
        if(cVar1S18S35N061N057P064P065(0)='1' AND  B( 2)='0' AND D(11)='0' AND B( 4)='0' )then
          cVar2S18S35P033P055P029nsss(0) <='1';
          else
          cVar2S18S35P033P055P029nsss(0) <='0';
          end if;
        if(cVar1S19S35N061N057P064P065(0)='1' AND  B( 2)='0' AND D(11)='1' AND A( 4)='1' )then
          cVar2S19S35P033P055P011nsss(0) <='1';
          else
          cVar2S19S35P033P055P011nsss(0) <='0';
          end if;
        if(cVar1S20S35N061N057P064P065(0)='1' AND  B( 2)='1' AND A( 1)='1' AND A( 0)='0' )then
          cVar2S20S35P033P017P019nsss(0) <='1';
          else
          cVar2S20S35P033P017P019nsss(0) <='0';
          end if;
        if(cVar1S21S35N061N057P064P065(0)='1' AND  B( 2)='1' AND A( 1)='0' AND A(11)='1' )then
          cVar2S21S35P033N017P016nsss(0) <='1';
          else
          cVar2S21S35P033N017P016nsss(0) <='0';
          end if;
        if(cVar1S22S35N061N057P064P065(0)='1' AND  A(10)='1' AND A( 2)='1' AND A( 4)='0' )then
          cVar2S22S35P018P015P011nsss(0) <='1';
          else
          cVar2S22S35P018P015P011nsss(0) <='0';
          end if;
        if(cVar1S23S35N061N057P064P065(0)='1' AND  A(10)='1' AND A( 2)='0' AND D( 9)='0' )then
          cVar2S23S35P018N015P063nsss(0) <='1';
          else
          cVar2S23S35P018N015P063nsss(0) <='0';
          end if;
        if(cVar1S24S35N061N057N064P063(0)='1' AND  B( 1)='1' AND B( 9)='0' AND E( 9)='1' )then
          cVar2S24S35P035P036P065nsss(0) <='1';
          else
          cVar2S24S35P035P036P065nsss(0) <='0';
          end if;
        if(cVar1S25S35N061N057N064P063(0)='1' AND  B( 1)='1' AND B( 9)='1' AND A( 0)='0' )then
          cVar2S25S35P035P036P019nsss(0) <='1';
          else
          cVar2S25S35P035P036P019nsss(0) <='0';
          end if;
        if(cVar1S26S35N061N057N064N063(0)='1' AND  E(13)='1' AND A( 5)='1' AND E( 5)='0' )then
          cVar2S26S35P049P009P048nsss(0) <='1';
          else
          cVar2S26S35P049P009P048nsss(0) <='0';
          end if;
        if(cVar1S27S35N061N057N064N063(0)='1' AND  E(13)='0' AND D( 8)='0' AND E( 2)='1' )then
          cVar2S27S35N049N067P060nsss(0) <='1';
          else
          cVar2S27S35N049N067P060nsss(0) <='0';
          end if;
        if(cVar1S0S36P063P062P065P066(0)='1' AND  B( 1)='1' AND A( 0)='0' )then
          cVar2S0S36P035P019nsss(0) <='1';
          else
          cVar2S0S36P035P019nsss(0) <='0';
          end if;
        if(cVar1S1S36P063P062P065P066(0)='1' AND  B( 1)='1' AND A( 0)='1' AND B( 9)='0' )then
          cVar2S1S36P035P019P036nsss(0) <='1';
          else
          cVar2S1S36P035P019P036nsss(0) <='0';
          end if;
        if(cVar1S2S36P063P062P065P066(0)='1' AND  B( 1)='0' AND B( 6)='0' AND D( 2)='0' )then
          cVar2S2S36N035P025P058nsss(0) <='1';
          else
          cVar2S2S36N035P025P058nsss(0) <='0';
          end if;
        if(cVar1S3S36P063P062P065P066(0)='1' AND  B( 1)='0' AND B( 6)='1' AND B(10)='0' )then
          cVar2S3S36N035P025P034nsss(0) <='1';
          else
          cVar2S3S36N035P025P034nsss(0) <='0';
          end if;
        if(cVar1S4S36P063P062P065P066(0)='1' AND  E( 4)='0' AND D(10)='0' )then
          cVar2S4S36P052P059nsss(0) <='1';
          else
          cVar2S4S36P052P059nsss(0) <='0';
          end if;
        if(cVar1S5S36P063P062N065P007(0)='1' AND  A( 1)='1' AND E(10)='1' )then
          cVar2S5S36P017P061nsss(0) <='1';
          else
          cVar2S5S36P017P061nsss(0) <='0';
          end if;
        if(cVar1S6S36P063P062N065P007(0)='1' AND  A( 1)='1' AND E(10)='0' AND E( 2)='1' )then
          cVar2S6S36P017N061P060nsss(0) <='1';
          else
          cVar2S6S36P017N061P060nsss(0) <='0';
          end if;
        if(cVar1S7S36P063P062N065P007(0)='1' AND  A( 1)='0' AND A( 0)='1' AND A( 2)='1' )then
          cVar2S7S36N017P019P015nsss(0) <='1';
          else
          cVar2S7S36N017P019P015nsss(0) <='0';
          end if;
        if(cVar1S8S36P063P062N065P007(0)='1' AND  B(10)='0' AND A( 5)='1' )then
          cVar2S8S36P034P009nsss(0) <='1';
          else
          cVar2S8S36P034P009nsss(0) <='0';
          end if;
        if(cVar1S9S36P063P062P048P054(0)='1' AND  A(13)='1' AND E( 2)='1' )then
          cVar2S9S36P012P060nsss(0) <='1';
          else
          cVar2S9S36P012P060nsss(0) <='0';
          end if;
        if(cVar1S10S36P063P062P048P054(0)='1' AND  A(13)='1' AND E( 2)='0' AND D(11)='0' )then
          cVar2S10S36P012N060P055nsss(0) <='1';
          else
          cVar2S10S36P012N060P055nsss(0) <='0';
          end if;
        if(cVar1S11S36P063P062P048P054(0)='1' AND  A(13)='0' AND E( 7)='1' )then
          cVar2S11S36N012P040nsss(0) <='1';
          else
          cVar2S11S36N012P040nsss(0) <='0';
          end if;
        if(cVar1S12S36P063P062P048P054(0)='1' AND  A(13)='0' AND E( 7)='0' AND D(13)='0' )then
          cVar2S12S36N012N040P047nsss(0) <='1';
          else
          cVar2S12S36N012N040P047nsss(0) <='0';
          end if;
        if(cVar1S13S36P063P062P048P054(0)='1' AND  D( 0)='1' )then
          cVar2S13S36P066nsss(0) <='1';
          else
          cVar2S13S36P066nsss(0) <='0';
          end if;
        if(cVar1S14S36P063P062P048P046(0)='1' AND  B( 1)='1' )then
          cVar2S14S36P035nsss(0) <='1';
          else
          cVar2S14S36P035nsss(0) <='0';
          end if;
        if(cVar1S15S36N063P067P064P019(0)='1' AND  D( 2)='0' AND D( 0)='0' AND D( 3)='0' )then
          cVar2S15S36P058P066P054nsss(0) <='1';
          else
          cVar2S15S36P058P066P054nsss(0) <='0';
          end if;
        if(cVar1S16S36N063P067P064P019(0)='1' AND  D( 2)='0' AND D( 0)='1' AND E(12)='0' )then
          cVar2S16S36P058P066P053nsss(0) <='1';
          else
          cVar2S16S36P058P066P053nsss(0) <='0';
          end if;
        if(cVar1S17S36N063P067P064P019(0)='1' AND  D( 2)='1' AND A(10)='0' )then
          cVar2S17S36P058P018nsss(0) <='1';
          else
          cVar2S17S36P058P018nsss(0) <='0';
          end if;
        if(cVar1S18S36N063P067P064P019(0)='1' AND  D( 2)='1' AND A(10)='1' AND A( 3)='1' )then
          cVar2S18S36P058P018P013nsss(0) <='1';
          else
          cVar2S18S36P058P018P013nsss(0) <='0';
          end if;
        if(cVar1S19S36N063P067P064N019(0)='1' AND  D( 1)='0' AND A(10)='1' AND E( 0)='0' )then
          cVar2S19S36P062P018P068nsss(0) <='1';
          else
          cVar2S19S36P062P018P068nsss(0) <='0';
          end if;
        if(cVar1S20S36N063P067P064N019(0)='1' AND  D( 1)='0' AND A(10)='0' AND E( 0)='1' )then
          cVar2S20S36P062N018P068nsss(0) <='1';
          else
          cVar2S20S36P062N018P068nsss(0) <='0';
          end if;
        if(cVar1S21S36N063P067P064N019(0)='1' AND  D( 1)='1' AND E( 2)='1' AND D( 0)='1' )then
          cVar2S21S36P062P060P066nsss(0) <='1';
          else
          cVar2S21S36P062P060P066nsss(0) <='0';
          end if;
        if(cVar1S22S36N063P067P064P037(0)='1' AND  B( 1)='0' AND B(10)='0' AND E( 0)='0' )then
          cVar2S22S36P035P034P068nsss(0) <='1';
          else
          cVar2S22S36P035P034P068nsss(0) <='0';
          end if;
        if(cVar1S23S36N063P067P064P037(0)='1' AND  B( 1)='1' AND A( 0)='0' AND A( 1)='1' )then
          cVar2S23S36P035P019P017nsss(0) <='1';
          else
          cVar2S23S36P035P019P017nsss(0) <='0';
          end if;
        if(cVar1S24S36N063P067P064N037(0)='1' AND  A(12)='1' AND A(14)='0' AND A(10)='1' )then
          cVar2S24S36P014P010P018nsss(0) <='1';
          else
          cVar2S24S36P014P010P018nsss(0) <='0';
          end if;
        if(cVar1S25S36N063P067P064N037(0)='1' AND  A(12)='0' AND A(11)='1' AND A( 0)='0' )then
          cVar2S25S36N014P016P019nsss(0) <='1';
          else
          cVar2S25S36N014P016P019nsss(0) <='0';
          end if;
        if(cVar1S26S36N063N067P053P051(0)='1' AND  E( 4)='0' AND B(14)='1' )then
          cVar2S26S36P052P026nsss(0) <='1';
          else
          cVar2S26S36P052P026nsss(0) <='0';
          end if;
        if(cVar1S27S36N063N067P053P051(0)='1' AND  E( 4)='0' AND B(14)='0' AND E( 2)='0' )then
          cVar2S27S36P052N026P060nsss(0) <='1';
          else
          cVar2S27S36P052N026P060nsss(0) <='0';
          end if;
        if(cVar1S28S36N063N067P053P051(0)='1' AND  E( 4)='1' AND A(10)='1' )then
          cVar2S28S36P052P018nsss(0) <='1';
          else
          cVar2S28S36P052P018nsss(0) <='0';
          end if;
        if(cVar1S29S36N063N067P053N051(0)='1' AND  B(14)='0' AND A( 0)='0' AND A(10)='0' )then
          cVar2S29S36P026P019P018nsss(0) <='1';
          else
          cVar2S29S36P026P019P018nsss(0) <='0';
          end if;
        if(cVar1S30S36N063N067N053P022(0)='1' AND  D(14)='1' )then
          cVar2S30S36P043nsss(0) <='1';
          else
          cVar2S30S36P043nsss(0) <='0';
          end if;
        if(cVar1S31S36N063N067N053P022(0)='1' AND  D(14)='0' AND B( 1)='0' AND B(14)='0' )then
          cVar2S31S36N043P035P026nsss(0) <='1';
          else
          cVar2S31S36N043P035P026nsss(0) <='0';
          end if;
        if(cVar1S32S36N063N067N053N022(0)='1' AND  E( 0)='1' AND D( 0)='1' AND D(15)='1' )then
          cVar2S32S36P068P066P039nsss(0) <='1';
          else
          cVar2S32S36P068P066P039nsss(0) <='0';
          end if;
        if(cVar1S33S36N063N067N053N022(0)='1' AND  E( 0)='0' AND E( 8)='0' AND D(13)='1' )then
          cVar2S33S36N068P069P047nsss(0) <='1';
          else
          cVar2S33S36N068P069P047nsss(0) <='0';
          end if;
        if(cVar1S0S37P065P067P000P068(0)='1' AND  D( 0)='1' AND B( 9)='1' AND A(10)='1' )then
          cVar2S0S37P066P036P018nsss(0) <='1';
          else
          cVar2S0S37P066P036P018nsss(0) <='0';
          end if;
        if(cVar1S1S37P065P067P000P068(0)='1' AND  D( 0)='1' AND B( 9)='0' AND A( 2)='0' )then
          cVar2S1S37P066N036P015nsss(0) <='1';
          else
          cVar2S1S37P066N036P015nsss(0) <='0';
          end if;
        if(cVar1S2S37P065P067P000P068(0)='1' AND  D( 0)='0' AND E( 1)='1' )then
          cVar2S2S37N066P064nsss(0) <='1';
          else
          cVar2S2S37N066P064nsss(0) <='0';
          end if;
        if(cVar1S3S37P065P067P000N068(0)='1' AND  A( 4)='1' AND A(11)='0' AND B( 9)='0' )then
          cVar2S3S37P011P016P036nsss(0) <='1';
          else
          cVar2S3S37P011P016P036nsss(0) <='0';
          end if;
        if(cVar1S4S37P065P067P000N068(0)='1' AND  A( 4)='0' AND D( 1)='1' AND E(13)='0' )then
          cVar2S4S37N011P062P049nsss(0) <='1';
          else
          cVar2S4S37N011P062P049nsss(0) <='0';
          end if;
        if(cVar1S5S37P065P067P000N068(0)='1' AND  A( 4)='0' AND D( 1)='0' AND D(10)='1' )then
          cVar2S5S37N011N062P059nsss(0) <='1';
          else
          cVar2S5S37N011N062P059nsss(0) <='0';
          end if;
        if(cVar1S6S37P065P067P000P053(0)='1' AND  E( 6)='0' AND E(15)='1' )then
          cVar2S6S37P044P041nsss(0) <='1';
          else
          cVar2S6S37P044P041nsss(0) <='0';
          end if;
        if(cVar1S7S37P065P067P062P056(0)='1' AND  E( 4)='0' AND E( 2)='0' AND E( 0)='0' )then
          cVar2S7S37P052P060P068nsss(0) <='1';
          else
          cVar2S7S37P052P060P068nsss(0) <='0';
          end if;
        if(cVar1S8S37P065P067P062N056(0)='1' AND  A(12)='0' AND B(10)='0' AND A( 0)='0' )then
          cVar2S8S37P014P034P019nsss(0) <='1';
          else
          cVar2S8S37P014P034P019nsss(0) <='0';
          end if;
        if(cVar1S9S37P065P067P062N056(0)='1' AND  A(12)='0' AND B(10)='1' AND A( 4)='1' )then
          cVar2S9S37P014P034P011nsss(0) <='1';
          else
          cVar2S9S37P014P034P011nsss(0) <='0';
          end if;
        if(cVar1S10S37P065P067P062N056(0)='1' AND  A(12)='1' AND D(13)='1' )then
          cVar2S10S37P014P047nsss(0) <='1';
          else
          cVar2S10S37P014P047nsss(0) <='0';
          end if;
        if(cVar1S11S37P065P067P062N056(0)='1' AND  A(12)='1' AND D(13)='0' AND D(11)='1' )then
          cVar2S11S37P014N047P055nsss(0) <='1';
          else
          cVar2S11S37P014N047P055nsss(0) <='0';
          end if;
        if(cVar1S12S37P065P067P062P018(0)='1' AND  D( 2)='0' AND A(12)='1' )then
          cVar2S12S37P058P014nsss(0) <='1';
          else
          cVar2S12S37P058P014nsss(0) <='0';
          end if;
        if(cVar1S13S37P065P067P062P018(0)='1' AND  D( 2)='0' AND A(12)='0' AND A( 0)='0' )then
          cVar2S13S37P058N014P019nsss(0) <='1';
          else
          cVar2S13S37P058N014P019nsss(0) <='0';
          end if;
        if(cVar1S14S37P065P067P062P018(0)='1' AND  D( 2)='1' AND A( 2)='1' )then
          cVar2S14S37P058P015nsss(0) <='1';
          else
          cVar2S14S37P058P015nsss(0) <='0';
          end if;
        if(cVar1S15S37P065P067P062P018(0)='1' AND  A( 0)='1' AND A(14)='0' AND E( 1)='1' )then
          cVar2S15S37P019P010P064nsss(0) <='1';
          else
          cVar2S15S37P019P010P064nsss(0) <='0';
          end if;
        if(cVar1S16S37P065P067P062P018(0)='1' AND  A( 0)='1' AND A(14)='1' AND D( 0)='1' )then
          cVar2S16S37P019P010P066nsss(0) <='1';
          else
          cVar2S16S37P019P010P066nsss(0) <='0';
          end if;
        if(cVar1S17S37P065P060P058P069(0)='1' AND  D( 9)='1' )then
          cVar2S17S37P063nsss(0) <='1';
          else
          cVar2S17S37P063nsss(0) <='0';
          end if;
        if(cVar1S18S37P065P060P058N069(0)='1' AND  A(13)='1' AND B( 2)='0' )then
          cVar2S18S37P012P033nsss(0) <='1';
          else
          cVar2S18S37P012P033nsss(0) <='0';
          end if;
        if(cVar1S19S37P065P060P058N069(0)='1' AND  A(13)='1' AND B( 2)='1' AND A(11)='0' )then
          cVar2S19S37P012P033P016nsss(0) <='1';
          else
          cVar2S19S37P012P033P016nsss(0) <='0';
          end if;
        if(cVar1S20S37P065P060P058N069(0)='1' AND  A(13)='0' AND A(12)='1' AND B( 9)='0' )then
          cVar2S20S37N012P014P036nsss(0) <='1';
          else
          cVar2S20S37N012P014P036nsss(0) <='0';
          end if;
        if(cVar1S21S37P065P060P058N069(0)='1' AND  A(13)='0' AND A(12)='0' AND A( 0)='1' )then
          cVar2S21S37N012N014P019nsss(0) <='1';
          else
          cVar2S21S37N012N014P019nsss(0) <='0';
          end if;
        if(cVar1S22S37P065P060N058P018(0)='1' AND  A( 2)='0' )then
          cVar2S22S37P015nsss(0) <='1';
          else
          cVar2S22S37P015nsss(0) <='0';
          end if;
        if(cVar1S23S37P065N060P062P063(0)='1' AND  D( 0)='0' AND E( 8)='0' AND E( 0)='0' )then
          cVar2S23S37P066P069P068nsss(0) <='1';
          else
          cVar2S23S37P066P069P068nsss(0) <='0';
          end if;
        if(cVar1S24S37P065N060P062P063(0)='1' AND  D( 0)='1' AND B( 9)='1' AND E( 4)='0' )then
          cVar2S24S37P066P036P052nsss(0) <='1';
          else
          cVar2S24S37P066P036P052nsss(0) <='0';
          end if;
        if(cVar1S25S37P065N060P062P063(0)='1' AND  D( 0)='1' AND B( 9)='0' AND E( 8)='1' )then
          cVar2S25S37P066N036P069nsss(0) <='1';
          else
          cVar2S25S37P066N036P069nsss(0) <='0';
          end if;
        if(cVar1S26S37P065N060P062N063(0)='1' AND  A(10)='1' AND E(11)='1' )then
          cVar2S26S37P018P057nsss(0) <='1';
          else
          cVar2S26S37P018P057nsss(0) <='0';
          end if;
        if(cVar1S27S37P065N060P062N063(0)='1' AND  A(10)='1' AND E(11)='0' AND A( 2)='1' )then
          cVar2S27S37P018N057P015nsss(0) <='1';
          else
          cVar2S27S37P018N057P015nsss(0) <='0';
          end if;
        if(cVar1S28S37P065N060P062N063(0)='1' AND  A(10)='0' AND A(19)='1' )then
          cVar2S28S37N018P000nsss(0) <='1';
          else
          cVar2S28S37N018P000nsss(0) <='0';
          end if;
        if(cVar1S29S37P065N060P062P063(0)='1' AND  A( 1)='1' AND A(10)='1' )then
          cVar2S29S37P017P018nsss(0) <='1';
          else
          cVar2S29S37P017P018nsss(0) <='0';
          end if;
        if(cVar1S30S37P065N060P062P063(0)='1' AND  A( 1)='1' AND A(10)='0' AND B( 0)='1' )then
          cVar2S30S37P017N018P037nsss(0) <='1';
          else
          cVar2S30S37P017N018P037nsss(0) <='0';
          end if;
        if(cVar1S31S37P065N060P062P063(0)='1' AND  A( 1)='0' AND E( 0)='1' )then
          cVar2S31S37N017P068nsss(0) <='1';
          else
          cVar2S31S37N017P068nsss(0) <='0';
          end if;
        if(cVar1S32S37P065N060P062P063(0)='1' AND  A( 1)='0' AND E( 0)='0' AND A(10)='0' )then
          cVar2S32S37N017N068P018nsss(0) <='1';
          else
          cVar2S32S37N017N068P018nsss(0) <='0';
          end if;
        if(cVar1S33S37P065N060P062P063(0)='1' AND  D( 2)='0' AND E(14)='1' )then
          cVar2S33S37P058P045nsss(0) <='1';
          else
          cVar2S33S37P058P045nsss(0) <='0';
          end if;
        if(cVar1S0S38P019P069P015P006(0)='1' AND  B(15)='0' AND B( 4)='0' AND D( 3)='0' )then
          cVar2S0S38P024P029P054nsss(0) <='1';
          else
          cVar2S0S38P024P029P054nsss(0) <='0';
          end if;
        if(cVar1S1S38P019P069P015P006(0)='1' AND  B(15)='0' AND B( 4)='1' AND A(11)='0' )then
          cVar2S1S38P024P029P016nsss(0) <='1';
          else
          cVar2S1S38P024P029P016nsss(0) <='0';
          end if;
        if(cVar1S2S38P019P069P015P006(0)='1' AND  D( 1)='1' )then
          cVar2S2S38P062nsss(0) <='1';
          else
          cVar2S2S38P062nsss(0) <='0';
          end if;
        if(cVar1S3S38P019P069P015P006(0)='1' AND  D( 1)='0' AND A(15)='1' )then
          cVar2S3S38N062P008nsss(0) <='1';
          else
          cVar2S3S38N062P008nsss(0) <='0';
          end if;
        if(cVar1S4S38P019P069N015P009(0)='1' AND  E( 1)='1' )then
          cVar2S4S38P064nsss(0) <='1';
          else
          cVar2S4S38P064nsss(0) <='0';
          end if;
        if(cVar1S5S38P019P069N015P009(0)='1' AND  E( 1)='0' AND A( 8)='0' AND D( 9)='0' )then
          cVar2S5S38N064P003P063nsss(0) <='1';
          else
          cVar2S5S38N064P003P063nsss(0) <='0';
          end if;
        if(cVar1S6S38P019P069N015N009(0)='1' AND  D( 1)='0' AND D( 2)='0' )then
          cVar2S6S38P062P058nsss(0) <='1';
          else
          cVar2S6S38P062P058nsss(0) <='0';
          end if;
        if(cVar1S7S38P019P069N015N009(0)='1' AND  D( 1)='0' AND D( 2)='1' AND A(10)='0' )then
          cVar2S7S38P062P058P018nsss(0) <='1';
          else
          cVar2S7S38P062P058P018nsss(0) <='0';
          end if;
        if(cVar1S8S38P019P069N015N009(0)='1' AND  D( 1)='1' AND D( 8)='0' )then
          cVar2S8S38P062P067nsss(0) <='1';
          else
          cVar2S8S38P062P067nsss(0) <='0';
          end if;
        if(cVar1S9S38P019P069N015N009(0)='1' AND  D( 1)='1' AND D( 8)='1' AND E( 2)='1' )then
          cVar2S9S38P062P067P060nsss(0) <='1';
          else
          cVar2S9S38P062P067P060nsss(0) <='0';
          end if;
        if(cVar1S10S38P019N069P008P034(0)='1' AND  A( 4)='0' AND A(14)='0' AND B(13)='0' )then
          cVar2S10S38P011P010P028nsss(0) <='1';
          else
          cVar2S10S38P011P010P028nsss(0) <='0';
          end if;
        if(cVar1S11S38P019N069P008P034(0)='1' AND  A( 4)='0' AND A(14)='1' AND A( 1)='0' )then
          cVar2S11S38P011P010P017nsss(0) <='1';
          else
          cVar2S11S38P011P010P017nsss(0) <='0';
          end if;
        if(cVar1S12S38P019N069P008P034(0)='1' AND  A( 4)='1' AND B( 5)='1' )then
          cVar2S12S38P011P027nsss(0) <='1';
          else
          cVar2S12S38P011P027nsss(0) <='0';
          end if;
        if(cVar1S13S38P019N069P008P034(0)='1' AND  A( 4)='1' AND B( 5)='0' AND B( 0)='0' )then
          cVar2S13S38P011N027P037nsss(0) <='1';
          else
          cVar2S13S38P011N027P037nsss(0) <='0';
          end if;
        if(cVar1S14S38P019N069P008P034(0)='1' AND  A( 6)='0' AND A( 4)='1' AND A(10)='0' )then
          cVar2S14S38P007P011P018nsss(0) <='1';
          else
          cVar2S14S38P007P011P018nsss(0) <='0';
          end if;
        if(cVar1S15S38P019N069N008P016(0)='1' AND  E(10)='0' AND A( 2)='0' AND E(12)='0' )then
          cVar2S15S38P061P015P053nsss(0) <='1';
          else
          cVar2S15S38P061P015P053nsss(0) <='0';
          end if;
        if(cVar1S16S38P019N069N008P016(0)='1' AND  E(10)='0' AND A( 2)='1' AND B( 7)='1' )then
          cVar2S16S38P061P015P023nsss(0) <='1';
          else
          cVar2S16S38P061P015P023nsss(0) <='0';
          end if;
        if(cVar1S17S38P019N069N008P016(0)='1' AND  E(10)='1' AND A( 1)='1' AND B(10)='0' )then
          cVar2S17S38P061P017P034nsss(0) <='1';
          else
          cVar2S17S38P061P017P034nsss(0) <='0';
          end if;
        if(cVar1S18S38P019N069N008N016(0)='1' AND  A( 2)='1' AND E(10)='1' AND B(11)='0' )then
          cVar2S18S38P015P061P032nsss(0) <='1';
          else
          cVar2S18S38P015P061P032nsss(0) <='0';
          end if;
        if(cVar1S19S38P019N069N008N016(0)='1' AND  A( 2)='1' AND E(10)='0' AND A(10)='0' )then
          cVar2S19S38P015N061P018nsss(0) <='1';
          else
          cVar2S19S38P015N061P018nsss(0) <='0';
          end if;
        if(cVar1S20S38P019N069N008N016(0)='1' AND  A( 2)='0' AND A(13)='1' AND A( 1)='1' )then
          cVar2S20S38N015P012P017nsss(0) <='1';
          else
          cVar2S20S38N015P012P017nsss(0) <='0';
          end if;
        if(cVar1S21S38N019P069P033P003(0)='1' AND  E( 3)='1' AND E(11)='0' AND A(11)='0' )then
          cVar2S21S38P056P057P016nsss(0) <='1';
          else
          cVar2S21S38P056P057P016nsss(0) <='0';
          end if;
        if(cVar1S22S38N019P069P033P003(0)='1' AND  E( 3)='1' AND E(11)='1' AND B( 3)='1' )then
          cVar2S22S38P056P057P031nsss(0) <='1';
          else
          cVar2S22S38P056P057P031nsss(0) <='0';
          end if;
        if(cVar1S23S38N019P069P033P003(0)='1' AND  E( 3)='0' AND A(10)='1' )then
          cVar2S23S38N056P018nsss(0) <='1';
          else
          cVar2S23S38N056P018nsss(0) <='0';
          end if;
        if(cVar1S24S38N019P069P033P003(0)='1' AND  E( 3)='0' AND A(10)='0' AND B(11)='0' )then
          cVar2S24S38N056N018P032nsss(0) <='1';
          else
          cVar2S24S38N056N018P032nsss(0) <='0';
          end if;
        if(cVar1S25S38N019P069P033P003(0)='1' AND  D( 0)='0' AND A( 6)='0' AND A( 1)='1' )then
          cVar2S25S38P066P007P017nsss(0) <='1';
          else
          cVar2S25S38P066P007P017nsss(0) <='0';
          end if;
        if(cVar1S26S38N019P069N033P041(0)='1' AND  B(17)='1' AND A( 7)='1' )then
          cVar2S26S38P020P005nsss(0) <='1';
          else
          cVar2S26S38P020P005nsss(0) <='0';
          end if;
        if(cVar1S27S38N019P069N033P041(0)='1' AND  B(17)='1' AND A( 7)='0' AND E( 7)='0' )then
          cVar2S27S38P020N005P040nsss(0) <='1';
          else
          cVar2S27S38P020N005P040nsss(0) <='0';
          end if;
        if(cVar1S28S38N019P069N033P041(0)='1' AND  B(17)='0' AND A( 3)='0' AND D( 1)='0' )then
          cVar2S28S38N020P013P062nsss(0) <='1';
          else
          cVar2S28S38N020P013P062nsss(0) <='0';
          end if;
        if(cVar1S29S38N019P069N033N041(0)='1' AND  A( 4)='1' AND E( 2)='1' AND B(13)='0' )then
          cVar2S29S38P011P060P028nsss(0) <='1';
          else
          cVar2S29S38P011P060P028nsss(0) <='0';
          end if;
        if(cVar1S30S38N019P069N033N041(0)='1' AND  A( 4)='1' AND E( 2)='0' )then
          cVar2S30S38P011N060psss(0) <='1';
          else
          cVar2S30S38P011N060psss(0) <='0';
          end if;
        if(cVar1S31S38N019P069N033N041(0)='1' AND  A( 4)='0' AND B(15)='1' AND B(14)='0' )then
          cVar2S31S38N011P024P026nsss(0) <='1';
          else
          cVar2S31S38N011P024P026nsss(0) <='0';
          end if;
        if(cVar1S32S38N019P069P058P054(0)='1' AND  E( 1)='0' AND A( 2)='0' )then
          cVar2S32S38P064P015nsss(0) <='1';
          else
          cVar2S32S38P064P015nsss(0) <='0';
          end if;
        if(cVar1S33S38N019P069P058P054(0)='1' AND  E( 1)='0' AND A( 2)='1' AND D(10)='0' )then
          cVar2S33S38P064P015P059nsss(0) <='1';
          else
          cVar2S33S38P064P015P059nsss(0) <='0';
          end if;
        if(cVar1S34S38N019P069P058P054(0)='1' AND  E( 1)='1' AND E( 9)='1' )then
          cVar2S34S38P064P065nsss(0) <='1';
          else
          cVar2S34S38P064P065nsss(0) <='0';
          end if;
        if(cVar1S35S38N019P069N058P011(0)='1' AND  D( 3)='1' AND B( 9)='0' )then
          cVar2S35S38P054P036nsss(0) <='1';
          else
          cVar2S35S38P054P036nsss(0) <='0';
          end if;
        if(cVar1S36S38N019P069N058P011(0)='1' AND  D( 3)='1' AND B( 9)='1' AND A(10)='0' )then
          cVar2S36S38P054P036P018nsss(0) <='1';
          else
          cVar2S36S38P054P036P018nsss(0) <='0';
          end if;
        if(cVar1S37S38N019P069N058P011(0)='1' AND  E( 9)='1' AND D( 9)='1' AND A( 1)='1' )then
          cVar2S37S38P065P063P017nsss(0) <='1';
          else
          cVar2S37S38P065P063P017nsss(0) <='0';
          end if;
        if(cVar1S38S38N019P069N058P011(0)='1' AND  E( 9)='0' AND B( 1)='0' AND A(14)='1' )then
          cVar2S38S38N065P035P010nsss(0) <='1';
          else
          cVar2S38S38N065P035P010nsss(0) <='0';
          end if;
        if(cVar1S0S39P011P069P058P067(0)='1' AND  A( 0)='0' AND D(10)='1' AND A( 5)='0' )then
          cVar2S0S39P019P059P009nsss(0) <='1';
          else
          cVar2S0S39P019P059P009nsss(0) <='0';
          end if;
        if(cVar1S1S39P011P069P058P067(0)='1' AND  A( 0)='0' AND D(10)='0' AND B( 2)='0' )then
          cVar2S1S39P019N059P033nsss(0) <='1';
          else
          cVar2S1S39P019N059P033nsss(0) <='0';
          end if;
        if(cVar1S2S39P011P069P058P067(0)='1' AND  A( 0)='1' AND E( 0)='1' AND B(11)='0' )then
          cVar2S2S39P019P068P032nsss(0) <='1';
          else
          cVar2S2S39P019P068P032nsss(0) <='0';
          end if;
        if(cVar1S3S39P011P069P058P067(0)='1' AND  A( 0)='1' AND E( 0)='0' AND E( 9)='1' )then
          cVar2S3S39P019N068P065nsss(0) <='1';
          else
          cVar2S3S39P019N068P065nsss(0) <='0';
          end if;
        if(cVar1S4S39P011P069P058P067(0)='1' AND  E( 0)='1' AND E( 9)='0' AND B( 0)='1' )then
          cVar2S4S39P068P065P037nsss(0) <='1';
          else
          cVar2S4S39P068P065P037nsss(0) <='0';
          end if;
        if(cVar1S5S39P011P069P058P067(0)='1' AND  E( 0)='1' AND E( 9)='1' AND B( 9)='0' )then
          cVar2S5S39P068P065P036nsss(0) <='1';
          else
          cVar2S5S39P068P065P036nsss(0) <='0';
          end if;
        if(cVar1S6S39P011P069P058P067(0)='1' AND  E( 0)='0' AND D(13)='1' )then
          cVar2S6S39N068P047nsss(0) <='1';
          else
          cVar2S6S39N068P047nsss(0) <='0';
          end if;
        if(cVar1S7S39P011P069P058P067(0)='1' AND  E( 0)='0' AND D(13)='0' AND E(14)='1' )then
          cVar2S7S39N068N047P045nsss(0) <='1';
          else
          cVar2S7S39N068N047P045nsss(0) <='0';
          end if;
        if(cVar1S8S39P011P069P058P062(0)='1' AND  E( 3)='1' AND E(11)='0' )then
          cVar2S8S39P056P057nsss(0) <='1';
          else
          cVar2S8S39P056P057nsss(0) <='0';
          end if;
        if(cVar1S9S39P011P069P058P062(0)='1' AND  E( 3)='1' AND E(11)='1' AND A(12)='0' )then
          cVar2S9S39P056P057P014nsss(0) <='1';
          else
          cVar2S9S39P056P057P014nsss(0) <='0';
          end if;
        if(cVar1S10S39P011P069P058P062(0)='1' AND  E( 3)='0' AND D( 3)='0' AND E( 2)='1' )then
          cVar2S10S39N056P054P060nsss(0) <='1';
          else
          cVar2S10S39N056P054P060nsss(0) <='0';
          end if;
        if(cVar1S11S39P011P069P058P062(0)='1' AND  A( 2)='1' AND B( 1)='1' AND B(10)='0' )then
          cVar2S11S39P015P035P034nsss(0) <='1';
          else
          cVar2S11S39P015P035P034nsss(0) <='0';
          end if;
        if(cVar1S12S39P011P069P058P062(0)='1' AND  A( 2)='1' AND B( 1)='0' AND A(11)='1' )then
          cVar2S12S39P015N035P016nsss(0) <='1';
          else
          cVar2S12S39P015N035P016nsss(0) <='0';
          end if;
        if(cVar1S13S39P011P069P017P068(0)='1' AND  B( 0)='0' AND A(10)='1' AND B( 2)='0' )then
          cVar2S13S39P037P018P033nsss(0) <='1';
          else
          cVar2S13S39P037P018P033nsss(0) <='0';
          end if;
        if(cVar1S14S39P011P069P017P068(0)='1' AND  B( 0)='0' AND A(10)='0' AND A(12)='0' )then
          cVar2S14S39P037N018P014nsss(0) <='1';
          else
          cVar2S14S39P037N018P014nsss(0) <='0';
          end if;
        if(cVar1S15S39P011P069P017P068(0)='1' AND  B( 0)='1' AND B( 9)='0' AND A(10)='0' )then
          cVar2S15S39P037P036P018nsss(0) <='1';
          else
          cVar2S15S39P037P036P018nsss(0) <='0';
          end if;
        if(cVar1S16S39P011P069P017P068(0)='1' AND  B( 0)='1' AND B( 9)='1' AND A(13)='1' )then
          cVar2S16S39P037P036P012nsss(0) <='1';
          else
          cVar2S16S39P037P036P012nsss(0) <='0';
          end if;
        if(cVar1S17S39P011P069P017N068(0)='1' AND  D( 5)='1' AND A(10)='0' )then
          cVar2S17S39P046P018nsss(0) <='1';
          else
          cVar2S17S39P046P018nsss(0) <='0';
          end if;
        if(cVar1S18S39P011P069P017N068(0)='1' AND  D( 5)='0' AND A( 2)='0' AND B( 2)='1' )then
          cVar2S18S39N046P015P033nsss(0) <='1';
          else
          cVar2S18S39N046P015P033nsss(0) <='0';
          end if;
        if(cVar1S19S39P011P069N017P047(0)='1' AND  D( 9)='0' )then
          cVar2S19S39P063nsss(0) <='1';
          else
          cVar2S19S39P063nsss(0) <='0';
          end if;
        if(cVar1S20S39P011P069N017N047(0)='1' AND  D( 8)='1' AND A( 9)='1' )then
          cVar2S20S39P067P001nsss(0) <='1';
          else
          cVar2S20S39P067P001nsss(0) <='0';
          end if;
        if(cVar1S21S39P011P069N017N047(0)='1' AND  D( 8)='0' AND A( 0)='1' AND D( 0)='1' )then
          cVar2S21S39N067P019P066nsss(0) <='1';
          else
          cVar2S21S39N067P019P066nsss(0) <='0';
          end if;
        if(cVar1S22S39P011P019P062P015(0)='1' AND  E(11)='1' )then
          cVar2S22S39P057nsss(0) <='1';
          else
          cVar2S22S39P057nsss(0) <='0';
          end if;
        if(cVar1S23S39P011P019P062P015(0)='1' AND  E(11)='0' AND B( 9)='1' )then
          cVar2S23S39N057P036nsss(0) <='1';
          else
          cVar2S23S39N057P036nsss(0) <='0';
          end if;
        if(cVar1S24S39P011P019P062P015(0)='1' AND  E(11)='0' AND B( 9)='0' AND A( 1)='1' )then
          cVar2S24S39N057N036P017nsss(0) <='1';
          else
          cVar2S24S39N057N036P017nsss(0) <='0';
          end if;
        if(cVar1S25S39P011P019P062P015(0)='1' AND  A( 5)='0' AND E( 8)='1' )then
          cVar2S25S39P009P069nsss(0) <='1';
          else
          cVar2S25S39P009P069nsss(0) <='0';
          end if;
        if(cVar1S26S39P011P019P062P015(0)='1' AND  A( 5)='0' AND E( 8)='0' AND B( 0)='0' )then
          cVar2S26S39P009N069P037nsss(0) <='1';
          else
          cVar2S26S39P009N069P037nsss(0) <='0';
          end if;
        if(cVar1S27S39P011P019P062P015(0)='1' AND  A( 5)='1' AND A(10)='0' AND D( 0)='0' )then
          cVar2S27S39P009P018P066nsss(0) <='1';
          else
          cVar2S27S39P009P018P066nsss(0) <='0';
          end if;
        if(cVar1S28S39P011P019N062P064(0)='1' AND  B( 0)='1' AND E( 8)='1' )then
          cVar2S28S39P037P069nsss(0) <='1';
          else
          cVar2S28S39P037P069nsss(0) <='0';
          end if;
        if(cVar1S29S39P011P019N062P064(0)='1' AND  B( 0)='1' AND E( 8)='0' AND D(11)='1' )then
          cVar2S29S39P037N069P055nsss(0) <='1';
          else
          cVar2S29S39P037N069P055nsss(0) <='0';
          end if;
        if(cVar1S30S39P011P019N062P064(0)='1' AND  B( 0)='0' AND E(10)='1' AND A(12)='0' )then
          cVar2S30S39N037P061P014nsss(0) <='1';
          else
          cVar2S30S39N037P061P014nsss(0) <='0';
          end if;
        if(cVar1S31S39P011P019N062P064(0)='1' AND  A(12)='0' AND A( 2)='0' AND B( 0)='1' )then
          cVar2S31S39P014P015P037nsss(0) <='1';
          else
          cVar2S31S39P014P015P037nsss(0) <='0';
          end if;
        if(cVar1S32S39P011N019P060P061(0)='1' AND  B(10)='1' )then
          cVar2S32S39P034nsss(0) <='1';
          else
          cVar2S32S39P034nsss(0) <='0';
          end if;
        if(cVar1S33S39P011N019P060P061(0)='1' AND  B(10)='0' AND A(10)='1' )then
          cVar2S33S39N034P018nsss(0) <='1';
          else
          cVar2S33S39N034P018nsss(0) <='0';
          end if;
        if(cVar1S34S39P011N019P060P061(0)='1' AND  B(10)='0' AND A(10)='0' AND B(11)='0' )then
          cVar2S34S39N034N018P032nsss(0) <='1';
          else
          cVar2S34S39N034N018P032nsss(0) <='0';
          end if;
        if(cVar1S35S39P011N019P060N061(0)='1' AND  B(14)='0' AND E(11)='1' )then
          cVar2S35S39P026P057nsss(0) <='1';
          else
          cVar2S35S39P026P057nsss(0) <='0';
          end if;
        if(cVar1S36S39P011N019P060N061(0)='1' AND  B(14)='0' AND E(11)='0' AND D( 9)='1' )then
          cVar2S36S39P026N057P063nsss(0) <='1';
          else
          cVar2S36S39P026N057P063nsss(0) <='0';
          end if;
        if(cVar1S37S39P011N019N060P049(0)='1' AND  B(14)='1' )then
          cVar2S37S39P026nsss(0) <='1';
          else
          cVar2S37S39P026nsss(0) <='0';
          end if;
        if(cVar1S38S39P011N019N060P049(0)='1' AND  B(14)='0' AND D( 0)='0' )then
          cVar2S38S39N026P066nsss(0) <='1';
          else
          cVar2S38S39N026P066nsss(0) <='0';
          end if;
        if(cVar1S39S39P011N019N060N049(0)='1' AND  D( 8)='0' AND D( 3)='1' AND B(11)='0' )then
          cVar2S39S39P067P054P032nsss(0) <='1';
          else
          cVar2S39S39P067P054P032nsss(0) <='0';
          end if;
        if(cVar1S40S39P011N019N060N049(0)='1' AND  D( 8)='1' AND D(11)='1' AND A(10)='1' )then
          cVar2S40S39P067P055P018nsss(0) <='1';
          else
          cVar2S40S39P067P055P018nsss(0) <='0';
          end if;
        if(cVar1S0S40P069P053P067P011(0)='1' AND  D( 2)='0' )then
          cVar2S0S40P058nsss(0) <='1';
          else
          cVar2S0S40P058nsss(0) <='0';
          end if;
        if(cVar1S1S40P069P053P067P011(0)='1' AND  D( 2)='1' AND A(13)='1' AND E( 9)='0' )then
          cVar2S1S40P058P012P065nsss(0) <='1';
          else
          cVar2S1S40P058P012P065nsss(0) <='0';
          end if;
        if(cVar1S2S40P069P053P067P011(0)='1' AND  D( 2)='1' AND A(13)='0' AND D( 9)='1' )then
          cVar2S2S40P058N012P063nsss(0) <='1';
          else
          cVar2S2S40P058N012P063nsss(0) <='0';
          end if;
        if(cVar1S3S40P069P053P067P011(0)='1' AND  A( 0)='1' AND D(13)='0' )then
          cVar2S3S40P019P047nsss(0) <='1';
          else
          cVar2S3S40P019P047nsss(0) <='0';
          end if;
        if(cVar1S4S40P069P053P067P011(0)='1' AND  A( 0)='0' AND D( 9)='1' )then
          cVar2S4S40N019P063nsss(0) <='1';
          else
          cVar2S4S40N019P063nsss(0) <='0';
          end if;
        if(cVar1S5S40P069P053N067P064(0)='1' AND  E( 0)='0' AND D( 9)='1' )then
          cVar2S5S40P068P063nsss(0) <='1';
          else
          cVar2S5S40P068P063nsss(0) <='0';
          end if;
        if(cVar1S6S40P069P053N067P064(0)='1' AND  E( 0)='0' AND D( 9)='0' AND A( 3)='1' )then
          cVar2S6S40P068N063P013nsss(0) <='1';
          else
          cVar2S6S40P068N063P013nsss(0) <='0';
          end if;
        if(cVar1S7S40P069P053N067P064(0)='1' AND  E( 0)='1' AND B( 0)='1' )then
          cVar2S7S40P068P037nsss(0) <='1';
          else
          cVar2S7S40P068P037nsss(0) <='0';
          end if;
        if(cVar1S8S40P069P053N067N064(0)='1' AND  E( 0)='1' AND A( 1)='1' )then
          cVar2S8S40P068P017nsss(0) <='1';
          else
          cVar2S8S40P068P017nsss(0) <='0';
          end if;
        if(cVar1S9S40P069P053N067N064(0)='1' AND  E( 0)='1' AND A( 1)='0' AND A( 0)='1' )then
          cVar2S9S40P068N017P019nsss(0) <='1';
          else
          cVar2S9S40P068N017P019nsss(0) <='0';
          end if;
        if(cVar1S10S40P069P053N067N064(0)='1' AND  E( 0)='0' AND E( 2)='1' AND E( 9)='1' )then
          cVar2S10S40N068P060P065nsss(0) <='1';
          else
          cVar2S10S40N068P060P065nsss(0) <='0';
          end if;
        if(cVar1S11S40P069P053N067N064(0)='1' AND  E( 0)='0' AND E( 2)='0' AND E( 4)='1' )then
          cVar2S11S40N068N060P052nsss(0) <='1';
          else
          cVar2S11S40N068N060P052nsss(0) <='0';
          end if;
        if(cVar1S13S40P069P053P059N060(0)='1' AND  E(11)='0' AND A(16)='0' AND D( 3)='1' )then
          cVar2S13S40P057P006P054nsss(0) <='1';
          else
          cVar2S13S40P057P006P054nsss(0) <='0';
          end if;
        if(cVar1S14S40N069P031P013P065(0)='1' AND  B(12)='0' AND D(10)='0' )then
          cVar2S14S40P030P059nsss(0) <='1';
          else
          cVar2S14S40P030P059nsss(0) <='0';
          end if;
        if(cVar1S15S40N069P031P013P065(0)='1' AND  B(12)='0' AND D(10)='1' AND A(13)='1' )then
          cVar2S15S40P030P059P012nsss(0) <='1';
          else
          cVar2S15S40P030P059P012nsss(0) <='0';
          end if;
        if(cVar1S16S40N069P031P013P065(0)='1' AND  B(12)='1' AND A( 4)='0' AND A(14)='1' )then
          cVar2S16S40P030P011P010nsss(0) <='1';
          else
          cVar2S16S40P030P011P010nsss(0) <='0';
          end if;
        if(cVar1S17S40N069P031P013P065(0)='1' AND  A( 4)='1' )then
          cVar2S17S40P011nsss(0) <='1';
          else
          cVar2S17S40P011nsss(0) <='0';
          end if;
        if(cVar1S18S40N069P031P013P065(0)='1' AND  A( 4)='0' AND E( 3)='0' AND E(11)='1' )then
          cVar2S18S40N011P056P057nsss(0) <='1';
          else
          cVar2S18S40N011P056P057nsss(0) <='0';
          end if;
        if(cVar1S19S40N069P031P013P065(0)='1' AND  A( 4)='0' AND E( 3)='1' AND A(10)='1' )then
          cVar2S19S40N011P056P018nsss(0) <='1';
          else
          cVar2S19S40N011P056P018nsss(0) <='0';
          end if;
        if(cVar1S20S40N069P031N013P058(0)='1' AND  B( 2)='0' )then
          cVar2S20S40P033nsss(0) <='1';
          else
          cVar2S20S40P033nsss(0) <='0';
          end if;
        if(cVar1S21S40N069P031N013P058(0)='1' AND  B( 2)='1' AND D( 3)='1' )then
          cVar2S21S40P033P054nsss(0) <='1';
          else
          cVar2S21S40P033P054nsss(0) <='0';
          end if;
        if(cVar1S22S40N069P031N013N058(0)='1' AND  D( 3)='1' AND B( 1)='1' )then
          cVar2S22S40P054P035nsss(0) <='1';
          else
          cVar2S22S40P054P035nsss(0) <='0';
          end if;
        if(cVar1S23S40N069P031N013N058(0)='1' AND  D( 3)='0' AND A( 4)='1' AND A(12)='0' )then
          cVar2S23S40N054P011P014nsss(0) <='1';
          else
          cVar2S23S40N054P011P014nsss(0) <='0';
          end if;
        if(cVar1S24S40N069P031N013N058(0)='1' AND  D( 3)='0' AND A( 4)='0' AND B( 4)='1' )then
          cVar2S24S40N054N011P029nsss(0) <='1';
          else
          cVar2S24S40N054N011P029nsss(0) <='0';
          end if;
        if(cVar1S25S40N069N031P030P061(0)='1' AND  A( 3)='1' )then
          cVar2S25S40P013nsss(0) <='1';
          else
          cVar2S25S40P013nsss(0) <='0';
          end if;
        if(cVar1S26S40N069N031P030P061(0)='1' AND  A( 3)='0' AND D( 1)='0' )then
          cVar2S26S40N013P062nsss(0) <='1';
          else
          cVar2S26S40N013P062nsss(0) <='0';
          end if;
        if(cVar1S27S40N069N031P030N061(0)='1' AND  E(14)='1' )then
          cVar2S27S40P045nsss(0) <='1';
          else
          cVar2S27S40P045nsss(0) <='0';
          end if;
        if(cVar1S28S40N069N031P030N061(0)='1' AND  E(14)='0' AND E( 1)='0' AND A( 3)='0' )then
          cVar2S28S40N045P064P013nsss(0) <='1';
          else
          cVar2S28S40N045P064P013nsss(0) <='0';
          end if;
        if(cVar1S29S40N069N031P030N061(0)='1' AND  E(14)='0' AND E( 1)='1' AND B( 0)='1' )then
          cVar2S29S40N045P064P037nsss(0) <='1';
          else
          cVar2S29S40N045P064P037nsss(0) <='0';
          end if;
        if(cVar1S30S40N069N031N030P000(0)='1' AND  D( 2)='0' AND A( 3)='0' AND B(14)='1' )then
          cVar2S30S40P058P013P026nsss(0) <='1';
          else
          cVar2S30S40P058P013P026nsss(0) <='0';
          end if;
        if(cVar1S31S40N069N031N030P000(0)='1' AND  D( 2)='0' AND A( 3)='1' AND D(10)='1' )then
          cVar2S31S40P058P013P059nsss(0) <='1';
          else
          cVar2S31S40P058P013P059nsss(0) <='0';
          end if;
        if(cVar1S32S40N069N031N030P000(0)='1' AND  D( 2)='1' AND A(12)='1' AND A(11)='0' )then
          cVar2S32S40P058P014P016nsss(0) <='1';
          else
          cVar2S32S40P058P014P016nsss(0) <='0';
          end if;
        if(cVar1S33S40N069N031N030P000(0)='1' AND  D( 1)='1' AND B( 1)='1' )then
          cVar2S33S40P062P035nsss(0) <='1';
          else
          cVar2S33S40P062P035nsss(0) <='0';
          end if;
        if(cVar1S34S40N069N031N030P000(0)='1' AND  D( 1)='1' AND B( 1)='0' AND B( 2)='1' )then
          cVar2S34S40P062N035P033nsss(0) <='1';
          else
          cVar2S34S40P062N035P033nsss(0) <='0';
          end if;
        if(cVar1S35S40N069N031N030P000(0)='1' AND  D( 1)='0' AND D(10)='1' AND A( 2)='1' )then
          cVar2S35S40N062P059P015nsss(0) <='1';
          else
          cVar2S35S40N062P059P015nsss(0) <='0';
          end if;
        if(cVar1S36S40N069N031N030P000(0)='1' AND  D( 1)='0' AND D(10)='0' AND B(17)='1' )then
          cVar2S36S40N062N059P020nsss(0) <='1';
          else
          cVar2S36S40N062N059P020nsss(0) <='0';
          end if;
        if(cVar1S2S41P025N004P007P067(0)='1' AND  E( 9)='0' AND A( 8)='0' )then
          cVar2S2S41P065P003nsss(0) <='1';
          else
          cVar2S2S41P065P003nsss(0) <='0';
          end if;
        if(cVar1S3S41P025N004P007P067(0)='1' AND  E( 9)='1' AND A(11)='0' )then
          cVar2S3S41P065P016nsss(0) <='1';
          else
          cVar2S3S41P065P016nsss(0) <='0';
          end if;
        if(cVar1S4S41P025N004P007P067(0)='1' AND  E( 6)='0' AND B( 9)='1' )then
          cVar2S4S41P044P036nsss(0) <='1';
          else
          cVar2S4S41P044P036nsss(0) <='0';
          end if;
        if(cVar1S5S41P025N004N007P037(0)='1' AND  A( 2)='1' AND A(11)='0' )then
          cVar2S5S41P015P016nsss(0) <='1';
          else
          cVar2S5S41P015P016nsss(0) <='0';
          end if;
        if(cVar1S6S41P025N004N007P037(0)='1' AND  A( 2)='0' AND A( 1)='1' )then
          cVar2S6S41N015P017nsss(0) <='1';
          else
          cVar2S6S41N015P017nsss(0) <='0';
          end if;
        if(cVar1S7S41P025N004N007N037(0)='1' AND  B( 2)='1' AND A(13)='0' )then
          cVar2S7S41P033P012nsss(0) <='1';
          else
          cVar2S7S41P033P012nsss(0) <='0';
          end if;
        if(cVar1S8S41P025N004N007N037(0)='1' AND  B( 2)='0' AND A(16)='1' )then
          cVar2S8S41N033P006nsss(0) <='1';
          else
          cVar2S8S41N033P006nsss(0) <='0';
          end if;
        if(cVar1S9S41P025N004N007N037(0)='1' AND  B( 2)='0' AND A(16)='0' AND A( 5)='1' )then
          cVar2S9S41N033N006P009nsss(0) <='1';
          else
          cVar2S9S41N033N006P009nsss(0) <='0';
          end if;
        if(cVar1S10S41N025P062P058P055(0)='1' AND  D( 8)='0' AND A(16)='0' )then
          cVar2S10S41P067P006nsss(0) <='1';
          else
          cVar2S10S41P067P006nsss(0) <='0';
          end if;
        if(cVar1S11S41N025P062P058P055(0)='1' AND  D( 8)='0' AND A(16)='1' AND E( 3)='1' )then
          cVar2S11S41P067P006P056nsss(0) <='1';
          else
          cVar2S11S41P067P006P056nsss(0) <='0';
          end if;
        if(cVar1S12S41N025P062P058P055(0)='1' AND  D( 8)='1' AND D( 5)='0' AND A(10)='0' )then
          cVar2S12S41P067P046P018nsss(0) <='1';
          else
          cVar2S12S41P067P046P018nsss(0) <='0';
          end if;
        if(cVar1S13S41N025P062P058P055(0)='1' AND  A( 3)='1' AND B( 3)='1' AND D( 3)='0' )then
          cVar2S13S41P013P031P054nsss(0) <='1';
          else
          cVar2S13S41P013P031P054nsss(0) <='0';
          end if;
        if(cVar1S14S41N025P062P058P055(0)='1' AND  A( 3)='1' AND B( 3)='0' AND A(10)='0' )then
          cVar2S14S41P013N031P018nsss(0) <='1';
          else
          cVar2S14S41P013N031P018nsss(0) <='0';
          end if;
        if(cVar1S15S41N025P062P058P055(0)='1' AND  A( 3)='0' AND E( 0)='1' )then
          cVar2S15S41N013P068nsss(0) <='1';
          else
          cVar2S15S41N013P068nsss(0) <='0';
          end if;
        if(cVar1S16S41N025P062P058P055(0)='1' AND  A( 3)='0' AND E( 0)='0' AND E( 3)='1' )then
          cVar2S16S41N013N068P056nsss(0) <='1';
          else
          cVar2S16S41N013N068P056nsss(0) <='0';
          end if;
        if(cVar1S17S41N025P062P058P049(0)='1' AND  E( 5)='0' AND D( 9)='1' AND D(10)='1' )then
          cVar2S17S41P048P063P059nsss(0) <='1';
          else
          cVar2S17S41P048P063P059nsss(0) <='0';
          end if;
        if(cVar1S18S41N025P062P058P049(0)='1' AND  E( 5)='0' AND D( 9)='0' AND B( 1)='1' )then
          cVar2S18S41P048N063P035nsss(0) <='1';
          else
          cVar2S18S41P048N063P035nsss(0) <='0';
          end if;
        if(cVar1S19S41N025N062P027P026(0)='1' AND  D( 5)='1' AND A(15)='1' )then
          cVar2S19S41P046P008nsss(0) <='1';
          else
          cVar2S19S41P046P008nsss(0) <='0';
          end if;
        if(cVar1S20S41N025N062P027P026(0)='1' AND  D( 5)='1' AND A(15)='0' AND B( 9)='1' )then
          cVar2S20S41P046N008P036nsss(0) <='1';
          else
          cVar2S20S41P046N008P036nsss(0) <='0';
          end if;
        if(cVar1S21S41N025N062P027P026(0)='1' AND  D( 5)='0' AND E( 8)='0' )then
          cVar2S21S41N046P069nsss(0) <='1';
          else
          cVar2S21S41N046P069nsss(0) <='0';
          end if;
        if(cVar1S22S41N025N062P027P026(0)='1' AND  D( 5)='0' AND E( 8)='1' AND E( 5)='0' )then
          cVar2S22S41N046P069P048nsss(0) <='1';
          else
          cVar2S22S41N046P069P048nsss(0) <='0';
          end if;
        if(cVar1S23S41N025N062P027P026(0)='1' AND  A( 5)='1' )then
          cVar2S23S41P009nsss(0) <='1';
          else
          cVar2S23S41P009nsss(0) <='0';
          end if;
        if(cVar1S24S41N025N062N027P048(0)='1' AND  E( 3)='1' AND B( 2)='1' AND A(15)='0' )then
          cVar2S24S41P056P033P008nsss(0) <='1';
          else
          cVar2S24S41P056P033P008nsss(0) <='0';
          end if;
        if(cVar1S25S41N025N062N027P048(0)='1' AND  E( 3)='1' AND B( 2)='0' AND D( 3)='1' )then
          cVar2S25S41P056N033P054nsss(0) <='1';
          else
          cVar2S25S41P056N033P054nsss(0) <='0';
          end if;
        if(cVar1S26S41N025N062N027P048(0)='1' AND  E( 3)='0' AND E( 0)='1' AND E( 1)='0' )then
          cVar2S26S41N056P068P064nsss(0) <='1';
          else
          cVar2S26S41N056P068P064nsss(0) <='0';
          end if;
        if(cVar1S27S41N025N062N027P048(0)='1' AND  E( 3)='0' AND E( 0)='0' AND D(11)='1' )then
          cVar2S27S41N056N068P055nsss(0) <='1';
          else
          cVar2S27S41N056N068P055nsss(0) <='0';
          end if;
        if(cVar1S28S41N025N062N027P048(0)='1' AND  E( 8)='1' AND A(14)='1' )then
          cVar2S28S41P069P010nsss(0) <='1';
          else
          cVar2S28S41P069P010nsss(0) <='0';
          end if;
        if(cVar1S29S41N025N062N027P048(0)='1' AND  E( 8)='1' AND A(14)='0' AND B(15)='1' )then
          cVar2S29S41P069N010P024nsss(0) <='1';
          else
          cVar2S29S41P069N010P024nsss(0) <='0';
          end if;
        if(cVar1S1S42P068P004P025N048(0)='1' AND  A(13)='0' )then
          cVar2S1S42P012nsss(0) <='1';
          else
          cVar2S1S42P012nsss(0) <='0';
          end if;
        if(cVar1S2S42P068P004N025P040(0)='1' AND  B( 8)='1' )then
          cVar2S2S42P021nsss(0) <='1';
          else
          cVar2S2S42P021nsss(0) <='0';
          end if;
        if(cVar1S3S42P068P004N025P040(0)='1' AND  B( 8)='0' AND B(17)='1' )then
          cVar2S3S42N021P020nsss(0) <='1';
          else
          cVar2S3S42N021P020nsss(0) <='0';
          end if;
        if(cVar1S4S42P068P004N025P040(0)='1' AND  B( 8)='0' AND B(17)='0' AND B( 7)='1' )then
          cVar2S4S42N021N020P023nsss(0) <='1';
          else
          cVar2S4S42N021N020P023nsss(0) <='0';
          end if;
        if(cVar1S5S42P068P004N025N040(0)='1' AND  E( 6)='1' )then
          cVar2S5S42P044nsss(0) <='1';
          else
          cVar2S5S42P044nsss(0) <='0';
          end if;
        if(cVar1S6S42P068P004N025N040(0)='1' AND  E( 6)='0' AND E( 5)='0' AND B(16)='1' )then
          cVar2S6S42N044P048P022nsss(0) <='1';
          else
          cVar2S6S42N044P048P022nsss(0) <='0';
          end if;
        if(cVar1S7S42P068N004P055P013(0)='1' AND  E(11)='0' )then
          cVar2S7S42P057nsss(0) <='1';
          else
          cVar2S7S42P057nsss(0) <='0';
          end if;
        if(cVar1S8S42P068N004P055P013(0)='1' AND  E(11)='1' AND B( 1)='1' AND D(10)='1' )then
          cVar2S8S42P057P035P059nsss(0) <='1';
          else
          cVar2S8S42P057P035P059nsss(0) <='0';
          end if;
        if(cVar1S9S42P068N004P055P013(0)='1' AND  D( 2)='1' AND A( 7)='0' )then
          cVar2S9S42P058P005nsss(0) <='1';
          else
          cVar2S9S42P058P005nsss(0) <='0';
          end if;
        if(cVar1S10S42P068N004P055P013(0)='1' AND  D( 2)='0' AND E( 4)='1' AND A(14)='1' )then
          cVar2S10S42N058P052P010nsss(0) <='1';
          else
          cVar2S10S42N058P052P010nsss(0) <='0';
          end if;
        if(cVar1S11S42P068N004P055P013(0)='1' AND  D( 2)='0' AND E( 4)='0' AND B(12)='1' )then
          cVar2S11S42N058N052P030nsss(0) <='1';
          else
          cVar2S11S42N058N052P030nsss(0) <='0';
          end if;
        if(cVar1S12S42P068N004P055P066(0)='1' AND  E(11)='1' AND A( 0)='1' AND B( 9)='0' )then
          cVar2S12S42P057P019P036nsss(0) <='1';
          else
          cVar2S12S42P057P019P036nsss(0) <='0';
          end if;
        if(cVar1S13S42P068N004P055P066(0)='1' AND  E(11)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar2S13S42P057N019P064nsss(0) <='1';
          else
          cVar2S13S42P057N019P064nsss(0) <='0';
          end if;
        if(cVar1S14S42P068N004P055P066(0)='1' AND  E(11)='0' AND E( 8)='1' AND E(10)='0' )then
          cVar2S14S42N057P069P061nsss(0) <='1';
          else
          cVar2S14S42N057P069P061nsss(0) <='0';
          end if;
        if(cVar1S15S42P068N004P055P066(0)='1' AND  E(11)='0' AND E( 8)='0' AND A(12)='1' )then
          cVar2S15S42N057N069P014nsss(0) <='1';
          else
          cVar2S15S42N057N069P014nsss(0) <='0';
          end if;
        if(cVar1S16S42P068N004P055P066(0)='1' AND  E( 9)='1' )then
          cVar2S16S42P065nsss(0) <='1';
          else
          cVar2S16S42P065nsss(0) <='0';
          end if;
        if(cVar1S17S42P068P015P061P069(0)='1' AND  B(11)='0' AND A( 6)='0' )then
          cVar2S17S42P032P007nsss(0) <='1';
          else
          cVar2S17S42P032P007nsss(0) <='0';
          end if;
        if(cVar1S18S42P068P015P061P069(0)='1' AND  B(11)='1' AND B( 0)='0' )then
          cVar2S18S42P032P037nsss(0) <='1';
          else
          cVar2S18S42P032P037nsss(0) <='0';
          end if;
        if(cVar1S19S42P068P015P061P069(0)='1' AND  B(11)='1' AND B( 0)='1' AND A(12)='1' )then
          cVar2S19S42P032P037P014nsss(0) <='1';
          else
          cVar2S19S42P032P037P014nsss(0) <='0';
          end if;
        if(cVar1S20S42P068P015P061P069(0)='1' AND  A(12)='1' )then
          cVar2S20S42P014nsss(0) <='1';
          else
          cVar2S20S42P014nsss(0) <='0';
          end if;
        if(cVar1S21S42P068P015P061P069(0)='1' AND  A(12)='0' AND A( 3)='1' )then
          cVar2S21S42N014P013nsss(0) <='1';
          else
          cVar2S21S42N014P013nsss(0) <='0';
          end if;
        if(cVar1S23S42P068P015N061N025(0)='1' AND  A(11)='1' AND B( 0)='1' AND A( 9)='0' )then
          cVar2S23S42P016P037P001nsss(0) <='1';
          else
          cVar2S23S42P016P037P001nsss(0) <='0';
          end if;
        if(cVar1S24S42P068P015N061N025(0)='1' AND  A(11)='1' AND B( 0)='0' AND B( 9)='1' )then
          cVar2S24S42P016N037P036nsss(0) <='1';
          else
          cVar2S24S42P016N037P036nsss(0) <='0';
          end if;
        if(cVar1S25S42P068P015N061N025(0)='1' AND  A(11)='0' AND D( 0)='1' AND E( 4)='1' )then
          cVar2S25S42N016P066P052nsss(0) <='1';
          else
          cVar2S25S42N016P066P052nsss(0) <='0';
          end if;
        if(cVar1S26S42P068N015P059P069(0)='1' AND  B( 2)='0' AND D( 9)='0' AND B( 9)='1' )then
          cVar2S26S42P033P063P036nsss(0) <='1';
          else
          cVar2S26S42P033P063P036nsss(0) <='0';
          end if;
        if(cVar1S27S42P068N015P059P069(0)='1' AND  B( 2)='1' AND B(10)='1' )then
          cVar2S27S42P033P034nsss(0) <='1';
          else
          cVar2S27S42P033P034nsss(0) <='0';
          end if;
        if(cVar1S28S42P068N015P059P069(0)='1' AND  A( 0)='0' AND D( 9)='1' AND A(15)='0' )then
          cVar2S28S42P019P063P008nsss(0) <='1';
          else
          cVar2S28S42P019P063P008nsss(0) <='0';
          end if;
        if(cVar1S29S42P068N015P059P069(0)='1' AND  A( 0)='1' AND A( 5)='1' )then
          cVar2S29S42P019P009nsss(0) <='1';
          else
          cVar2S29S42P019P009nsss(0) <='0';
          end if;
        if(cVar1S30S42P068N015P059P069(0)='1' AND  A( 0)='1' AND A( 5)='0' AND B( 2)='1' )then
          cVar2S30S42P019N009P033nsss(0) <='1';
          else
          cVar2S30S42P019N009P033nsss(0) <='0';
          end if;
        if(cVar1S31S42P068N015P059P032(0)='1' AND  E( 2)='0' AND E(11)='1' )then
          cVar2S31S42P060P057nsss(0) <='1';
          else
          cVar2S31S42P060P057nsss(0) <='0';
          end if;
        if(cVar1S32S42P068N015P059P032(0)='1' AND  E( 2)='0' AND E(11)='0' AND A(11)='1' )then
          cVar2S32S42P060N057P016nsss(0) <='1';
          else
          cVar2S32S42P060N057P016nsss(0) <='0';
          end if;
        if(cVar1S33S42P068N015P059P032(0)='1' AND  E( 2)='1' AND A( 1)='1' )then
          cVar2S33S42P060P017nsss(0) <='1';
          else
          cVar2S33S42P060P017nsss(0) <='0';
          end if;
        if(cVar1S34S42P068N015P059P032(0)='1' AND  E( 2)='1' AND A( 1)='0' AND A(13)='1' )then
          cVar2S34S42P060N017P012nsss(0) <='1';
          else
          cVar2S34S42P060N017P012nsss(0) <='0';
          end if;
        if(cVar1S35S42P068N015P059N032(0)='1' AND  D( 1)='1' AND B( 9)='0' AND E( 1)='1' )then
          cVar2S35S42P062P036P064nsss(0) <='1';
          else
          cVar2S35S42P062P036P064nsss(0) <='0';
          end if;
        if(cVar1S36S42P068N015P059N032(0)='1' AND  D( 1)='0' AND E( 8)='1' AND A(12)='1' )then
          cVar2S36S42N062P069P014nsss(0) <='1';
          else
          cVar2S36S42N062P069P014nsss(0) <='0';
          end if;
        if(cVar1S0S43P068P069P000P047(0)='1' AND  D(14)='1' AND A( 0)='0' AND A( 3)='0' )then
          cVar2S0S43P043P019P013nsss(0) <='1';
          else
          cVar2S0S43P043P019P013nsss(0) <='0';
          end if;
        if(cVar1S1S43P068P069P000P047(0)='1' AND  D(14)='1' AND A( 0)='1' AND A(17)='0' )then
          cVar2S1S43P043P019P004nsss(0) <='1';
          else
          cVar2S1S43P043P019P004nsss(0) <='0';
          end if;
        if(cVar1S2S43P068P069P000P047(0)='1' AND  D(14)='0' AND B(15)='0' )then
          cVar2S2S43N043P024nsss(0) <='1';
          else
          cVar2S2S43N043P024nsss(0) <='0';
          end if;
        if(cVar1S3S43P068P069P000P047(0)='1' AND  D(14)='0' AND B(15)='1' AND E( 3)='1' )then
          cVar2S3S43N043P024P056nsss(0) <='1';
          else
          cVar2S3S43N043P024P056nsss(0) <='0';
          end if;
        if(cVar1S4S43P068P069P000P047(0)='1' AND  B(15)='1' AND E(13)='0' )then
          cVar2S4S43P024P049nsss(0) <='1';
          else
          cVar2S4S43P024P049nsss(0) <='0';
          end if;
        if(cVar1S5S43P068P069P000P047(0)='1' AND  B(15)='1' AND E(13)='1' AND A(16)='1' )then
          cVar2S5S43P024P049P006nsss(0) <='1';
          else
          cVar2S5S43P024P049P006nsss(0) <='0';
          end if;
        if(cVar1S6S43P068P069P000P047(0)='1' AND  B(15)='0' AND E( 1)='0' AND A( 3)='1' )then
          cVar2S6S43N024P064P013nsss(0) <='1';
          else
          cVar2S6S43N024P064P013nsss(0) <='0';
          end if;
        if(cVar1S7S43P068P069P000P064(0)='1' AND  B( 0)='1' )then
          cVar2S7S43P037nsss(0) <='1';
          else
          cVar2S7S43P037nsss(0) <='0';
          end if;
        if(cVar1S8S43P068P069P000N064(0)='1' AND  A(10)='1' AND A(13)='1' )then
          cVar2S8S43P018P012nsss(0) <='1';
          else
          cVar2S8S43P018P012nsss(0) <='0';
          end if;
        if(cVar1S9S43P068P069P000N064(0)='1' AND  A(10)='0' AND A( 1)='0' AND A(14)='0' )then
          cVar2S9S43N018P017P010nsss(0) <='1';
          else
          cVar2S9S43N018P017P010nsss(0) <='0';
          end if;
        if(cVar1S10S43P068P069P023P019(0)='1' AND  B(16)='0' AND A( 2)='0' AND B( 4)='0' )then
          cVar2S10S43P022P015P029nsss(0) <='1';
          else
          cVar2S10S43P022P015P029nsss(0) <='0';
          end if;
        if(cVar1S11S43P068P069P023P019(0)='1' AND  B(16)='0' AND A( 2)='1' AND A( 5)='1' )then
          cVar2S11S43P022P015P009nsss(0) <='1';
          else
          cVar2S11S43P022P015P009nsss(0) <='0';
          end if;
        if(cVar1S12S43P068P069P023P019(0)='1' AND  E( 1)='1' AND A( 1)='0' )then
          cVar2S12S43P064P017nsss(0) <='1';
          else
          cVar2S12S43P064P017nsss(0) <='0';
          end if;
        if(cVar1S13S43P068P069P023P019(0)='1' AND  E( 1)='1' AND A( 1)='1' AND A(11)='1' )then
          cVar2S13S43P064P017P016nsss(0) <='1';
          else
          cVar2S13S43P064P017P016nsss(0) <='0';
          end if;
        if(cVar1S14S43P068P069P023P019(0)='1' AND  E( 1)='0' AND D( 0)='0' AND A(13)='0' )then
          cVar2S14S43N064P066P012nsss(0) <='1';
          else
          cVar2S14S43N064P066P012nsss(0) <='0';
          end if;
        if(cVar1S16S43N068P004P025N048(0)='1' AND  A(13)='0' )then
          cVar2S16S43P012nsss(0) <='1';
          else
          cVar2S16S43P012nsss(0) <='0';
          end if;
        if(cVar1S17S43N068P004N025P040(0)='1' AND  A( 0)='1' )then
          cVar2S17S43P019nsss(0) <='1';
          else
          cVar2S17S43P019nsss(0) <='0';
          end if;
        if(cVar1S18S43N068P004N025P040(0)='1' AND  A( 0)='0' AND B( 8)='1' )then
          cVar2S18S43N019P021nsss(0) <='1';
          else
          cVar2S18S43N019P021nsss(0) <='0';
          end if;
        if(cVar1S19S43N068P004N025P040(0)='1' AND  A( 0)='0' AND B( 8)='0' AND B(17)='1' )then
          cVar2S19S43N019N021P020nsss(0) <='1';
          else
          cVar2S19S43N019N021P020nsss(0) <='0';
          end if;
        if(cVar1S20S43N068P004N025N040(0)='1' AND  D( 6)='1' AND A( 1)='1' )then
          cVar2S20S43P042P017nsss(0) <='1';
          else
          cVar2S20S43P042P017nsss(0) <='0';
          end if;
        if(cVar1S21S43N068P004N025N040(0)='1' AND  D( 6)='1' AND A( 1)='0' AND B( 9)='0' )then
          cVar2S21S43P042N017P036nsss(0) <='1';
          else
          cVar2S21S43P042N017P036nsss(0) <='0';
          end if;
        if(cVar1S22S43N068P004N025N040(0)='1' AND  D( 6)='0' AND B( 8)='0' AND A(10)='0' )then
          cVar2S22S43N042P021P018nsss(0) <='1';
          else
          cVar2S22S43N042P021P018nsss(0) <='0';
          end if;
        if(cVar1S23S43N068N004P013P064(0)='1' AND  B( 7)='0' AND E(11)='1' )then
          cVar2S23S43P023P057nsss(0) <='1';
          else
          cVar2S23S43P023P057nsss(0) <='0';
          end if;
        if(cVar1S24S43N068N004P013P064(0)='1' AND  B( 7)='0' AND E(11)='0' AND B( 9)='1' )then
          cVar2S24S43P023N057P036nsss(0) <='1';
          else
          cVar2S24S43P023N057P036nsss(0) <='0';
          end if;
        if(cVar1S25S43N068N004P013N064(0)='1' AND  D( 0)='0' AND E( 4)='1' AND E( 9)='0' )then
          cVar2S25S43P066P052P065nsss(0) <='1';
          else
          cVar2S25S43P066P052P065nsss(0) <='0';
          end if;
        if(cVar1S26S43N068N004P013N064(0)='1' AND  D( 0)='0' AND E( 4)='0' AND D( 2)='1' )then
          cVar2S26S43P066N052P058nsss(0) <='1';
          else
          cVar2S26S43P066N052P058nsss(0) <='0';
          end if;
        if(cVar1S27S43N068N004P013N064(0)='1' AND  D( 0)='1' AND D( 8)='1' AND A( 2)='1' )then
          cVar2S27S43P066P067P015nsss(0) <='1';
          else
          cVar2S27S43P066P067P015nsss(0) <='0';
          end if;
        if(cVar1S28S43N068N004N013P032(0)='1' AND  E( 4)='0' AND B( 1)='0' AND A( 1)='1' )then
          cVar2S28S43P052P035P017nsss(0) <='1';
          else
          cVar2S28S43P052P035P017nsss(0) <='0';
          end if;
        if(cVar1S29S43N068N004N013P032(0)='1' AND  E( 4)='0' AND B( 1)='1' AND A(11)='1' )then
          cVar2S29S43P052P035P016nsss(0) <='1';
          else
          cVar2S29S43P052P035P016nsss(0) <='0';
          end if;
        if(cVar1S30S43N068N004N013P032(0)='1' AND  E( 4)='1' AND A(14)='1' )then
          cVar2S30S43P052P010nsss(0) <='1';
          else
          cVar2S30S43P052P010nsss(0) <='0';
          end if;
        if(cVar1S31S43N068N004N013P032(0)='1' AND  E( 4)='1' AND A(14)='0' AND D(10)='0' )then
          cVar2S31S43P052N010P059nsss(0) <='1';
          else
          cVar2S31S43P052N010P059nsss(0) <='0';
          end if;
        if(cVar1S32S43N068N004N013N032(0)='1' AND  B(15)='1' AND A( 6)='1' )then
          cVar2S32S43P024P007nsss(0) <='1';
          else
          cVar2S32S43P024P007nsss(0) <='0';
          end if;
        if(cVar1S33S43N068N004N013N032(0)='1' AND  B(15)='1' AND A( 6)='0' AND A(16)='1' )then
          cVar2S33S43P024N007P006nsss(0) <='1';
          else
          cVar2S33S43P024N007P006nsss(0) <='0';
          end if;
        if(cVar1S0S44P068P001P018P065(0)='1' AND  B(14)='0' AND B( 4)='0' AND E( 2)='0' )then
          cVar2S0S44P026P029P060nsss(0) <='1';
          else
          cVar2S0S44P026P029P060nsss(0) <='0';
          end if;
        if(cVar1S1S44P068P001P018N065(0)='1' AND  D( 3)='0' AND B( 1)='0' AND E( 8)='1' )then
          cVar2S1S44P054P035P069nsss(0) <='1';
          else
          cVar2S1S44P054P035P069nsss(0) <='0';
          end if;
        if(cVar1S2S44P068P001P018N065(0)='1' AND  D( 3)='0' AND B( 1)='1' AND E(13)='1' )then
          cVar2S2S44P054P035P049nsss(0) <='1';
          else
          cVar2S2S44P054P035P049nsss(0) <='0';
          end if;
        if(cVar1S3S44P068P001P018N065(0)='1' AND  D( 3)='1' AND A(13)='1' AND B( 0)='0' )then
          cVar2S3S44P054P012P037nsss(0) <='1';
          else
          cVar2S3S44P054P012P037nsss(0) <='0';
          end if;
        if(cVar1S4S44P068P001P018N065(0)='1' AND  D( 3)='1' AND A(13)='0' AND A(14)='1' )then
          cVar2S4S44P054N012P010nsss(0) <='1';
          else
          cVar2S4S44P054N012P010nsss(0) <='0';
          end if;
        if(cVar1S5S44P068P001N018P046(0)='1' AND  D( 6)='0' AND D(13)='0' AND E( 9)='0' )then
          cVar2S5S44P042P047P065nsss(0) <='1';
          else
          cVar2S5S44P042P047P065nsss(0) <='0';
          end if;
        if(cVar1S6S44P068P001N018P046(0)='1' AND  D( 6)='0' AND D(13)='1' AND A( 1)='1' )then
          cVar2S6S44P042P047P017nsss(0) <='1';
          else
          cVar2S6S44P042P047P017nsss(0) <='0';
          end if;
        if(cVar1S7S44P068P001N018N046(0)='1' AND  D( 7)='1' AND A(18)='1' )then
          cVar2S7S44P038P002nsss(0) <='1';
          else
          cVar2S7S44P038P002nsss(0) <='0';
          end if;
        if(cVar1S8S44P068P001N018N046(0)='1' AND  D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar2S8S44P038N002P004nsss(0) <='1';
          else
          cVar2S8S44P038N002P004nsss(0) <='0';
          end if;
        if(cVar1S9S44P068P001N018N046(0)='1' AND  D( 7)='0' AND E( 6)='1' )then
          cVar2S9S44N038P044nsss(0) <='1';
          else
          cVar2S9S44N038P044nsss(0) <='0';
          end if;
        if(cVar1S10S44P068P001N018N046(0)='1' AND  D( 7)='0' AND E( 6)='0' AND A(12)='1' )then
          cVar2S10S44N038N044P014nsss(0) <='1';
          else
          cVar2S10S44N038N044P014nsss(0) <='0';
          end if;
        if(cVar1S11S44P068P001P054P036(0)='1' AND  B( 2)='0' AND A(12)='1' AND A( 2)='0' )then
          cVar2S11S44P033P014P015nsss(0) <='1';
          else
          cVar2S11S44P033P014P015nsss(0) <='0';
          end if;
        if(cVar1S12S44P068P001P054P036(0)='1' AND  B( 2)='0' AND A(12)='0' AND E( 7)='1' )then
          cVar2S12S44P033N014P040nsss(0) <='1';
          else
          cVar2S12S44P033N014P040nsss(0) <='0';
          end if;
        if(cVar1S13S44P068P001P054P036(0)='1' AND  B( 2)='1' AND A( 5)='0' AND A( 1)='1' )then
          cVar2S13S44P033P009P017nsss(0) <='1';
          else
          cVar2S13S44P033P009P017nsss(0) <='0';
          end if;
        if(cVar1S14S44P068P001P054P036(0)='1' AND  D( 8)='1' AND A(10)='1' )then
          cVar2S14S44P067P018nsss(0) <='1';
          else
          cVar2S14S44P067P018nsss(0) <='0';
          end if;
        if(cVar1S15S44P068P067P057P023(0)='1' AND  D( 7)='0' )then
          cVar2S15S44P038nsss(0) <='1';
          else
          cVar2S15S44P038nsss(0) <='0';
          end if;
        if(cVar1S17S44P068P067P057N032(0)='1' AND  B( 1)='1' )then
          cVar2S17S44P035nsss(0) <='1';
          else
          cVar2S17S44P035nsss(0) <='0';
          end if;
        if(cVar1S18S44P068P067P057N032(0)='1' AND  B( 1)='0' AND B( 0)='1' AND B(12)='1' )then
          cVar2S18S44N035P037P030nsss(0) <='1';
          else
          cVar2S18S44N035P037P030nsss(0) <='0';
          end if;
        if(cVar1S19S44P068N067P025P016(0)='1' AND  B( 0)='1' )then
          cVar2S19S44P037nsss(0) <='1';
          else
          cVar2S19S44P037nsss(0) <='0';
          end if;
        if(cVar1S20S44P068N067P025P016(0)='1' AND  B( 0)='0' AND A( 1)='1' )then
          cVar2S20S44N037P017nsss(0) <='1';
          else
          cVar2S20S44N037P017nsss(0) <='0';
          end if;
        if(cVar1S21S44P068N067P025P016(0)='1' AND  B( 0)='0' AND A( 1)='0' AND A( 3)='0' )then
          cVar2S21S44N037N017P013nsss(0) <='1';
          else
          cVar2S21S44N037N017P013nsss(0) <='0';
          end if;
        if(cVar1S22S44P068N067P025P016(0)='1' AND  A( 2)='0' AND A(10)='0' )then
          cVar2S22S44P015P018nsss(0) <='1';
          else
          cVar2S22S44P015P018nsss(0) <='0';
          end if;
        if(cVar1S23S44P068N067N025P066(0)='1' AND  A( 2)='1' AND D(10)='1' AND B(11)='0' )then
          cVar2S23S44P015P059P032nsss(0) <='1';
          else
          cVar2S23S44P015P059P032nsss(0) <='0';
          end if;
        if(cVar1S24S44P068N067N025N066(0)='1' AND  A( 8)='1' AND A(13)='0' AND A(11)='1' )then
          cVar2S24S44P003P012P016nsss(0) <='1';
          else
          cVar2S24S44P003P012P016nsss(0) <='0';
          end if;
        if(cVar1S25S44P068N067N025N066(0)='1' AND  A( 8)='1' AND A(13)='1' AND A(12)='1' )then
          cVar2S25S44P003P012P014nsss(0) <='1';
          else
          cVar2S25S44P003P012P014nsss(0) <='0';
          end if;
        if(cVar1S0S45P014P068P016P067(0)='1' AND  D( 1)='0' AND D( 0)='1' AND E( 1)='1' )then
          cVar2S0S45P062P066P064nsss(0) <='1';
          else
          cVar2S0S45P062P066P064nsss(0) <='0';
          end if;
        if(cVar1S1S45P014P068P016P067(0)='1' AND  D( 1)='0' AND D( 0)='0' AND E( 1)='0' )then
          cVar2S1S45P062N066P064nsss(0) <='1';
          else
          cVar2S1S45P062N066P064nsss(0) <='0';
          end if;
        if(cVar1S2S45P014P068P016P067(0)='1' AND  D( 1)='1' )then
          cVar2S2S45P062psss(0) <='1';
          else
          cVar2S2S45P062psss(0) <='0';
          end if;
        if(cVar1S3S45P014P068P016P067(0)='1' AND  B(15)='1' )then
          cVar2S3S45P024nsss(0) <='1';
          else
          cVar2S3S45P024nsss(0) <='0';
          end if;
        if(cVar1S4S45P014P068P016P067(0)='1' AND  B(15)='0' AND D( 0)='0' AND D( 6)='0' )then
          cVar2S4S45N024P066P042nsss(0) <='1';
          else
          cVar2S4S45N024P066P042nsss(0) <='0';
          end if;
        if(cVar1S5S45P014P068N016P036(0)='1' AND  A( 0)='1' AND B(10)='0' AND D( 3)='0' )then
          cVar2S5S45P019P034P054nsss(0) <='1';
          else
          cVar2S5S45P019P034P054nsss(0) <='0';
          end if;
        if(cVar1S6S45P014P068N016P036(0)='1' AND  A( 0)='1' AND B(10)='1' AND E( 2)='1' )then
          cVar2S6S45P019P034P060nsss(0) <='1';
          else
          cVar2S6S45P019P034P060nsss(0) <='0';
          end if;
        if(cVar1S7S45P014P068N016P036(0)='1' AND  A( 0)='0' AND B( 4)='1' AND D(10)='0' )then
          cVar2S7S45N019P029P059nsss(0) <='1';
          else
          cVar2S7S45N019P029P059nsss(0) <='0';
          end if;
        if(cVar1S8S45P014P068N016P036(0)='1' AND  A( 0)='0' AND B( 4)='0' AND A(13)='1' )then
          cVar2S8S45N019N029P012nsss(0) <='1';
          else
          cVar2S8S45N019N029P012nsss(0) <='0';
          end if;
        if(cVar1S9S45P014P068N016P036(0)='1' AND  A( 1)='1' AND E(14)='0' AND E( 2)='0' )then
          cVar2S9S45P017P045P060nsss(0) <='1';
          else
          cVar2S9S45P017P045P060nsss(0) <='0';
          end if;
        if(cVar1S10S45P014P068N016P036(0)='1' AND  A( 1)='0' AND A( 0)='1' AND B(10)='0' )then
          cVar2S10S45N017P019P034nsss(0) <='1';
          else
          cVar2S10S45N017P019P034nsss(0) <='0';
          end if;
        if(cVar1S11S45P014P068N016P036(0)='1' AND  A( 1)='0' AND A( 0)='0' AND E( 2)='1' )then
          cVar2S11S45N017N019P060nsss(0) <='1';
          else
          cVar2S11S45N017N019P060nsss(0) <='0';
          end if;
        if(cVar1S12S45P014P068P067P045(0)='1' AND  A(15)='1' )then
          cVar2S12S45P008nsss(0) <='1';
          else
          cVar2S12S45P008nsss(0) <='0';
          end if;
        if(cVar1S13S45P014P068P067P045(0)='1' AND  A(15)='0' AND B( 9)='0' )then
          cVar2S13S45N008P036nsss(0) <='1';
          else
          cVar2S13S45N008P036nsss(0) <='0';
          end if;
        if(cVar1S14S45P014P068P067N045(0)='1' AND  B( 5)='1' AND E( 9)='0' )then
          cVar2S14S45P027P065nsss(0) <='1';
          else
          cVar2S14S45P027P065nsss(0) <='0';
          end if;
        if(cVar1S15S45P014P068P067N045(0)='1' AND  B( 5)='0' AND A( 5)='0' AND A(14)='0' )then
          cVar2S15S45N027P009P010nsss(0) <='1';
          else
          cVar2S15S45N027P009P010nsss(0) <='0';
          end if;
        if(cVar1S16S45P014P068P067N045(0)='1' AND  B( 5)='0' AND A( 5)='1' AND A(17)='1' )then
          cVar2S16S45N027P009P004nsss(0) <='1';
          else
          cVar2S16S45N027P009P004nsss(0) <='0';
          end if;
        if(cVar1S17S45P014P068P067P035(0)='1' AND  D( 1)='1' )then
          cVar2S17S45P062nsss(0) <='1';
          else
          cVar2S17S45P062nsss(0) <='0';
          end if;
        if(cVar1S18S45P014P068P067P035(0)='1' AND  D( 1)='0' AND A( 2)='0' AND A(11)='1' )then
          cVar2S18S45N062P015P016nsss(0) <='1';
          else
          cVar2S18S45N062P015P016nsss(0) <='0';
          end if;
        if(cVar1S19S45P014P015P021P034(0)='1' AND  A(15)='0' )then
          cVar2S19S45P008nsss(0) <='1';
          else
          cVar2S19S45P008nsss(0) <='0';
          end if;
        if(cVar1S20S45P014P015P021P034(0)='1' AND  A(15)='1' AND E( 9)='0' AND B( 1)='1' )then
          cVar2S20S45P008P065P035nsss(0) <='1';
          else
          cVar2S20S45P008P065P035nsss(0) <='0';
          end if;
        if(cVar1S21S45P014P015P021N034(0)='1' AND  A(14)='1' AND E( 2)='1' )then
          cVar2S21S45P010P060nsss(0) <='1';
          else
          cVar2S21S45P010P060nsss(0) <='0';
          end if;
        if(cVar1S22S45P014P015P021N034(0)='1' AND  A(14)='1' AND E( 2)='0' AND B( 4)='1' )then
          cVar2S22S45P010N060P029nsss(0) <='1';
          else
          cVar2S22S45P010N060P029nsss(0) <='0';
          end if;
        if(cVar1S23S45P014P015P021N034(0)='1' AND  A(14)='0' AND A( 7)='1' AND E(12)='0' )then
          cVar2S23S45N010P005P053nsss(0) <='1';
          else
          cVar2S23S45N010P005P053nsss(0) <='0';
          end if;
        if(cVar1S24S45P014P015P021P037(0)='1' AND  A( 1)='0' )then
          cVar2S24S45P017nsss(0) <='1';
          else
          cVar2S24S45P017nsss(0) <='0';
          end if;
        if(cVar1S25S45P014P015P021N037(0)='1' AND  A(14)='0' AND A(13)='0' AND B(11)='1' )then
          cVar2S25S45P010P012P032nsss(0) <='1';
          else
          cVar2S25S45P010P012P032nsss(0) <='0';
          end if;
        if(cVar1S26S45P014P015P018P061(0)='1' AND  D( 0)='1' )then
          cVar2S26S45P066nsss(0) <='1';
          else
          cVar2S26S45P066nsss(0) <='0';
          end if;
        if(cVar1S27S45P014P015P018P061(0)='1' AND  D( 0)='0' AND A(11)='0' AND B(10)='0' )then
          cVar2S27S45N066P016P034nsss(0) <='1';
          else
          cVar2S27S45N066P016P034nsss(0) <='0';
          end if;
        if(cVar1S28S45P014P015P018N061(0)='1' AND  E( 9)='1' AND D(10)='0' AND A( 3)='0' )then
          cVar2S28S45P065P059P013nsss(0) <='1';
          else
          cVar2S28S45P065P059P013nsss(0) <='0';
          end if;
        if(cVar1S29S45P014P015P018N061(0)='1' AND  E( 9)='0' AND D( 5)='0' AND D( 1)='1' )then
          cVar2S29S45N065P046P062nsss(0) <='1';
          else
          cVar2S29S45N065P046P062nsss(0) <='0';
          end if;
        if(cVar1S30S45P014P015N018P034(0)='1' AND  E(12)='1' )then
          cVar2S30S45P053nsss(0) <='1';
          else
          cVar2S30S45P053nsss(0) <='0';
          end if;
        if(cVar1S1S46P016P038N021P019(0)='1' AND  D( 2)='1' )then
          cVar2S1S46P058nsss(0) <='1';
          else
          cVar2S1S46P058nsss(0) <='0';
          end if;
        if(cVar1S2S46P016P038N021P019(0)='1' AND  D( 2)='0' AND A( 6)='1' )then
          cVar2S2S46N058P007nsss(0) <='1';
          else
          cVar2S2S46N058P007nsss(0) <='0';
          end if;
        if(cVar1S3S46P016P038N021P019(0)='1' AND  D( 2)='0' AND A( 6)='0' AND E( 9)='1' )then
          cVar2S3S46N058N007P065nsss(0) <='1';
          else
          cVar2S3S46N058N007P065nsss(0) <='0';
          end if;
        if(cVar1S4S46P016P038N021P019(0)='1' AND  E( 8)='0' AND B( 0)='0' AND A(12)='1' )then
          cVar2S4S46N069N037P014nsss(0) <='1';
          else
          cVar2S4S46N069N037P014nsss(0) <='0';
          end if;
        if(cVar1S5S46P016N038P010P036(0)='1' AND  B(10)='0' AND A( 4)='0' )then
          cVar2S5S46P034P011nsss(0) <='1';
          else
          cVar2S5S46P034P011nsss(0) <='0';
          end if;
        if(cVar1S6S46P016N038P010P036(0)='1' AND  B(10)='0' AND A( 4)='1' AND D( 0)='0' )then
          cVar2S6S46P034P011P066nsss(0) <='1';
          else
          cVar2S6S46P034P011P066nsss(0) <='0';
          end if;
        if(cVar1S7S46P016N038P010P036(0)='1' AND  B(10)='1' AND A(12)='0' AND E( 9)='1' )then
          cVar2S7S46P034P014P065nsss(0) <='1';
          else
          cVar2S7S46P034P014P065nsss(0) <='0';
          end if;
        if(cVar1S8S46P016N038P010P036(0)='1' AND  B(10)='1' AND A(12)='1' AND B( 2)='1' )then
          cVar2S8S46P034P014P033nsss(0) <='1';
          else
          cVar2S8S46P034P014P033nsss(0) <='0';
          end if;
        if(cVar1S9S46P016N038P010P036(0)='1' AND  A( 0)='1' AND D( 4)='1' )then
          cVar2S9S46P019P050nsss(0) <='1';
          else
          cVar2S9S46P019P050nsss(0) <='0';
          end if;
        if(cVar1S10S46P016N038P010P036(0)='1' AND  A( 0)='1' AND D( 4)='0' AND A( 2)='0' )then
          cVar2S10S46P019N050P015nsss(0) <='1';
          else
          cVar2S10S46P019N050P015nsss(0) <='0';
          end if;
        if(cVar1S11S46P016N038N010P008(0)='1' AND  D( 5)='1' AND B(10)='0' )then
          cVar2S11S46P046P034nsss(0) <='1';
          else
          cVar2S11S46P046P034nsss(0) <='0';
          end if;
        if(cVar1S12S46P016N038N010P008(0)='1' AND  D( 5)='0' AND A( 1)='1' AND A(18)='0' )then
          cVar2S12S46N046P017P002nsss(0) <='1';
          else
          cVar2S12S46N046P017P002nsss(0) <='0';
          end if;
        if(cVar1S13S46P016N038N010P008(0)='1' AND  D( 5)='0' AND A( 1)='0' AND D( 3)='1' )then
          cVar2S13S46N046N017P054nsss(0) <='1';
          else
          cVar2S13S46N046N017P054nsss(0) <='0';
          end if;
        if(cVar1S14S46P016N038N010N008(0)='1' AND  D( 8)='1' AND B( 4)='0' AND D( 4)='0' )then
          cVar2S14S46P067P029P050nsss(0) <='1';
          else
          cVar2S14S46P067P029P050nsss(0) <='0';
          end if;
        if(cVar1S15S46P016N038N010N008(0)='1' AND  D( 8)='0' AND E( 1)='1' AND E( 0)='0' )then
          cVar2S15S46N067P064P068nsss(0) <='1';
          else
          cVar2S15S46N067P064P068nsss(0) <='0';
          end if;
        if(cVar1S16S46P016N038N010N008(0)='1' AND  D( 8)='0' AND E( 1)='0' AND A(16)='1' )then
          cVar2S16S46N067N064P006nsss(0) <='1';
          else
          cVar2S16S46N067N064P006nsss(0) <='0';
          end if;
        if(cVar1S17S46P016P032P049P056(0)='1' AND  A( 7)='0' AND B( 0)='1' )then
          cVar2S17S46P005P037nsss(0) <='1';
          else
          cVar2S17S46P005P037nsss(0) <='0';
          end if;
        if(cVar1S18S46P016P032P049P056(0)='1' AND  A( 7)='0' AND B( 0)='0' AND A( 2)='0' )then
          cVar2S18S46P005N037P015nsss(0) <='1';
          else
          cVar2S18S46P005N037P015nsss(0) <='0';
          end if;
        if(cVar1S19S46P016P032P049P056(0)='1' AND  A( 4)='0' AND A(12)='1' )then
          cVar2S19S46P011P014nsss(0) <='1';
          else
          cVar2S19S46P011P014nsss(0) <='0';
          end if;
        if(cVar1S20S46P016N032P018P035(0)='1' AND  E( 3)='0' AND B( 0)='0' AND E( 5)='0' )then
          cVar2S20S46P056P037P048nsss(0) <='1';
          else
          cVar2S20S46P056P037P048nsss(0) <='0';
          end if;
        if(cVar1S21S46P016N032P018P035(0)='1' AND  E( 3)='0' AND B( 0)='1' AND E( 1)='1' )then
          cVar2S21S46P056P037P064nsss(0) <='1';
          else
          cVar2S21S46P056P037P064nsss(0) <='0';
          end if;
        if(cVar1S22S46P016N032P018P035(0)='1' AND  E( 3)='1' AND E( 9)='0' AND B( 3)='1' )then
          cVar2S22S46P056P065P031nsss(0) <='1';
          else
          cVar2S22S46P056P065P031nsss(0) <='0';
          end if;
        if(cVar1S23S46P016N032P018P035(0)='1' AND  E( 3)='1' AND E( 9)='1' AND B( 4)='1' )then
          cVar2S23S46P056P065P029nsss(0) <='1';
          else
          cVar2S23S46P056P065P029nsss(0) <='0';
          end if;
        if(cVar1S24S46P016N032P018P035(0)='1' AND  E( 1)='0' AND A(13)='0' )then
          cVar2S24S46P064P012nsss(0) <='1';
          else
          cVar2S24S46P064P012nsss(0) <='0';
          end if;
        if(cVar1S25S46P016N032P018P035(0)='1' AND  E( 1)='1' AND D( 1)='1' AND A( 5)='1' )then
          cVar2S25S46P064P062P009nsss(0) <='1';
          else
          cVar2S25S46P064P062P009nsss(0) <='0';
          end if;
        if(cVar1S26S46P016N032P018P058(0)='1' AND  D( 1)='0' AND A( 2)='0' AND E( 2)='1' )then
          cVar2S26S46P062P015P060nsss(0) <='1';
          else
          cVar2S26S46P062P015P060nsss(0) <='0';
          end if;
        if(cVar1S27S46P016N032P018P058(0)='1' AND  D( 1)='0' AND A( 2)='1' AND B( 1)='0' )then
          cVar2S27S46P062P015P035nsss(0) <='1';
          else
          cVar2S27S46P062P015P035nsss(0) <='0';
          end if;
        if(cVar1S28S46P016N032P018P058(0)='1' AND  D( 1)='1' AND E( 0)='0' AND E( 1)='1' )then
          cVar2S28S46P062P068P064nsss(0) <='1';
          else
          cVar2S28S46P062P068P064nsss(0) <='0';
          end if;
        if(cVar1S29S46P016N032P018N058(0)='1' AND  A( 2)='1' AND D( 0)='0' AND B( 4)='0' )then
          cVar2S29S46P015P066P029nsss(0) <='1';
          else
          cVar2S29S46P015P066P029nsss(0) <='0';
          end if;
        if(cVar1S30S46P016N032P018N058(0)='1' AND  A( 2)='1' AND D( 0)='1' AND D( 9)='0' )then
          cVar2S30S46P015P066P063nsss(0) <='1';
          else
          cVar2S30S46P015P066P063nsss(0) <='0';
          end if;
        if(cVar1S31S46P016N032P018N058(0)='1' AND  A( 2)='0' AND A( 0)='1' AND D( 1)='1' )then
          cVar2S31S46N015P019P062nsss(0) <='1';
          else
          cVar2S31S46N015P019P062nsss(0) <='0';
          end if;
        if(cVar1S32S46P016N032P018N058(0)='1' AND  A( 2)='0' AND A( 0)='0' AND A( 5)='1' )then
          cVar2S32S46N015N019P009nsss(0) <='1';
          else
          cVar2S32S46N015N019P009nsss(0) <='0';
          end if;
        if(cVar1S0S47P067P016P064P047(0)='1' AND  E( 5)='0' AND B( 3)='0' )then
          cVar2S0S47P048P031nsss(0) <='1';
          else
          cVar2S0S47P048P031nsss(0) <='0';
          end if;
        if(cVar1S1S47P067P016P064P047(0)='1' AND  E( 5)='1' AND A(10)='1' )then
          cVar2S1S47P048P018nsss(0) <='1';
          else
          cVar2S1S47P048P018nsss(0) <='0';
          end if;
        if(cVar1S2S47P067P016P064P047(0)='1' AND  E( 5)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar2S2S47P048N018P019nsss(0) <='1';
          else
          cVar2S2S47P048N018P019nsss(0) <='0';
          end if;
        if(cVar1S3S47P067P016P064N047(0)='1' AND  B( 5)='1' AND E( 5)='1' AND B(10)='0' )then
          cVar2S3S47P027P048P034nsss(0) <='1';
          else
          cVar2S3S47P027P048P034nsss(0) <='0';
          end if;
        if(cVar1S4S47P067P016P064N047(0)='1' AND  B( 5)='1' AND E( 5)='0' AND E( 0)='1' )then
          cVar2S4S47P027N048P068nsss(0) <='1';
          else
          cVar2S4S47P027N048P068nsss(0) <='0';
          end if;
        if(cVar1S5S47P067P016P064N047(0)='1' AND  B( 5)='0' AND D(12)='1' )then
          cVar2S5S47N027P051nsss(0) <='1';
          else
          cVar2S5S47N027P051nsss(0) <='0';
          end if;
        if(cVar1S6S47P067P016P064N047(0)='1' AND  B( 5)='0' AND D(12)='0' AND B(14)='0' )then
          cVar2S6S47N027N051P026nsss(0) <='1';
          else
          cVar2S6S47N027N051P026nsss(0) <='0';
          end if;
        if(cVar1S7S47P067P016P064P048(0)='1' AND  D(13)='0' AND A( 3)='1' AND E( 3)='0' )then
          cVar2S7S47P047P013P056nsss(0) <='1';
          else
          cVar2S7S47P047P013P056nsss(0) <='0';
          end if;
        if(cVar1S8S47P067P016P064P048(0)='1' AND  D(13)='0' AND A( 3)='0' AND D(11)='0' )then
          cVar2S8S47P047N013P055nsss(0) <='1';
          else
          cVar2S8S47P047N013P055nsss(0) <='0';
          end if;
        if(cVar1S9S47P067P016P064P048(0)='1' AND  D(13)='1' AND B( 1)='0' AND D( 0)='0' )then
          cVar2S9S47P047P035P066nsss(0) <='1';
          else
          cVar2S9S47P047P035P066nsss(0) <='0';
          end if;
        if(cVar1S10S47P067P016P064P048(0)='1' AND  D( 5)='1' AND B( 6)='1' )then
          cVar2S10S47P046P025nsss(0) <='1';
          else
          cVar2S10S47P046P025nsss(0) <='0';
          end if;
        if(cVar1S11S47P067P016P064P048(0)='1' AND  D( 5)='1' AND B( 6)='0' AND A( 1)='1' )then
          cVar2S11S47P046N025P017nsss(0) <='1';
          else
          cVar2S11S47P046N025P017nsss(0) <='0';
          end if;
        if(cVar1S12S47P067P016P002P006(0)='1' AND  A( 9)='0' AND B( 9)='1' )then
          cVar2S12S47P001P036nsss(0) <='1';
          else
          cVar2S12S47P001P036nsss(0) <='0';
          end if;
        if(cVar1S13S47P067P016P002P006(0)='1' AND  A( 9)='0' AND B( 9)='0' AND B(11)='1' )then
          cVar2S13S47P001N036P032nsss(0) <='1';
          else
          cVar2S13S47P001N036P032nsss(0) <='0';
          end if;
        if(cVar1S14S47P067P016P002P006(0)='1' AND  E( 9)='1' AND A(12)='1' )then
          cVar2S14S47P065P014nsss(0) <='1';
          else
          cVar2S14S47P065P014nsss(0) <='0';
          end if;
        if(cVar1S15S47P067P016P002P006(0)='1' AND  E( 9)='1' AND A(12)='0' AND B( 9)='0' )then
          cVar2S15S47P065N014P036nsss(0) <='1';
          else
          cVar2S15S47P065N014P036nsss(0) <='0';
          end if;
        if(cVar1S16S47P067P016P002P006(0)='1' AND  E( 9)='0' AND B( 1)='1' AND A(12)='0' )then
          cVar2S16S47N065P035P014nsss(0) <='1';
          else
          cVar2S16S47N065P035P014nsss(0) <='0';
          end if;
        if(cVar1S17S47P067P016P002P050(0)='1' AND  D(11)='1' )then
          cVar2S17S47P055nsss(0) <='1';
          else
          cVar2S17S47P055nsss(0) <='0';
          end if;
        if(cVar1S18S47P067P016P002P050(0)='1' AND  D(11)='0' AND A(14)='1' AND A( 3)='0' )then
          cVar2S18S47N055P010P013nsss(0) <='1';
          else
          cVar2S18S47N055P010P013nsss(0) <='0';
          end if;
        if(cVar1S19S47P067P062P058P033(0)='1' AND  A(10)='0' AND B( 9)='1' )then
          cVar2S19S47P018P036nsss(0) <='1';
          else
          cVar2S19S47P018P036nsss(0) <='0';
          end if;
        if(cVar1S20S47P067P062P058P033(0)='1' AND  A(10)='0' AND B( 9)='0' AND A( 2)='1' )then
          cVar2S20S47P018N036P015nsss(0) <='1';
          else
          cVar2S20S47P018N036P015nsss(0) <='0';
          end if;
        if(cVar1S21S47P067P062P058P033(0)='1' AND  A(10)='1' AND A( 0)='0' )then
          cVar2S21S47P018P019nsss(0) <='1';
          else
          cVar2S21S47P018P019nsss(0) <='0';
          end if;
        if(cVar1S22S47P067P062P058N033(0)='1' AND  A(10)='1' AND A(13)='1' AND E( 2)='1' )then
          cVar2S22S47P018P012P060nsss(0) <='1';
          else
          cVar2S22S47P018P012P060nsss(0) <='0';
          end if;
        if(cVar1S23S47P067P062P058N033(0)='1' AND  A(10)='1' AND A(13)='0' AND B(11)='1' )then
          cVar2S23S47P018N012P032nsss(0) <='1';
          else
          cVar2S23S47P018N012P032nsss(0) <='0';
          end if;
        if(cVar1S24S47P067P062P058N033(0)='1' AND  A(10)='0' AND A( 3)='1' )then
          cVar2S24S47N018P013nsss(0) <='1';
          else
          cVar2S24S47N018P013nsss(0) <='0';
          end if;
        if(cVar1S25S47P067P062N058P033(0)='1' AND  B(11)='1' AND E(10)='1' )then
          cVar2S25S47P032P061nsss(0) <='1';
          else
          cVar2S25S47P032P061nsss(0) <='0';
          end if;
        if(cVar1S26S47P067P062N058P033(0)='1' AND  B(11)='1' AND E(10)='0' AND D( 0)='1' )then
          cVar2S26S47P032N061P066nsss(0) <='1';
          else
          cVar2S26S47P032N061P066nsss(0) <='0';
          end if;
        if(cVar1S27S47P067P062N058P033(0)='1' AND  B(11)='0' AND D(10)='1' AND B(12)='1' )then
          cVar2S27S47N032P059P030nsss(0) <='1';
          else
          cVar2S27S47N032P059P030nsss(0) <='0';
          end if;
        if(cVar1S28S47P067P062N058P033(0)='1' AND  A(10)='1' AND B(11)='0' AND A(14)='1' )then
          cVar2S28S47P018P032P010nsss(0) <='1';
          else
          cVar2S28S47P018P032P010nsss(0) <='0';
          end if;
        if(cVar1S29S47P067P062N058P033(0)='1' AND  A(10)='0' AND E(10)='1' )then
          cVar2S29S47N018P061nsss(0) <='1';
          else
          cVar2S29S47N018P061nsss(0) <='0';
          end if;
        if(cVar1S30S47P067P062P044P035(0)='1' AND  E( 1)='0' AND B( 0)='0' )then
          cVar2S30S47P064P037nsss(0) <='1';
          else
          cVar2S30S47P064P037nsss(0) <='0';
          end if;
        if(cVar1S31S47P067P062P044P035(0)='1' AND  E( 1)='1' AND A( 0)='0' AND A( 1)='0' )then
          cVar2S31S47P064P019P017nsss(0) <='1';
          else
          cVar2S31S47P064P019P017nsss(0) <='0';
          end if;
        if(cVar1S32S47P067P062P044N035(0)='1' AND  B( 0)='1' AND A(14)='1' )then
          cVar2S32S47P037P010nsss(0) <='1';
          else
          cVar2S32S47P037P010nsss(0) <='0';
          end if;
        if(cVar1S33S47P067P062P044N035(0)='1' AND  B( 0)='0' AND A( 3)='0' AND E( 0)='1' )then
          cVar2S33S47N037P013P068nsss(0) <='1';
          else
          cVar2S33S47N037P013P068nsss(0) <='0';
          end if;
        if(cVar1S0S48P067P062P057P049(0)='1' AND  A(13)='0' AND D( 9)='0' AND A( 6)='0' )then
          cVar2S0S48P012P063P007nsss(0) <='1';
          else
          cVar2S0S48P012P063P007nsss(0) <='0';
          end if;
        if(cVar1S1S48P067P062P057P049(0)='1' AND  A(13)='1' AND A( 0)='0' )then
          cVar2S1S48P012P019nsss(0) <='1';
          else
          cVar2S1S48P012P019nsss(0) <='0';
          end if;
        if(cVar1S2S48P067P062P057N049(0)='1' AND  E( 8)='1' AND E(15)='1' AND B( 9)='1' )then
          cVar2S2S48P069P041P036nsss(0) <='1';
          else
          cVar2S2S48P069P041P036nsss(0) <='0';
          end if;
        if(cVar1S3S48P067P062P057N049(0)='1' AND  E( 8)='1' AND E(15)='0' AND A( 7)='0' )then
          cVar2S3S48P069N041P005nsss(0) <='1';
          else
          cVar2S3S48P069N041P005nsss(0) <='0';
          end if;
        if(cVar1S4S48P067P062P057N049(0)='1' AND  E( 8)='0' AND D( 5)='0' AND A(11)='0' )then
          cVar2S4S48N069P046P016nsss(0) <='1';
          else
          cVar2S4S48N069P046P016nsss(0) <='0';
          end if;
        if(cVar1S5S48P067P062P057P051(0)='1' AND  D( 0)='0' AND D(10)='0' AND D( 9)='0' )then
          cVar2S5S48P066P059P063nsss(0) <='1';
          else
          cVar2S5S48P066P059P063nsss(0) <='0';
          end if;
        if(cVar1S6S48P067P062P057P051(0)='1' AND  D( 0)='0' AND D(10)='1' AND A(12)='1' )then
          cVar2S6S48P066P059P014nsss(0) <='1';
          else
          cVar2S6S48P066P059P014nsss(0) <='0';
          end if;
        if(cVar1S7S48P067P062P057P051(0)='1' AND  D( 0)='1' AND D(10)='1' )then
          cVar2S7S48P066P059nsss(0) <='1';
          else
          cVar2S7S48P066P059nsss(0) <='0';
          end if;
        if(cVar1S8S48P067P062P057P051(0)='1' AND  D( 0)='1' AND D(10)='0' AND A(12)='1' )then
          cVar2S8S48P066N059P014nsss(0) <='1';
          else
          cVar2S8S48P066N059P014nsss(0) <='0';
          end if;
        if(cVar1S9S48P067P062P044P042(0)='1' AND  B(12)='1' AND A( 0)='1' )then
          cVar2S9S48P030P019nsss(0) <='1';
          else
          cVar2S9S48P030P019nsss(0) <='0';
          end if;
        if(cVar1S10S48N067P036P027P050(0)='1' AND  B(12)='1' )then
          cVar2S10S48P030nsss(0) <='1';
          else
          cVar2S10S48P030nsss(0) <='0';
          end if;
        if(cVar1S11S48N067P036P027P050(0)='1' AND  B(12)='0' AND E(12)='0' )then
          cVar2S11S48N030P053nsss(0) <='1';
          else
          cVar2S11S48N030P053nsss(0) <='0';
          end if;
        if(cVar1S12S48N067P036P027P050(0)='1' AND  B(12)='0' AND E(12)='1' AND A( 5)='1' )then
          cVar2S12S48N030P053P009nsss(0) <='1';
          else
          cVar2S12S48N030P053P009nsss(0) <='0';
          end if;
        if(cVar1S13S48N067P036P027N050(0)='1' AND  A(15)='1' AND E( 9)='0' AND E( 5)='1' )then
          cVar2S13S48P008P065P048nsss(0) <='1';
          else
          cVar2S13S48P008P065P048nsss(0) <='0';
          end if;
        if(cVar1S14S48N067P036P027N050(0)='1' AND  A(15)='0' AND D( 0)='1' AND A(10)='1' )then
          cVar2S14S48N008P066P018nsss(0) <='1';
          else
          cVar2S14S48N008P066P018nsss(0) <='0';
          end if;
        if(cVar1S15S48N067P036N027P016(0)='1' AND  A(18)='0' AND A(16)='0' )then
          cVar2S15S48P002P006nsss(0) <='1';
          else
          cVar2S15S48P002P006nsss(0) <='0';
          end if;
        if(cVar1S16S48N067P036N027P016(0)='1' AND  A(18)='0' AND A(16)='1' AND D(12)='1' )then
          cVar2S16S48P002P006P051nsss(0) <='1';
          else
          cVar2S16S48P002P006P051nsss(0) <='0';
          end if;
        if(cVar1S17S48N067P036N027P016(0)='1' AND  A(18)='1' AND B(12)='1' )then
          cVar2S17S48P002P030nsss(0) <='1';
          else
          cVar2S17S48P002P030nsss(0) <='0';
          end if;
        if(cVar1S18S48N067P036N027N016(0)='1' AND  B( 6)='1' AND A( 6)='1' AND D( 6)='0' )then
          cVar2S18S48P025P007P042nsss(0) <='1';
          else
          cVar2S18S48P025P007P042nsss(0) <='0';
          end if;
        if(cVar1S19S48N067P036N027N016(0)='1' AND  B( 6)='1' AND A( 6)='0' AND E(10)='1' )then
          cVar2S19S48P025N007P061nsss(0) <='1';
          else
          cVar2S19S48P025N007P061nsss(0) <='0';
          end if;
        if(cVar1S20S48N067P036N027N016(0)='1' AND  B( 6)='0' AND E( 5)='0' AND B(14)='1' )then
          cVar2S20S48N025P048P026nsss(0) <='1';
          else
          cVar2S20S48N025P048P026nsss(0) <='0';
          end if;
        if(cVar1S21S48N067P036N027N016(0)='1' AND  B( 6)='0' AND E( 5)='1' AND A(16)='1' )then
          cVar2S21S48N025P048P006nsss(0) <='1';
          else
          cVar2S21S48N025P048P006nsss(0) <='0';
          end if;
        if(cVar1S22S48N067P036P005P043(0)='1' AND  A(11)='1' )then
          cVar2S22S48P016nsss(0) <='1';
          else
          cVar2S22S48P016nsss(0) <='0';
          end if;
        if(cVar1S23S48N067P036P005P043(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S23S48N016P018nsss(0) <='1';
          else
          cVar2S23S48N016P018nsss(0) <='0';
          end if;
        if(cVar1S24S48N067P036P005N043(0)='1' AND  E(15)='0' AND B( 2)='1' AND A( 6)='0' )then
          cVar2S24S48P041P033P007nsss(0) <='1';
          else
          cVar2S24S48P041P033P007nsss(0) <='0';
          end if;
        if(cVar1S26S48N067P036P005N032(0)='1' AND  E(10)='1' )then
          cVar2S26S48P061nsss(0) <='1';
          else
          cVar2S26S48P061nsss(0) <='0';
          end if;
        if(cVar1S27S48N067P036P005N032(0)='1' AND  E(10)='0' AND B( 2)='0' AND A(14)='1' )then
          cVar2S27S48N061P033P010nsss(0) <='1';
          else
          cVar2S27S48N061P033P010nsss(0) <='0';
          end if;
        if(cVar1S0S49P036P011P010P013(0)='1' AND  B(13)='1' AND A( 0)='1' )then
          cVar2S0S49P028P019nsss(0) <='1';
          else
          cVar2S0S49P028P019nsss(0) <='0';
          end if;
        if(cVar1S1S49P036P011P010P013(0)='1' AND  B(13)='1' AND A( 0)='0' AND E( 1)='0' )then
          cVar2S1S49P028N019P064nsss(0) <='1';
          else
          cVar2S1S49P028N019P064nsss(0) <='0';
          end if;
        if(cVar1S2S49P036P011P010P013(0)='1' AND  B(13)='0' )then
          cVar2S2S49N028psss(0) <='1';
          else
          cVar2S2S49N028psss(0) <='0';
          end if;
        if(cVar1S3S49P036P011P010P013(0)='1' AND  A( 2)='1' AND B(11)='1' AND D(10)='1' )then
          cVar2S3S49P015P032P059nsss(0) <='1';
          else
          cVar2S3S49P015P032P059nsss(0) <='0';
          end if;
        if(cVar1S4S49P036P011P010P013(0)='1' AND  A( 2)='1' AND B(11)='0' AND E( 0)='1' )then
          cVar2S4S49P015N032P068nsss(0) <='1';
          else
          cVar2S4S49P015N032P068nsss(0) <='0';
          end if;
        if(cVar1S5S49P036P011P010P013(0)='1' AND  A( 2)='0' AND A( 6)='0' AND B( 1)='1' )then
          cVar2S5S49N015P007P035nsss(0) <='1';
          else
          cVar2S5S49N015P007P035nsss(0) <='0';
          end if;
        if(cVar1S7S49P036P011P010N042(0)='1' AND  D( 0)='0' AND A( 7)='0' AND A( 1)='1' )then
          cVar2S7S49P066P005P017nsss(0) <='1';
          else
          cVar2S7S49P066P005P017nsss(0) <='0';
          end if;
        if(cVar1S8S49P036P011P010N042(0)='1' AND  D( 0)='1' AND E( 3)='0' AND E( 8)='1' )then
          cVar2S8S49P066P056P069nsss(0) <='1';
          else
          cVar2S8S49P066P056P069nsss(0) <='0';
          end if;
        if(cVar1S9S49P036N011P005P039(0)='1' AND  B(17)='1' )then
          cVar2S9S49P020nsss(0) <='1';
          else
          cVar2S9S49P020nsss(0) <='0';
          end if;
        if(cVar1S10S49P036N011P005P039(0)='1' AND  B(17)='0' AND A(11)='1' )then
          cVar2S10S49N020P016nsss(0) <='1';
          else
          cVar2S10S49N020P016nsss(0) <='0';
          end if;
        if(cVar1S11S49P036N011P005P039(0)='1' AND  B(17)='0' AND A(11)='0' AND B( 8)='1' )then
          cVar2S11S49N020N016P021nsss(0) <='1';
          else
          cVar2S11S49N020N016P021nsss(0) <='0';
          end if;
        if(cVar1S12S49P036N011P005N039(0)='1' AND  D( 4)='1' AND A( 0)='0' )then
          cVar2S12S49P050P019nsss(0) <='1';
          else
          cVar2S12S49P050P019nsss(0) <='0';
          end if;
        if(cVar1S13S49P036N011P005N039(0)='1' AND  D( 4)='0' AND D(11)='0' AND E(10)='0' )then
          cVar2S13S49N050P055P061nsss(0) <='1';
          else
          cVar2S13S49N050P055P061nsss(0) <='0';
          end if;
        if(cVar1S14S49P036N011N005P016(0)='1' AND  A( 2)='1' AND D( 3)='1' )then
          cVar2S14S49P015P054nsss(0) <='1';
          else
          cVar2S14S49P015P054nsss(0) <='0';
          end if;
        if(cVar1S15S49P036N011N005P016(0)='1' AND  A( 2)='1' AND D( 3)='0' AND A( 3)='0' )then
          cVar2S15S49P015N054P013nsss(0) <='1';
          else
          cVar2S15S49P015N054P013nsss(0) <='0';
          end if;
        if(cVar1S16S49P036N011N005P016(0)='1' AND  A( 2)='0' AND A( 5)='1' AND E( 1)='0' )then
          cVar2S16S49N015P009P064nsss(0) <='1';
          else
          cVar2S16S49N015P009P064nsss(0) <='0';
          end if;
        if(cVar1S17S49P036N011N005P016(0)='1' AND  A( 2)='0' AND A( 5)='0' AND A( 3)='1' )then
          cVar2S17S49N015N009P013nsss(0) <='1';
          else
          cVar2S17S49N015N009P013nsss(0) <='0';
          end if;
        if(cVar1S18S49P036N011N005P016(0)='1' AND  D( 8)='1' AND E( 0)='1' )then
          cVar2S18S49P067P068nsss(0) <='1';
          else
          cVar2S18S49P067P068nsss(0) <='0';
          end if;
        if(cVar1S19S49P036N011N005P016(0)='1' AND  D( 8)='1' AND E( 0)='0' AND E( 3)='1' )then
          cVar2S19S49P067N068P056nsss(0) <='1';
          else
          cVar2S19S49P067N068P056nsss(0) <='0';
          end if;
        if(cVar1S20S49P036N011N005P016(0)='1' AND  D( 8)='0' AND A(18)='1' AND A(17)='1' )then
          cVar2S20S49N067P002P004nsss(0) <='1';
          else
          cVar2S20S49N067P002P004nsss(0) <='0';
          end if;
        if(cVar1S22S49P036P043N022P015(0)='1' AND  A(11)='1' )then
          cVar2S22S49P016nsss(0) <='1';
          else
          cVar2S22S49P016nsss(0) <='0';
          end if;
        if(cVar1S23S49P036P043N022P015(0)='1' AND  A(11)='0' AND A( 0)='1' )then
          cVar2S23S49N016P019nsss(0) <='1';
          else
          cVar2S23S49N016P019nsss(0) <='0';
          end if;
        if(cVar1S24S49P036P043N022P015(0)='1' AND  A(11)='0' AND A( 0)='0' AND E( 8)='0' )then
          cVar2S24S49N016N019P069nsss(0) <='1';
          else
          cVar2S24S49N016N019P069nsss(0) <='0';
          end if;
        if(cVar1S25S49P036N043P045P016(0)='1' AND  E( 9)='0' AND B(16)='0' AND D( 7)='0' )then
          cVar2S25S49P065P022P038nsss(0) <='1';
          else
          cVar2S25S49P065P022P038nsss(0) <='0';
          end if;
        if(cVar1S26S49P036N043P045P016(0)='1' AND  E( 9)='1' AND B(11)='1' AND A( 0)='0' )then
          cVar2S26S49P065P032P019nsss(0) <='1';
          else
          cVar2S26S49P065P032P019nsss(0) <='0';
          end if;
        if(cVar1S27S49P036N043P045N016(0)='1' AND  A(12)='1' AND E( 9)='1' )then
          cVar2S27S49P014P065nsss(0) <='1';
          else
          cVar2S27S49P014P065nsss(0) <='0';
          end if;
        if(cVar1S28S49P036N043P045N016(0)='1' AND  A(12)='1' AND E( 9)='0' AND B( 1)='1' )then
          cVar2S28S49P014N065P035nsss(0) <='1';
          else
          cVar2S28S49P014N065P035nsss(0) <='0';
          end if;
        if(cVar1S29S49P036N043P045N016(0)='1' AND  A(12)='0' AND E( 0)='1' AND B( 2)='0' )then
          cVar2S29S49N014P068P033nsss(0) <='1';
          else
          cVar2S29S49N014P068P033nsss(0) <='0';
          end if;
        if(cVar1S30S49P036N043P045P016(0)='1' AND  B( 0)='1' )then
          cVar2S30S49P037nsss(0) <='1';
          else
          cVar2S30S49P037nsss(0) <='0';
          end if;
        if(cVar1S0S50P036P033P015P038(0)='1' AND  A(18)='1' )then
          cVar2S0S50P002nsss(0) <='1';
          else
          cVar2S0S50P002nsss(0) <='0';
          end if;
        if(cVar1S1S50P036P033P015P038(0)='1' AND  A(18)='0' AND A(17)='1' AND B( 8)='1' )then
          cVar2S1S50N002P004P021nsss(0) <='1';
          else
          cVar2S1S50N002P004P021nsss(0) <='0';
          end if;
        if(cVar1S2S50P036P033P015P038(0)='1' AND  A(18)='0' AND A(17)='0' AND D(15)='0' )then
          cVar2S2S50N002N004P039nsss(0) <='1';
          else
          cVar2S2S50N002N004P039nsss(0) <='0';
          end if;
        if(cVar1S3S50P036P033P015N038(0)='1' AND  B( 7)='1' AND D( 6)='1' AND E( 7)='0' )then
          cVar2S3S50P023P042P040nsss(0) <='1';
          else
          cVar2S3S50P023P042P040nsss(0) <='0';
          end if;
        if(cVar1S4S50P036P033P015N038(0)='1' AND  B( 7)='1' AND D( 6)='0' AND E(14)='1' )then
          cVar2S4S50P023N042P045nsss(0) <='1';
          else
          cVar2S4S50P023N042P045nsss(0) <='0';
          end if;
        if(cVar1S5S50P036P033P015N038(0)='1' AND  B( 7)='0' AND E( 6)='0' )then
          cVar2S5S50N023P044nsss(0) <='1';
          else
          cVar2S5S50N023P044nsss(0) <='0';
          end if;
        if(cVar1S6S50P036P033P015N038(0)='1' AND  B( 7)='0' AND E( 6)='1' AND E(12)='1' )then
          cVar2S6S50N023P044P053nsss(0) <='1';
          else
          cVar2S6S50N023P044P053nsss(0) <='0';
          end if;
        if(cVar1S7S50P036P033P015P049(0)='1' AND  B(13)='1' AND A(14)='1' )then
          cVar2S7S50P028P010nsss(0) <='1';
          else
          cVar2S7S50P028P010nsss(0) <='0';
          end if;
        if(cVar1S8S50P036P033P015P049(0)='1' AND  B(13)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar2S8S50P028N010P011nsss(0) <='1';
          else
          cVar2S8S50P028N010P011nsss(0) <='0';
          end if;
        if(cVar1S9S50P036P033P015P049(0)='1' AND  B(13)='0' AND D( 9)='1' )then
          cVar2S9S50N028P063nsss(0) <='1';
          else
          cVar2S9S50N028P063nsss(0) <='0';
          end if;
        if(cVar1S10S50P036P033P015P049(0)='1' AND  B(13)='0' AND D( 9)='0' AND A( 3)='1' )then
          cVar2S10S50N028N063P013nsss(0) <='1';
          else
          cVar2S10S50N028N063P013nsss(0) <='0';
          end if;
        if(cVar1S11S50P036P033P015P049(0)='1' AND  A( 6)='1' )then
          cVar2S11S50P007nsss(0) <='1';
          else
          cVar2S11S50P007nsss(0) <='0';
          end if;
        if(cVar1S12S50P036P033P015P049(0)='1' AND  A( 6)='0' AND D(13)='1' AND A( 5)='1' )then
          cVar2S12S50N007P047P009nsss(0) <='1';
          else
          cVar2S12S50N007P047P009nsss(0) <='0';
          end if;
        if(cVar1S13S50P036P033P026P001(0)='1' AND  E( 3)='1' AND A(15)='0' AND D(11)='0' )then
          cVar2S13S50P056P008P055nsss(0) <='1';
          else
          cVar2S13S50P056P008P055nsss(0) <='0';
          end if;
        if(cVar1S14S50P036P033P026P001(0)='1' AND  E( 3)='0' AND B( 3)='0' AND A( 8)='0' )then
          cVar2S14S50N056P031P003nsss(0) <='1';
          else
          cVar2S14S50N056P031P003nsss(0) <='0';
          end if;
        if(cVar1S15S50P036P033P026P001(0)='1' AND  E( 3)='0' AND B( 3)='1' AND B(10)='1' )then
          cVar2S15S50N056P031P034nsss(0) <='1';
          else
          cVar2S15S50N056P031P034nsss(0) <='0';
          end if;
        if(cVar1S16S50P036P033P026P001(0)='1' AND  A( 5)='0' AND D( 2)='1' )then
          cVar2S16S50P009P058nsss(0) <='1';
          else
          cVar2S16S50P009P058nsss(0) <='0';
          end if;
        if(cVar1S18S50P036P033P026N047(0)='1' AND  D( 3)='0' AND A(17)='0' AND A(10)='1' )then
          cVar2S18S50P054P004P018nsss(0) <='1';
          else
          cVar2S18S50P054P004P018nsss(0) <='0';
          end if;
        if(cVar1S19S50P036P068P065P018(0)='1' AND  D( 4)='0' AND B(14)='0' AND A(13)='0' )then
          cVar2S19S50P050P026P012nsss(0) <='1';
          else
          cVar2S19S50P050P026P012nsss(0) <='0';
          end if;
        if(cVar1S20S50P036P068P065N018(0)='1' AND  A(13)='1' )then
          cVar2S20S50P012nsss(0) <='1';
          else
          cVar2S20S50P012nsss(0) <='0';
          end if;
        if(cVar1S21S50P036P068P065N018(0)='1' AND  A(13)='0' AND A(11)='1' AND D( 2)='0' )then
          cVar2S21S50N012P016P058nsss(0) <='1';
          else
          cVar2S21S50N012P016P058nsss(0) <='0';
          end if;
        if(cVar1S22S50P036P068P065N018(0)='1' AND  A(13)='0' AND A(11)='0' AND B( 2)='1' )then
          cVar2S22S50N012N016P033nsss(0) <='1';
          else
          cVar2S22S50N012N016P033nsss(0) <='0';
          end if;
        if(cVar1S23S50P036P068N065P018(0)='1' AND  B( 0)='0' AND D( 0)='1' AND D( 8)='0' )then
          cVar2S23S50P037P066P067nsss(0) <='1';
          else
          cVar2S23S50P037P066P067nsss(0) <='0';
          end if;
        if(cVar1S24S50P036P068N065P018(0)='1' AND  B( 0)='0' AND D( 0)='0' AND E( 8)='1' )then
          cVar2S24S50P037N066P069nsss(0) <='1';
          else
          cVar2S24S50P037N066P069nsss(0) <='0';
          end if;
        if(cVar1S25S50P036P068N065P018(0)='1' AND  A(19)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar2S25S50P000P010P069nsss(0) <='1';
          else
          cVar2S25S50P000P010P069nsss(0) <='0';
          end if;
        if(cVar1S26S50P036P068N065P018(0)='1' AND  A(19)='0' AND A(15)='1' AND A( 5)='0' )then
          cVar2S26S50N000P008P009nsss(0) <='1';
          else
          cVar2S26S50N000P008P009nsss(0) <='0';
          end if;
        if(cVar1S28S50P036P068P019N025(0)='1' AND  A( 7)='0' AND D( 3)='1' )then
          cVar2S28S50P005P054nsss(0) <='1';
          else
          cVar2S28S50P005P054nsss(0) <='0';
          end if;
        if(cVar1S29S50P036P068P019N025(0)='1' AND  A( 7)='0' AND D( 3)='0' AND A(10)='1' )then
          cVar2S29S50P005N054P018nsss(0) <='1';
          else
          cVar2S29S50P005N054P018nsss(0) <='0';
          end if;
        if(cVar1S30S50P036P068N019P066(0)='1' AND  B( 0)='1' AND A(10)='1' )then
          cVar2S30S50P037P018nsss(0) <='1';
          else
          cVar2S30S50P037P018nsss(0) <='0';
          end if;
        if(cVar1S31S50P036P068N019P066(0)='1' AND  B( 0)='1' AND A(10)='0' AND A( 1)='0' )then
          cVar2S31S50P037N018P017nsss(0) <='1';
          else
          cVar2S31S50P037N018P017nsss(0) <='0';
          end if;
        if(cVar1S32S50P036P068N019P066(0)='1' AND  B( 0)='0' AND A(13)='0' AND A( 1)='1' )then
          cVar2S32S50N037P012P017nsss(0) <='1';
          else
          cVar2S32S50N037P012P017nsss(0) <='0';
          end if;
        if(cVar1S33S50P036P068N019P066(0)='1' AND  B( 0)='0' AND A(13)='1' AND B( 1)='1' )then
          cVar2S33S50N037P012P035nsss(0) <='1';
          else
          cVar2S33S50N037P012P035nsss(0) <='0';
          end if;
        if(cVar1S34S50P036P068N019N066(0)='1' AND  E( 9)='1' AND E( 8)='1' )then
          cVar2S34S50P065P069nsss(0) <='1';
          else
          cVar2S34S50P065P069nsss(0) <='0';
          end if;
        if(cVar1S0S51P033P015P032P035(0)='1' AND  E( 0)='0' AND D( 4)='0' )then
          cVar2S0S51P068P050nsss(0) <='1';
          else
          cVar2S0S51P068P050nsss(0) <='0';
          end if;
        if(cVar1S1S51P033P015P032P035(0)='1' AND  E( 0)='1' AND E( 2)='1' )then
          cVar2S1S51P068P060nsss(0) <='1';
          else
          cVar2S1S51P068P060nsss(0) <='0';
          end if;
        if(cVar1S2S51P033P015P032P035(0)='1' AND  E(10)='0' AND E( 1)='1' )then
          cVar2S2S51P061P064nsss(0) <='1';
          else
          cVar2S2S51P061P064nsss(0) <='0';
          end if;
        if(cVar1S3S51P033P015P032P035(0)='1' AND  E(10)='0' AND E( 1)='0' AND A(11)='1' )then
          cVar2S3S51P061N064P016nsss(0) <='1';
          else
          cVar2S3S51P061N064P016nsss(0) <='0';
          end if;
        if(cVar1S4S51P033P015P032P035(0)='1' AND  E(10)='1' AND E( 0)='1' )then
          cVar2S4S51P061P068nsss(0) <='1';
          else
          cVar2S4S51P061P068nsss(0) <='0';
          end if;
        if(cVar1S5S51P033P015N032P017(0)='1' AND  A(12)='0' )then
          cVar2S5S51P014nsss(0) <='1';
          else
          cVar2S5S51P014nsss(0) <='0';
          end if;
        if(cVar1S6S51P033P015N032P017(0)='1' AND  A(12)='1' AND B( 0)='0' AND B( 4)='0' )then
          cVar2S6S51P014P037P029nsss(0) <='1';
          else
          cVar2S6S51P014P037P029nsss(0) <='0';
          end if;
        if(cVar1S7S51P033P015N032P017(0)='1' AND  A(16)='0' AND D(12)='1' AND D( 1)='0' )then
          cVar2S7S51P006P051P062nsss(0) <='1';
          else
          cVar2S7S51P006P051P062nsss(0) <='0';
          end if;
        if(cVar1S8S51P033P015N032P017(0)='1' AND  A(16)='0' AND D(12)='0' AND E( 3)='1' )then
          cVar2S8S51P006N051P056nsss(0) <='1';
          else
          cVar2S8S51P006N051P056nsss(0) <='0';
          end if;
        if(cVar1S9S51P033P015N032P017(0)='1' AND  A(16)='1' AND D( 8)='1' AND A( 0)='1' )then
          cVar2S9S51P006P067P019nsss(0) <='1';
          else
          cVar2S9S51P006P067P019nsss(0) <='0';
          end if;
        if(cVar1S10S51P033N015P059P049(0)='1' AND  A(10)='1' AND A(12)='0' )then
          cVar2S10S51P018P014nsss(0) <='1';
          else
          cVar2S10S51P018P014nsss(0) <='0';
          end if;
        if(cVar1S11S51P033N015P059P049(0)='1' AND  A(10)='1' AND A(12)='1' AND E( 0)='1' )then
          cVar2S11S51P018P014P068nsss(0) <='1';
          else
          cVar2S11S51P018P014P068nsss(0) <='0';
          end if;
        if(cVar1S12S51P033N015P059P049(0)='1' AND  A(10)='0' AND A( 6)='1' AND A(11)='0' )then
          cVar2S12S51N018P007P016nsss(0) <='1';
          else
          cVar2S12S51N018P007P016nsss(0) <='0';
          end if;
        if(cVar1S13S51P033N015P059P049(0)='1' AND  A(10)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar2S13S51N018N007P009nsss(0) <='1';
          else
          cVar2S13S51N018N007P009nsss(0) <='0';
          end if;
        if(cVar1S14S51P033N015P059N049(0)='1' AND  D( 5)='1' AND D( 6)='0' AND E( 4)='0' )then
          cVar2S14S51P046P042P052nsss(0) <='1';
          else
          cVar2S14S51P046P042P052nsss(0) <='0';
          end if;
        if(cVar1S15S51P033N015P059N049(0)='1' AND  D( 5)='0' AND E( 7)='1' )then
          cVar2S15S51N046P040nsss(0) <='1';
          else
          cVar2S15S51N046P040nsss(0) <='0';
          end if;
        if(cVar1S16S51P033N015P059N049(0)='1' AND  D( 5)='0' AND E( 7)='0' AND E( 6)='1' )then
          cVar2S16S51N046N040P044nsss(0) <='1';
          else
          cVar2S16S51N046N040P044nsss(0) <='0';
          end if;
        if(cVar1S17S51P033N015P059P032(0)='1' AND  D( 1)='0' AND A( 1)='1' AND E(11)='0' )then
          cVar2S17S51P062P017P057nsss(0) <='1';
          else
          cVar2S17S51P062P017P057nsss(0) <='0';
          end if;
        if(cVar1S18S51P033N015P059P032(0)='1' AND  D( 1)='0' AND A( 1)='0' AND A(12)='1' )then
          cVar2S18S51P062N017P014nsss(0) <='1';
          else
          cVar2S18S51P062N017P014nsss(0) <='0';
          end if;
        if(cVar1S19S51P033N015P059P032(0)='1' AND  D( 1)='1' AND E( 8)='1' )then
          cVar2S19S51P062P069nsss(0) <='1';
          else
          cVar2S19S51P062P069nsss(0) <='0';
          end if;
        if(cVar1S20S51P033N015P059N032(0)='1' AND  B(12)='1' AND D(11)='0' )then
          cVar2S20S51P030P055nsss(0) <='1';
          else
          cVar2S20S51P030P055nsss(0) <='0';
          end if;
        if(cVar1S21S51P033N015P059N032(0)='1' AND  B(12)='1' AND D(11)='1' AND A(13)='1' )then
          cVar2S21S51P030P055P012nsss(0) <='1';
          else
          cVar2S21S51P030P055P012nsss(0) <='0';
          end if;
        if(cVar1S22S51P033N015P059N032(0)='1' AND  B(12)='0' AND B(10)='1' AND E( 2)='1' )then
          cVar2S22S51N030P034P060nsss(0) <='1';
          else
          cVar2S22S51N030P034P060nsss(0) <='0';
          end if;
        if(cVar1S23S51P033N015P059N032(0)='1' AND  B(12)='0' AND B(10)='0' AND A(15)='1' )then
          cVar2S23S51N030N034P008nsss(0) <='1';
          else
          cVar2S23S51N030N034P008nsss(0) <='0';
          end if;
        if(cVar1S24S51P033P056P016P060(0)='1' AND  A( 4)='0' AND B(12)='0' )then
          cVar2S24S51P011P030nsss(0) <='1';
          else
          cVar2S24S51P011P030nsss(0) <='0';
          end if;
        if(cVar1S25S51P033P056P016P060(0)='1' AND  A( 4)='1' AND D( 3)='1' )then
          cVar2S25S51P011P054nsss(0) <='1';
          else
          cVar2S25S51P011P054nsss(0) <='0';
          end if;
        if(cVar1S26S51P033P056P016P060(0)='1' AND  E(11)='0' AND A( 3)='1' )then
          cVar2S26S51P057P013nsss(0) <='1';
          else
          cVar2S26S51P057P013nsss(0) <='0';
          end if;
        if(cVar1S27S51P033P056P016P060(0)='1' AND  E(11)='0' AND A( 3)='0' AND D( 3)='1' )then
          cVar2S27S51P057N013P054nsss(0) <='1';
          else
          cVar2S27S51P057N013P054nsss(0) <='0';
          end if;
        if(cVar1S28S51P033P056P016P058(0)='1' AND  E( 9)='0' AND A( 1)='0' )then
          cVar2S28S51P065P017nsss(0) <='1';
          else
          cVar2S28S51P065P017nsss(0) <='0';
          end if;
        if(cVar1S30S51P033N056P006N042(0)='1' AND  B(13)='1' )then
          cVar2S30S51P028nsss(0) <='1';
          else
          cVar2S30S51P028nsss(0) <='0';
          end if;
        if(cVar1S31S51P033N056P006N042(0)='1' AND  B(13)='0' AND A(13)='0' AND D(10)='1' )then
          cVar2S31S51N028P012P059nsss(0) <='1';
          else
          cVar2S31S51N028P012P059nsss(0) <='0';
          end if;
        if(cVar1S0S52P006P017P064P037(0)='1' AND  E(13)='0' AND E( 3)='0' )then
          cVar2S0S52P049P056nsss(0) <='1';
          else
          cVar2S0S52P049P056nsss(0) <='0';
          end if;
        if(cVar1S1S52P006P017P064P037(0)='1' AND  E(13)='0' AND E( 3)='1' AND B( 1)='1' )then
          cVar2S1S52P049P056P035nsss(0) <='1';
          else
          cVar2S1S52P049P056P035nsss(0) <='0';
          end if;
        if(cVar1S2S52P006P017P064N037(0)='1' AND  A( 8)='1' AND E( 8)='0' )then
          cVar2S2S52P003P069nsss(0) <='1';
          else
          cVar2S2S52P003P069nsss(0) <='0';
          end if;
        if(cVar1S3S52P006P017P064N037(0)='1' AND  A( 8)='0' AND D( 5)='1' )then
          cVar2S3S52N003P046nsss(0) <='1';
          else
          cVar2S3S52N003P046nsss(0) <='0';
          end if;
        if(cVar1S4S52P006P017P064N037(0)='1' AND  A( 8)='0' AND D( 5)='0' AND D( 1)='1' )then
          cVar2S4S52N003N046P062nsss(0) <='1';
          else
          cVar2S4S52N003N046P062nsss(0) <='0';
          end if;
        if(cVar1S5S52P006P017N064P005(0)='1' AND  A( 3)='0' AND B(12)='0' )then
          cVar2S5S52P013P030nsss(0) <='1';
          else
          cVar2S5S52P013P030nsss(0) <='0';
          end if;
        if(cVar1S6S52P006P017N064P005(0)='1' AND  A( 3)='0' AND B(12)='1' AND D( 1)='1' )then
          cVar2S6S52P013P030P062nsss(0) <='1';
          else
          cVar2S6S52P013P030P062nsss(0) <='0';
          end if;
        if(cVar1S7S52P006P017N064P005(0)='1' AND  A( 3)='1' AND A( 8)='0' AND B( 3)='1' )then
          cVar2S7S52P013P003P031nsss(0) <='1';
          else
          cVar2S7S52P013P003P031nsss(0) <='0';
          end if;
        if(cVar1S8S52P006P017N064P005(0)='1' AND  B( 5)='1' )then
          cVar2S8S52P027nsss(0) <='1';
          else
          cVar2S8S52P027nsss(0) <='0';
          end if;
        if(cVar1S9S52P006P017N064P005(0)='1' AND  B( 5)='0' AND B(15)='1' )then
          cVar2S9S52N027P024nsss(0) <='1';
          else
          cVar2S9S52N027P024nsss(0) <='0';
          end if;
        if(cVar1S10S52P006N017P059P044(0)='1' AND  A(12)='1' AND A( 2)='0' )then
          cVar2S10S52P014P015nsss(0) <='1';
          else
          cVar2S10S52P014P015nsss(0) <='0';
          end if;
        if(cVar1S11S52P006N017P059P044(0)='1' AND  A(12)='1' AND A( 2)='1' AND D( 2)='1' )then
          cVar2S11S52P014P015P058nsss(0) <='1';
          else
          cVar2S11S52P014P015P058nsss(0) <='0';
          end if;
        if(cVar1S12S52P006N017P059P044(0)='1' AND  A(12)='0' AND A( 6)='1' AND A( 2)='0' )then
          cVar2S12S52N014P007P015nsss(0) <='1';
          else
          cVar2S12S52N014P007P015nsss(0) <='0';
          end if;
        if(cVar1S13S52P006N017P059P044(0)='1' AND  A(12)='0' AND A( 6)='0' AND A(11)='1' )then
          cVar2S13S52N014N007P016nsss(0) <='1';
          else
          cVar2S13S52N014N007P016nsss(0) <='0';
          end if;
        if(cVar1S14S52P006N017P059P044(0)='1' AND  A(17)='1' AND B( 9)='0' AND E(14)='0' )then
          cVar2S14S52P004P036P045nsss(0) <='1';
          else
          cVar2S14S52P004P036P045nsss(0) <='0';
          end if;
        if(cVar1S15S52P006N017P059P044(0)='1' AND  A(17)='0' AND A( 7)='1' AND D( 8)='0' )then
          cVar2S15S52N004P005P067nsss(0) <='1';
          else
          cVar2S15S52N004P005P067nsss(0) <='0';
          end if;
        if(cVar1S16S52P006N017P059P060(0)='1' AND  B( 2)='1' )then
          cVar2S16S52P033nsss(0) <='1';
          else
          cVar2S16S52P033nsss(0) <='0';
          end if;
        if(cVar1S17S52P006N017P059P060(0)='1' AND  B( 2)='0' AND B(11)='1' AND E(13)='0' )then
          cVar2S17S52N033P032P049nsss(0) <='1';
          else
          cVar2S17S52N033P032P049nsss(0) <='0';
          end if;
        if(cVar1S18S52P006N017P059P060(0)='1' AND  E( 1)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar2S18S52P064P012P054nsss(0) <='1';
          else
          cVar2S18S52P064P012P054nsss(0) <='0';
          end if;
        if(cVar1S19S52P006N017P059P060(0)='1' AND  E( 1)='1' AND A(12)='0' AND A( 2)='1' )then
          cVar2S19S52P064P014P015nsss(0) <='1';
          else
          cVar2S19S52P064P014P015nsss(0) <='0';
          end if;
        if(cVar1S22S52P006N042P047P064(0)='1' AND  A( 5)='1' )then
          cVar2S22S52P009nsss(0) <='1';
          else
          cVar2S22S52P009nsss(0) <='0';
          end if;
        if(cVar1S23S52P006N042P047P064(0)='1' AND  A( 5)='0' AND B(15)='1' AND D( 5)='0' )then
          cVar2S23S52N009P024P046nsss(0) <='1';
          else
          cVar2S23S52N009P024P046nsss(0) <='0';
          end if;
        if(cVar1S24S52P006N042P047P064(0)='1' AND  A( 5)='0' AND B(15)='0' AND E( 5)='1' )then
          cVar2S24S52N009N024P048nsss(0) <='1';
          else
          cVar2S24S52N009N024P048nsss(0) <='0';
          end if;
        if(cVar1S25S52P006N042N047P043(0)='1' AND  E(14)='1' )then
          cVar2S25S52P045nsss(0) <='1';
          else
          cVar2S25S52P045nsss(0) <='0';
          end if;
        if(cVar1S26S52P006N042N047N043(0)='1' AND  D(12)='1' AND B( 9)='0' AND B( 0)='1' )then
          cVar2S26S52P051P036P037nsss(0) <='1';
          else
          cVar2S26S52P051P036P037nsss(0) <='0';
          end if;
        if(cVar1S27S52P006N042N047N043(0)='1' AND  D(12)='0' AND B( 2)='0' AND D( 2)='1' )then
          cVar2S27S52N051P033P058nsss(0) <='1';
          else
          cVar2S27S52N051P033P058nsss(0) <='0';
          end if;
        if(cVar1S0S53P016P059P017P061(0)='1' AND  B( 4)='1' AND B(12)='0' )then
          cVar2S0S53P029P030nsss(0) <='1';
          else
          cVar2S0S53P029P030nsss(0) <='0';
          end if;
        if(cVar1S1S53P016P059P017P061(0)='1' AND  B( 4)='1' AND B(12)='1' AND A(13)='1' )then
          cVar2S1S53P029P030P012nsss(0) <='1';
          else
          cVar2S1S53P029P030P012nsss(0) <='0';
          end if;
        if(cVar1S2S53P016P059P017P061(0)='1' AND  B( 4)='0' AND A( 0)='1' AND E( 6)='0' )then
          cVar2S2S53N029P019P044nsss(0) <='1';
          else
          cVar2S2S53N029P019P044nsss(0) <='0';
          end if;
        if(cVar1S3S53P016P059P017P061(0)='1' AND  B( 4)='0' AND A( 0)='0' )then
          cVar2S3S53N029N019psss(0) <='1';
          else
          cVar2S3S53N029N019psss(0) <='0';
          end if;
        if(cVar1S4S53P016P059P017P061(0)='1' AND  A(10)='1' AND A(14)='0' AND B( 9)='0' )then
          cVar2S4S53P018P010P036nsss(0) <='1';
          else
          cVar2S4S53P018P010P036nsss(0) <='0';
          end if;
        if(cVar1S5S53P016P059P017P061(0)='1' AND  A(10)='0' AND D( 3)='1' )then
          cVar2S5S53N018P054nsss(0) <='1';
          else
          cVar2S5S53N018P054nsss(0) <='0';
          end if;
        if(cVar1S6S53P016P059P017P061(0)='1' AND  A(10)='0' AND D( 3)='0' AND E(12)='1' )then
          cVar2S6S53N018N054P053nsss(0) <='1';
          else
          cVar2S6S53N018N054P053nsss(0) <='0';
          end if;
        if(cVar1S7S53P016P059P017P015(0)='1' AND  A( 0)='0' AND A(10)='1' AND B( 1)='0' )then
          cVar2S7S53P019P018P035nsss(0) <='1';
          else
          cVar2S7S53P019P018P035nsss(0) <='0';
          end if;
        if(cVar1S8S53P016P059P017P015(0)='1' AND  A( 0)='0' AND A(10)='0' AND B( 0)='1' )then
          cVar2S8S53P019N018P037nsss(0) <='1';
          else
          cVar2S8S53P019N018P037nsss(0) <='0';
          end if;
        if(cVar1S9S53P016P059P017P015(0)='1' AND  A( 0)='1' AND A(10)='0' )then
          cVar2S9S53P019P018nsss(0) <='1';
          else
          cVar2S9S53P019P018nsss(0) <='0';
          end if;
        if(cVar1S10S53P016P059P017P015(0)='1' AND  A( 0)='1' AND A(10)='1' AND A(17)='1' )then
          cVar2S10S53P019P018P004nsss(0) <='1';
          else
          cVar2S10S53P019P018P004nsss(0) <='0';
          end if;
        if(cVar1S11S53P016P059P017P015(0)='1' AND  D( 0)='1' AND B(10)='0' )then
          cVar2S11S53P066P034nsss(0) <='1';
          else
          cVar2S11S53P066P034nsss(0) <='0';
          end if;
        if(cVar1S12S53P016P059P017P015(0)='1' AND  D( 0)='1' AND B(10)='1' AND A(13)='1' )then
          cVar2S12S53P066P034P012nsss(0) <='1';
          else
          cVar2S12S53P066P034P012nsss(0) <='0';
          end if;
        if(cVar1S13S53P016P059P017P015(0)='1' AND  D( 0)='0' AND E(12)='1' )then
          cVar2S13S53N066P053nsss(0) <='1';
          else
          cVar2S13S53N066P053nsss(0) <='0';
          end if;
        if(cVar1S14S53P016P059P017P015(0)='1' AND  D( 0)='0' AND E(12)='0' AND E(13)='1' )then
          cVar2S14S53N066N053P049nsss(0) <='1';
          else
          cVar2S14S53N066N053P049nsss(0) <='0';
          end if;
        if(cVar1S15S53P016P059P015P019(0)='1' AND  B( 2)='1' )then
          cVar2S15S53P033nsss(0) <='1';
          else
          cVar2S15S53P033nsss(0) <='0';
          end if;
        if(cVar1S16S53P016P059P015P019(0)='1' AND  B( 2)='0' AND E(10)='1' )then
          cVar2S16S53N033P061nsss(0) <='1';
          else
          cVar2S16S53N033P061nsss(0) <='0';
          end if;
        if(cVar1S17S53P016P059P015P019(0)='1' AND  B( 2)='0' AND E(10)='0' AND A(10)='0' )then
          cVar2S17S53N033N061P018nsss(0) <='1';
          else
          cVar2S17S53N033N061P018nsss(0) <='0';
          end if;
        if(cVar1S18S53P016P059P015N019(0)='1' AND  D( 2)='0' AND E( 8)='0' )then
          cVar2S18S53P058P069nsss(0) <='1';
          else
          cVar2S18S53P058P069nsss(0) <='0';
          end if;
        if(cVar1S19S53P016P059P015N019(0)='1' AND  D( 2)='0' AND E( 8)='1' AND A( 3)='1' )then
          cVar2S19S53P058P069P013nsss(0) <='1';
          else
          cVar2S19S53P058P069P013nsss(0) <='0';
          end if;
        if(cVar1S20S53P016P059P015N019(0)='1' AND  D( 2)='1' AND B(10)='0' AND B( 0)='1' )then
          cVar2S20S53P058P034P037nsss(0) <='1';
          else
          cVar2S20S53P058P034P037nsss(0) <='0';
          end if;
        if(cVar1S21S53P016P059N015P066(0)='1' AND  D( 1)='0' AND E(10)='1' )then
          cVar2S21S53P062P061nsss(0) <='1';
          else
          cVar2S21S53P062P061nsss(0) <='0';
          end if;
        if(cVar1S22S53P016P059N015P066(0)='1' AND  D( 1)='0' AND E(10)='0' AND D( 4)='1' )then
          cVar2S22S53P062N061P050nsss(0) <='1';
          else
          cVar2S22S53P062N061P050nsss(0) <='0';
          end if;
        if(cVar1S23S53P016P059N015P066(0)='1' AND  D( 1)='1' AND A( 3)='1' AND B(11)='1' )then
          cVar2S23S53P062P013P032nsss(0) <='1';
          else
          cVar2S23S53P062P013P032nsss(0) <='0';
          end if;
        if(cVar1S24S53P016P059N015P066(0)='1' AND  D( 1)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar2S24S53P062N013P011nsss(0) <='1';
          else
          cVar2S24S53P062N013P011nsss(0) <='0';
          end if;
        if(cVar1S25S53P016P059N015P066(0)='1' AND  A(12)='1' AND E(10)='0' )then
          cVar2S25S53P014P061nsss(0) <='1';
          else
          cVar2S25S53P014P061nsss(0) <='0';
          end if;
        if(cVar1S26S53P016P038P002P021(0)='1' AND  D( 3)='0' AND E( 2)='1' AND B( 1)='1' )then
          cVar2S26S53P054P060P035nsss(0) <='1';
          else
          cVar2S26S53P054P060P035nsss(0) <='0';
          end if;
        if(cVar1S27S53P016P038P002P021(0)='1' AND  D( 3)='0' AND E( 2)='0' AND B( 0)='1' )then
          cVar2S27S53P054N060P037nsss(0) <='1';
          else
          cVar2S27S53P054N060P037nsss(0) <='0';
          end if;
        if(cVar1S28S53P016P038P002P021(0)='1' AND  D( 3)='1' AND B( 1)='1' AND E( 3)='1' )then
          cVar2S28S53P054P035P056nsss(0) <='1';
          else
          cVar2S28S53P054P035P056nsss(0) <='0';
          end if;
        if(cVar1S29S53P016P038P002P021(0)='1' AND  D( 3)='1' AND B( 1)='0' AND A(14)='1' )then
          cVar2S29S53P054N035P010nsss(0) <='1';
          else
          cVar2S29S53P054N035P010nsss(0) <='0';
          end if;
        if(cVar1S30S53P016P038P002P021(0)='1' AND  B(14)='0' AND A( 7)='1' AND D( 0)='0' )then
          cVar2S30S53P026P005P066nsss(0) <='1';
          else
          cVar2S30S53P026P005P066nsss(0) <='0';
          end if;
        if(cVar1S31S53P016P038P002P019(0)='1' AND  B( 2)='0' AND E( 9)='1' )then
          cVar2S31S53P033P065nsss(0) <='1';
          else
          cVar2S31S53P033P065nsss(0) <='0';
          end if;
        if(cVar1S32S53P016P038P002P019(0)='1' AND  B( 2)='0' AND E( 9)='0' AND A( 6)='1' )then
          cVar2S32S53P033N065P007nsss(0) <='1';
          else
          cVar2S32S53P033N065P007nsss(0) <='0';
          end if;
        if(cVar1S33S53P016P038P002N019(0)='1' AND  D( 1)='1' AND D( 9)='0' )then
          cVar2S33S53P062P063nsss(0) <='1';
          else
          cVar2S33S53P062P063nsss(0) <='0';
          end if;
        if(cVar1S34S53P016P038P002N019(0)='1' AND  D( 1)='0' AND E(10)='0' AND A(15)='1' )then
          cVar2S34S53N062P061P008nsss(0) <='1';
          else
          cVar2S34S53N062P061P008nsss(0) <='0';
          end if;
        if(cVar1S35S53P016P038P033P064(0)='1' AND  A(15)='1' )then
          cVar2S35S53P008nsss(0) <='1';
          else
          cVar2S35S53P008nsss(0) <='0';
          end if;
        if(cVar1S36S53P016P038P033P064(0)='1' AND  A(15)='0' AND E( 8)='1' )then
          cVar2S36S53N008P069nsss(0) <='1';
          else
          cVar2S36S53N008P069nsss(0) <='0';
          end if;
        if(cVar1S37S53P016P038P033P064(0)='1' AND  A(15)='0' AND E( 8)='0' AND D( 0)='1' )then
          cVar2S37S53N008N069P066nsss(0) <='1';
          else
          cVar2S37S53N008N069P066nsss(0) <='0';
          end if;
        if(cVar1S0S54P037P016P038P002(0)='1' AND  B( 9)='1' AND E( 6)='0' AND A(13)='0' )then
          cVar2S0S54P036P044P012nsss(0) <='1';
          else
          cVar2S0S54P036P044P012nsss(0) <='0';
          end if;
        if(cVar1S1S54P037P016P038P002(0)='1' AND  B( 9)='0' AND A(17)='0' AND E( 7)='0' )then
          cVar2S1S54N036P004P040nsss(0) <='1';
          else
          cVar2S1S54N036P004P040nsss(0) <='0';
          end if;
        if(cVar1S2S54P037P016P038P002(0)='1' AND  B( 9)='0' AND A(17)='1' AND D( 6)='1' )then
          cVar2S2S54N036P004P042nsss(0) <='1';
          else
          cVar2S2S54N036P004P042nsss(0) <='0';
          end if;
        if(cVar1S3S54P037P016P038P002(0)='1' AND  B(15)='0' AND B( 7)='1' )then
          cVar2S3S54P024P023nsss(0) <='1';
          else
          cVar2S3S54P024P023nsss(0) <='0';
          end if;
        if(cVar1S4S54P037P016P038P002(0)='1' AND  B(15)='0' AND B( 7)='0' AND B( 4)='1' )then
          cVar2S4S54P024N023P029nsss(0) <='1';
          else
          cVar2S4S54P024N023P029nsss(0) <='0';
          end if;
        if(cVar1S5S54P037P016P038P033(0)='1' AND  E( 8)='1' )then
          cVar2S5S54P069nsss(0) <='1';
          else
          cVar2S5S54P069nsss(0) <='0';
          end if;
        if(cVar1S6S54P037P016P038P033(0)='1' AND  E( 8)='0' AND E( 7)='1' AND A(10)='1' )then
          cVar2S6S54N069P040P018nsss(0) <='1';
          else
          cVar2S6S54N069P040P018nsss(0) <='0';
          end if;
        if(cVar1S7S54P037N016P050P046(0)='1' AND  B(11)='0' AND A(18)='0' )then
          cVar2S7S54P032P002nsss(0) <='1';
          else
          cVar2S7S54P032P002nsss(0) <='0';
          end if;
        if(cVar1S8S54P037N016P050P046(0)='1' AND  B(11)='1' AND A( 2)='0' AND A(12)='0' )then
          cVar2S8S54P032P015P014nsss(0) <='1';
          else
          cVar2S8S54P032P015P014nsss(0) <='0';
          end if;
        if(cVar1S9S54P037N016P050P046(0)='1' AND  E( 5)='1' AND E( 4)='1' )then
          cVar2S9S54P048P052nsss(0) <='1';
          else
          cVar2S9S54P048P052nsss(0) <='0';
          end if;
        if(cVar1S10S54P037N016N050P039(0)='1' AND  B(17)='1' AND A( 7)='1' )then
          cVar2S10S54P020P005nsss(0) <='1';
          else
          cVar2S10S54P020P005nsss(0) <='0';
          end if;
        if(cVar1S11S54P037N016N050P039(0)='1' AND  B(17)='1' AND A( 7)='0' AND D( 7)='0' )then
          cVar2S11S54P020N005P038nsss(0) <='1';
          else
          cVar2S11S54P020N005P038nsss(0) <='0';
          end if;
        if(cVar1S12S54P037N016N050P039(0)='1' AND  B(17)='0' AND A(15)='0' AND D( 8)='1' )then
          cVar2S12S54N020P008P067nsss(0) <='1';
          else
          cVar2S12S54N020P008P067nsss(0) <='0';
          end if;
        if(cVar1S13S54P037N016N050N039(0)='1' AND  D(12)='1' AND E( 1)='0' )then
          cVar2S13S54P051P064nsss(0) <='1';
          else
          cVar2S13S54P051P064nsss(0) <='0';
          end if;
        if(cVar1S14S54P037N016N050N039(0)='1' AND  D(12)='0' AND A( 1)='1' AND A(10)='1' )then
          cVar2S14S54N051P017P018nsss(0) <='1';
          else
          cVar2S14S54N051P017P018nsss(0) <='0';
          end if;
        if(cVar1S15S54P037P018P060P031(0)='1' AND  A(19)='1' AND A( 5)='0' )then
          cVar2S15S54P000P009nsss(0) <='1';
          else
          cVar2S15S54P000P009nsss(0) <='0';
          end if;
        if(cVar1S16S54P037P018P060P031(0)='1' AND  A(19)='0' AND A(11)='0' AND A( 1)='0' )then
          cVar2S16S54N000P016P017nsss(0) <='1';
          else
          cVar2S16S54N000P016P017nsss(0) <='0';
          end if;
        if(cVar1S17S54P037P018P060P031(0)='1' AND  A(19)='0' AND A(11)='1' AND E( 8)='0' )then
          cVar2S17S54N000P016P069nsss(0) <='1';
          else
          cVar2S17S54N000P016P069nsss(0) <='0';
          end if;
        if(cVar1S18S54P037P018P060P031(0)='1' AND  A( 3)='1' AND D( 1)='1' )then
          cVar2S18S54P013P062nsss(0) <='1';
          else
          cVar2S18S54P013P062nsss(0) <='0';
          end if;
        if(cVar1S19S54P037P018P060P031(0)='1' AND  A( 3)='1' AND D( 1)='0' AND A( 2)='1' )then
          cVar2S19S54P013N062P015nsss(0) <='1';
          else
          cVar2S19S54P013N062P015nsss(0) <='0';
          end if;
        if(cVar1S20S54P037P018P060P031(0)='1' AND  A( 3)='0' AND A( 0)='1' AND A( 2)='0' )then
          cVar2S20S54N013P019P015nsss(0) <='1';
          else
          cVar2S20S54N013P019P015nsss(0) <='0';
          end if;
        if(cVar1S21S54P037P018P060P066(0)='1' AND  D(10)='1' )then
          cVar2S21S54P059nsss(0) <='1';
          else
          cVar2S21S54P059nsss(0) <='0';
          end if;
        if(cVar1S22S54P037P018P060P066(0)='1' AND  D(10)='0' AND D( 9)='1' )then
          cVar2S22S54N059P063nsss(0) <='1';
          else
          cVar2S22S54N059P063nsss(0) <='0';
          end if;
        if(cVar1S23S54P037P018P060P066(0)='1' AND  D(10)='0' AND D( 9)='0' AND A( 5)='1' )then
          cVar2S23S54N059N063P009nsss(0) <='1';
          else
          cVar2S23S54N059N063P009nsss(0) <='0';
          end if;
        if(cVar1S24S54P037P018P060N066(0)='1' AND  A(12)='1' AND A( 2)='0' )then
          cVar2S24S54P014P015nsss(0) <='1';
          else
          cVar2S24S54P014P015nsss(0) <='0';
          end if;
        if(cVar1S25S54P037N018P017P065(0)='1' AND  B( 9)='0' AND A( 6)='0' AND A(17)='0' )then
          cVar2S25S54P036P007P004nsss(0) <='1';
          else
          cVar2S25S54P036P007P004nsss(0) <='0';
          end if;
        if(cVar1S26S54P037N018P017P065(0)='1' AND  B( 9)='0' AND A( 6)='1' AND D( 0)='0' )then
          cVar2S26S54P036P007P066nsss(0) <='1';
          else
          cVar2S26S54P036P007P066nsss(0) <='0';
          end if;
        if(cVar1S27S54P037N018P017P065(0)='1' AND  B( 9)='1' AND A(14)='1' AND A( 0)='1' )then
          cVar2S27S54P036P010P019nsss(0) <='1';
          else
          cVar2S27S54P036P010P019nsss(0) <='0';
          end if;
        if(cVar1S28S54P037N018P017P065(0)='1' AND  A(13)='1' AND D( 0)='1' )then
          cVar2S28S54P012P066nsss(0) <='1';
          else
          cVar2S28S54P012P066nsss(0) <='0';
          end if;
        if(cVar1S29S54P037N018P017P065(0)='1' AND  A(13)='1' AND D( 0)='0' AND A(12)='1' )then
          cVar2S29S54P012N066P014nsss(0) <='1';
          else
          cVar2S29S54P012N066P014nsss(0) <='0';
          end if;
        if(cVar1S30S54P037N018P017P065(0)='1' AND  A(13)='0' AND A(14)='1' )then
          cVar2S30S54N012P010nsss(0) <='1';
          else
          cVar2S30S54N012P010nsss(0) <='0';
          end if;
        if(cVar1S31S54P037N018P017P065(0)='1' AND  A(13)='0' AND A(14)='0' AND B(11)='1' )then
          cVar2S31S54N012N010P032nsss(0) <='1';
          else
          cVar2S31S54N012N010P032nsss(0) <='0';
          end if;
        if(cVar1S32S54P037N018N017P064(0)='1' AND  B(10)='1' AND A(16)='0' AND A( 7)='0' )then
          cVar2S32S54P034P006P005nsss(0) <='1';
          else
          cVar2S32S54P034P006P005nsss(0) <='0';
          end if;
        if(cVar1S33S54P037N018N017P064(0)='1' AND  B(10)='0' AND D( 9)='1' AND E( 8)='0' )then
          cVar2S33S54N034P063P069nsss(0) <='1';
          else
          cVar2S33S54N034P063P069nsss(0) <='0';
          end if;
        if(cVar1S34S54P037N018N017P064(0)='1' AND  B( 6)='1' )then
          cVar2S34S54P025nsss(0) <='1';
          else
          cVar2S34S54P025nsss(0) <='0';
          end if;
        if(cVar1S35S54P037N018N017P064(0)='1' AND  B( 6)='0' AND A(17)='1' AND A(12)='1' )then
          cVar2S35S54N025P004P014nsss(0) <='1';
          else
          cVar2S35S54N025P004P014nsss(0) <='0';
          end if;
        if(cVar1S0S55P016P037P062P001(0)='1' AND  E(15)='1' AND E( 9)='0' )then
          cVar2S0S55P041P065nsss(0) <='1';
          else
          cVar2S0S55P041P065nsss(0) <='0';
          end if;
        if(cVar1S1S55P016P037P062P001(0)='1' AND  E(15)='1' AND E( 9)='1' AND A(10)='0' )then
          cVar2S1S55P041P065P018nsss(0) <='1';
          else
          cVar2S1S55P041P065P018nsss(0) <='0';
          end if;
        if(cVar1S2S55P016P037P062P001(0)='1' AND  E(15)='0' AND A( 8)='0' AND B(17)='0' )then
          cVar2S2S55N041P003P020nsss(0) <='1';
          else
          cVar2S2S55N041P003P020nsss(0) <='0';
          end if;
        if(cVar1S3S55P016P037P062P001(0)='1' AND  E(15)='0' AND A( 8)='1' AND D(14)='1' )then
          cVar2S3S55N041P003P043nsss(0) <='1';
          else
          cVar2S3S55N041P003P043nsss(0) <='0';
          end if;
        if(cVar1S4S55P016P037P062P001(0)='1' AND  D( 8)='1' AND A(14)='0' AND E( 9)='1' )then
          cVar2S4S55P067P010P065nsss(0) <='1';
          else
          cVar2S4S55P067P010P065nsss(0) <='0';
          end if;
        if(cVar1S5S55P016P037P062P047(0)='1' AND  B( 1)='1' AND B(15)='0' )then
          cVar2S5S55P035P024nsss(0) <='1';
          else
          cVar2S5S55P035P024nsss(0) <='0';
          end if;
        if(cVar1S6S55P016P037P062P047(0)='1' AND  B( 1)='0' AND D( 2)='0' AND B( 2)='1' )then
          cVar2S6S55N035P058P033nsss(0) <='1';
          else
          cVar2S6S55N035P058P033nsss(0) <='0';
          end if;
        if(cVar1S7S55P016P037P062P047(0)='1' AND  B(14)='1' )then
          cVar2S7S55P026nsss(0) <='1';
          else
          cVar2S7S55P026nsss(0) <='0';
          end if;
        if(cVar1S9S55P016P037P017N008(0)='1' AND  D( 8)='0' AND B( 1)='1' AND E( 0)='0' )then
          cVar2S9S55P067P035P068nsss(0) <='1';
          else
          cVar2S9S55P067P035P068nsss(0) <='0';
          end if;
        if(cVar1S10S55P016P037P017N008(0)='1' AND  D( 8)='0' AND B( 1)='0' AND E( 0)='1' )then
          cVar2S10S55P067N035P068nsss(0) <='1';
          else
          cVar2S10S55P067N035P068nsss(0) <='0';
          end if;
        if(cVar1S11S55P016P037P017N008(0)='1' AND  D( 8)='1' AND D( 1)='1' AND E( 1)='1' )then
          cVar2S11S55P067P062P064nsss(0) <='1';
          else
          cVar2S11S55P067P062P064nsss(0) <='0';
          end if;
        if(cVar1S12S55P016P037P017N008(0)='1' AND  D( 8)='1' AND D( 1)='0' AND A(12)='1' )then
          cVar2S12S55P067N062P014nsss(0) <='1';
          else
          cVar2S12S55P067N062P014nsss(0) <='0';
          end if;
        if(cVar1S13S55P016P037N017P067(0)='1' AND  D( 9)='0' AND E( 5)='0' )then
          cVar2S13S55P063P048nsss(0) <='1';
          else
          cVar2S13S55P063P048nsss(0) <='0';
          end if;
        if(cVar1S14S55P016P037N017P067(0)='1' AND  D( 9)='1' AND B(10)='1' AND D( 0)='0' )then
          cVar2S14S55P063P034P066nsss(0) <='1';
          else
          cVar2S14S55P063P034P066nsss(0) <='0';
          end if;
        if(cVar1S15S55P016P037N017N067(0)='1' AND  A( 0)='1' AND A( 2)='0' AND B(10)='1' )then
          cVar2S15S55P019P015P034nsss(0) <='1';
          else
          cVar2S15S55P019P015P034nsss(0) <='0';
          end if;
        if(cVar1S16S55P016P037N017N067(0)='1' AND  A( 0)='1' AND A( 2)='1' AND A( 3)='1' )then
          cVar2S16S55P019P015P013nsss(0) <='1';
          else
          cVar2S16S55P019P015P013nsss(0) <='0';
          end if;
        if(cVar1S17S55P016P037N017N067(0)='1' AND  A( 0)='0' AND E( 9)='0' AND A(17)='1' )then
          cVar2S17S55N019P065P004nsss(0) <='1';
          else
          cVar2S17S55N019P065P004nsss(0) <='0';
          end if;
        if(cVar1S18S55P016P036P038P037(0)='1' AND  D( 5)='0' AND D(11)='1' AND B(10)='0' )then
          cVar2S18S55P046P055P034nsss(0) <='1';
          else
          cVar2S18S55P046P055P034nsss(0) <='0';
          end if;
        if(cVar1S19S55P016P036P038P037(0)='1' AND  D( 5)='0' AND D(11)='0' AND B( 5)='0' )then
          cVar2S19S55P046N055P027nsss(0) <='1';
          else
          cVar2S19S55P046N055P027nsss(0) <='0';
          end if;
        if(cVar1S20S55P016P036P038P037(0)='1' AND  D( 5)='1' AND A( 0)='1' )then
          cVar2S20S55P046P019nsss(0) <='1';
          else
          cVar2S20S55P046P019nsss(0) <='0';
          end if;
        if(cVar1S21S55P016P036P038P037(0)='1' AND  A(14)='1' AND E( 9)='1' )then
          cVar2S21S55P010P065nsss(0) <='1';
          else
          cVar2S21S55P010P065nsss(0) <='0';
          end if;
        if(cVar1S22S55P016P036P038P037(0)='1' AND  A(14)='1' AND E( 9)='0' AND D( 8)='1' )then
          cVar2S22S55P010N065P067nsss(0) <='1';
          else
          cVar2S22S55P010N065P067nsss(0) <='0';
          end if;
        if(cVar1S23S55P016P036P038P037(0)='1' AND  A(14)='0' AND B( 4)='0' AND D( 1)='1' )then
          cVar2S23S55N010P029P062nsss(0) <='1';
          else
          cVar2S23S55N010P029P062nsss(0) <='0';
          end if;
        if(cVar1S25S55P016N036P046N024(0)='1' AND  D(13)='0' AND A(10)='0' )then
          cVar2S25S55P047P018nsss(0) <='1';
          else
          cVar2S25S55P047P018nsss(0) <='0';
          end if;
        if(cVar1S26S55P016N036P046N024(0)='1' AND  D(13)='0' AND A(10)='1' AND B( 0)='0' )then
          cVar2S26S55P047P018P037nsss(0) <='1';
          else
          cVar2S26S55P047P018P037nsss(0) <='0';
          end if;
        if(cVar1S27S55P016N036N046P025(0)='1' AND  D( 3)='0' AND A(19)='0' AND D( 6)='1' )then
          cVar2S27S55P054P000P042nsss(0) <='1';
          else
          cVar2S27S55P054P000P042nsss(0) <='0';
          end if;
        if(cVar1S28S55P016N036N046P025(0)='1' AND  D( 3)='1' AND B( 1)='1' AND A( 3)='0' )then
          cVar2S28S55P054P035P013nsss(0) <='1';
          else
          cVar2S28S55P054P035P013nsss(0) <='0';
          end if;
        if(cVar1S29S55P016N036N046P025(0)='1' AND  D( 3)='1' AND B( 1)='0' AND A(14)='1' )then
          cVar2S29S55P054N035P010nsss(0) <='1';
          else
          cVar2S29S55P054N035P010nsss(0) <='0';
          end if;
        if(cVar1S30S55P016N036N046P025(0)='1' AND  A(16)='1' )then
          cVar2S30S55P006nsss(0) <='1';
          else
          cVar2S30S55P006nsss(0) <='0';
          end if;
        if(cVar1S31S55P016N036N046P025(0)='1' AND  A(16)='0' AND A(15)='1' )then
          cVar2S31S55N006P008nsss(0) <='1';
          else
          cVar2S31S55N006P008nsss(0) <='0';
          end if;
        if(cVar1S0S56P016P036P054P000(0)='1' AND  E( 2)='1' AND E( 7)='0' AND E( 5)='0' )then
          cVar2S0S56P060P040P048nsss(0) <='1';
          else
          cVar2S0S56P060P040P048nsss(0) <='0';
          end if;
        if(cVar1S1S56P016P036P054P000(0)='1' AND  E( 2)='0' AND D( 2)='0' AND B( 3)='0' )then
          cVar2S1S56N060P058P031nsss(0) <='1';
          else
          cVar2S1S56N060P058P031nsss(0) <='0';
          end if;
        if(cVar1S2S56P016P036P054P000(0)='1' AND  E( 2)='0' AND D( 2)='1' AND E(11)='1' )then
          cVar2S2S56N060P058P057nsss(0) <='1';
          else
          cVar2S2S56N060P058P057nsss(0) <='0';
          end if;
        if(cVar1S3S56P016P036P054P000(0)='1' AND  D( 1)='1' AND A( 1)='1' )then
          cVar2S3S56P062P017nsss(0) <='1';
          else
          cVar2S3S56P062P017nsss(0) <='0';
          end if;
        if(cVar1S4S56P016P036P054P000(0)='1' AND  D( 1)='0' AND E( 9)='0' AND B( 0)='1' )then
          cVar2S4S56N062P065P037nsss(0) <='1';
          else
          cVar2S4S56N062P065P037nsss(0) <='0';
          end if;
        if(cVar1S5S56P016P036P054P052(0)='1' AND  B( 0)='0' AND E( 9)='0' )then
          cVar2S5S56P037P065nsss(0) <='1';
          else
          cVar2S5S56P037P065nsss(0) <='0';
          end if;
        if(cVar1S6S56P016P036P054P052(0)='1' AND  B( 0)='0' AND E( 9)='1' AND A(10)='1' )then
          cVar2S6S56P037P065P018nsss(0) <='1';
          else
          cVar2S6S56P037P065P018nsss(0) <='0';
          end if;
        if(cVar1S7S56P016P036P054P052(0)='1' AND  B( 0)='1' AND E( 9)='1' )then
          cVar2S7S56P037P065nsss(0) <='1';
          else
          cVar2S7S56P037P065nsss(0) <='0';
          end if;
        if(cVar1S8S56P016P036P054P052(0)='1' AND  D( 0)='0' AND A( 3)='1' )then
          cVar2S8S56P066P013nsss(0) <='1';
          else
          cVar2S8S56P066P013nsss(0) <='0';
          end if;
        if(cVar1S9S56P016P036P054P052(0)='1' AND  D( 0)='0' AND A( 3)='0' AND A( 0)='1' )then
          cVar2S9S56P066N013P019nsss(0) <='1';
          else
          cVar2S9S56P066N013P019nsss(0) <='0';
          end if;
        if(cVar1S11S56P016P036N043P005(0)='1' AND  B(17)='0' AND D(11)='1' AND D(10)='0' )then
          cVar2S11S56P020P055P059nsss(0) <='1';
          else
          cVar2S11S56P020P055P059nsss(0) <='0';
          end if;
        if(cVar1S12S56P016P036N043P005(0)='1' AND  D( 1)='1' AND A(12)='0' )then
          cVar2S12S56P062P014nsss(0) <='1';
          else
          cVar2S12S56P062P014nsss(0) <='0';
          end if;
        if(cVar1S13S56P016P036N043P005(0)='1' AND  D( 1)='0' AND A( 8)='1' )then
          cVar2S13S56N062P003nsss(0) <='1';
          else
          cVar2S13S56N062P003nsss(0) <='0';
          end if;
        if(cVar1S14S56N016P053P051P057(0)='1' AND  E( 2)='0' )then
          cVar2S14S56P060nsss(0) <='1';
          else
          cVar2S14S56P060nsss(0) <='0';
          end if;
        if(cVar1S15S56N016P053P051P057(0)='1' AND  E( 2)='1' AND A( 4)='1' )then
          cVar2S15S56P060P011nsss(0) <='1';
          else
          cVar2S15S56P060P011nsss(0) <='0';
          end if;
        if(cVar1S16S56N016P053P051N057(0)='1' AND  E( 3)='1' AND D( 0)='1' )then
          cVar2S16S56P056P066nsss(0) <='1';
          else
          cVar2S16S56P056P066nsss(0) <='0';
          end if;
        if(cVar1S17S56N016P053P051N057(0)='1' AND  E( 3)='1' AND D( 0)='0' AND E( 1)='0' )then
          cVar2S17S56P056N066P064nsss(0) <='1';
          else
          cVar2S17S56P056N066P064nsss(0) <='0';
          end if;
        if(cVar1S18S56N016P053P051P057(0)='1' AND  D(10)='1' )then
          cVar2S18S56P059nsss(0) <='1';
          else
          cVar2S18S56P059nsss(0) <='0';
          end if;
        if(cVar1S19S56N016P053P051P057(0)='1' AND  D(10)='0' AND A(10)='1' AND E(13)='1' )then
          cVar2S19S56N059P018P049nsss(0) <='1';
          else
          cVar2S19S56N059P018P049nsss(0) <='0';
          end if;
        if(cVar1S20S56N016P053P028P066(0)='1' AND  E( 2)='0' AND A( 3)='1' )then
          cVar2S20S56P060P013nsss(0) <='1';
          else
          cVar2S20S56P060P013nsss(0) <='0';
          end if;
        if(cVar1S21S56N016P053P028P066(0)='1' AND  E( 2)='0' AND A( 3)='0' AND E( 4)='0' )then
          cVar2S21S56P060N013P052nsss(0) <='1';
          else
          cVar2S21S56P060N013P052nsss(0) <='0';
          end if;
        if(cVar1S22S56N016P053P028P066(0)='1' AND  E( 2)='1' AND A( 2)='1' )then
          cVar2S22S56P060P015nsss(0) <='1';
          else
          cVar2S22S56P060P015nsss(0) <='0';
          end if;
        if(cVar1S23S56N016P053P028P066(0)='1' AND  D(12)='0' )then
          cVar2S23S56P051nsss(0) <='1';
          else
          cVar2S23S56P051nsss(0) <='0';
          end if;
        if(cVar1S24S56N016P053P028P066(0)='1' AND  D(12)='1' AND A( 1)='1' )then
          cVar2S24S56P051P017nsss(0) <='1';
          else
          cVar2S24S56P051P017nsss(0) <='0';
          end if;
        if(cVar1S25S56N016P053N028P066(0)='1' AND  D(12)='1' AND E( 8)='0' )then
          cVar2S25S56P051P069nsss(0) <='1';
          else
          cVar2S25S56P051P069nsss(0) <='0';
          end if;
        if(cVar1S26S56N016P053N028P066(0)='1' AND  D(12)='0' AND B( 9)='1' )then
          cVar2S26S56N051P036nsss(0) <='1';
          else
          cVar2S26S56N051P036nsss(0) <='0';
          end if;
        if(cVar1S27S56N016P053N028P066(0)='1' AND  D(12)='0' AND B( 9)='0' AND B(10)='1' )then
          cVar2S27S56N051N036P034nsss(0) <='1';
          else
          cVar2S27S56N051N036P034nsss(0) <='0';
          end if;
        if(cVar1S28S56N016P053N028N066(0)='1' AND  E(13)='0' AND B(14)='1' AND A( 4)='0' )then
          cVar2S28S56P049P026P011nsss(0) <='1';
          else
          cVar2S28S56P049P026P011nsss(0) <='0';
          end if;
        if(cVar1S29S56N016P053N028N066(0)='1' AND  E(13)='0' AND B(14)='0' AND B(10)='1' )then
          cVar2S29S56P049N026P034nsss(0) <='1';
          else
          cVar2S29S56P049N026P034nsss(0) <='0';
          end if;
        if(cVar1S0S57P056P051P016P053(0)='1' AND  B(17)='1' AND A( 7)='1' AND A( 3)='0' )then
          cVar2S0S57P020P005P013nsss(0) <='1';
          else
          cVar2S0S57P020P005P013nsss(0) <='0';
          end if;
        if(cVar1S1S57P056P051P016P053(0)='1' AND  B(17)='1' AND A( 7)='0' AND A( 1)='0' )then
          cVar2S1S57P020N005P017nsss(0) <='1';
          else
          cVar2S1S57P020N005P017nsss(0) <='0';
          end if;
        if(cVar1S2S57P056P051P016P053(0)='1' AND  B(17)='0' AND A( 0)='1' AND E(15)='0' )then
          cVar2S2S57N020P019P041nsss(0) <='1';
          else
          cVar2S2S57N020P019P041nsss(0) <='0';
          end if;
        if(cVar1S3S57P056P051P016P053(0)='1' AND  B(17)='0' AND A( 0)='0' AND A( 1)='1' )then
          cVar2S3S57N020N019P017nsss(0) <='1';
          else
          cVar2S3S57N020N019P017nsss(0) <='0';
          end if;
        if(cVar1S4S57P056P051P016P053(0)='1' AND  B(13)='1' AND D(11)='1' AND E(11)='0' )then
          cVar2S4S57P028P055P057nsss(0) <='1';
          else
          cVar2S4S57P028P055P057nsss(0) <='0';
          end if;
        if(cVar1S5S57P056P051P016P053(0)='1' AND  B(13)='0' AND B( 4)='1' AND A(10)='0' )then
          cVar2S5S57N028P029P018nsss(0) <='1';
          else
          cVar2S5S57N028P029P018nsss(0) <='0';
          end if;
        if(cVar1S6S57P056P051P016P036(0)='1' AND  A( 7)='0' AND B(17)='0' AND A( 0)='1' )then
          cVar2S6S57P005P020P019nsss(0) <='1';
          else
          cVar2S6S57P005P020P019nsss(0) <='0';
          end if;
        if(cVar1S7S57P056P051P016P036(0)='1' AND  A( 7)='1' AND D( 1)='1' AND A(12)='0' )then
          cVar2S7S57P005P062P014nsss(0) <='1';
          else
          cVar2S7S57P005P062P014nsss(0) <='0';
          end if;
        if(cVar1S8S57P056P051P016P036(0)='1' AND  A( 7)='1' AND D( 1)='0' AND A(14)='1' )then
          cVar2S8S57P005N062P010nsss(0) <='1';
          else
          cVar2S8S57P005N062P010nsss(0) <='0';
          end if;
        if(cVar1S9S57P056P051P016N036(0)='1' AND  D( 3)='0' AND E( 2)='1' AND A(15)='0' )then
          cVar2S9S57P054P060P008nsss(0) <='1';
          else
          cVar2S9S57P054P060P008nsss(0) <='0';
          end if;
        if(cVar1S10S57P056P051P016N036(0)='1' AND  D( 3)='0' AND E( 2)='0' AND E(11)='1' )then
          cVar2S10S57P054N060P057nsss(0) <='1';
          else
          cVar2S10S57P054N060P057nsss(0) <='0';
          end if;
        if(cVar1S11S57P056P051P016N036(0)='1' AND  D( 3)='1' AND A(12)='1' AND A( 1)='1' )then
          cVar2S11S57P054P014P017nsss(0) <='1';
          else
          cVar2S11S57P054P014P017nsss(0) <='0';
          end if;
        if(cVar1S12S57P056P051P016N036(0)='1' AND  D( 3)='1' AND A(12)='0' AND B(10)='1' )then
          cVar2S12S57P054N014P034nsss(0) <='1';
          else
          cVar2S12S57P054N014P034nsss(0) <='0';
          end if;
        if(cVar1S13S57P056P051P008P036(0)='1' AND  B(14)='1' )then
          cVar2S13S57P026nsss(0) <='1';
          else
          cVar2S13S57P026nsss(0) <='0';
          end if;
        if(cVar1S14S57P056P051P008P036(0)='1' AND  B(14)='0' AND A( 0)='0' )then
          cVar2S14S57N026P019nsss(0) <='1';
          else
          cVar2S14S57N026P019nsss(0) <='0';
          end if;
        if(cVar1S15S57P056P051P008N036(0)='1' AND  D( 8)='1' )then
          cVar2S15S57P067nsss(0) <='1';
          else
          cVar2S15S57P067nsss(0) <='0';
          end if;
        if(cVar1S16S57P056P051P008N036(0)='1' AND  D( 8)='0' AND D(11)='1' )then
          cVar2S16S57N067P055nsss(0) <='1';
          else
          cVar2S16S57N067P055nsss(0) <='0';
          end if;
        if(cVar1S17S57P056P051P008N036(0)='1' AND  D( 8)='0' AND D(11)='0' AND D(10)='1' )then
          cVar2S17S57N067N055P059nsss(0) <='1';
          else
          cVar2S17S57N067N055P059nsss(0) <='0';
          end if;
        if(cVar1S18S57P056P051N008P064(0)='1' AND  A(11)='1' AND D(10)='0' AND B( 2)='0' )then
          cVar2S18S57P016P059P033nsss(0) <='1';
          else
          cVar2S18S57P016P059P033nsss(0) <='0';
          end if;
        if(cVar1S19S57P056P051N008P064(0)='1' AND  A(11)='0' AND A( 2)='1' AND A(10)='1' )then
          cVar2S19S57N016P015P018nsss(0) <='1';
          else
          cVar2S19S57N016P015P018nsss(0) <='0';
          end if;
        if(cVar1S20S57P056P051N008P064(0)='1' AND  E( 0)='0' AND B( 1)='1' AND A( 3)='1' )then
          cVar2S20S57P068P035P013nsss(0) <='1';
          else
          cVar2S20S57P068P035P013nsss(0) <='0';
          end if;
        if(cVar1S21S57P056P051N008P064(0)='1' AND  E( 0)='0' AND B( 1)='0' AND B(14)='1' )then
          cVar2S21S57P068N035P026nsss(0) <='1';
          else
          cVar2S21S57P068N035P026nsss(0) <='0';
          end if;
        if(cVar1S22S57P056P052P027P050(0)='1' AND  A( 7)='0' AND B( 1)='1' )then
          cVar2S22S57P005P035nsss(0) <='1';
          else
          cVar2S22S57P005P035nsss(0) <='0';
          end if;
        if(cVar1S23S57P056P052P027P050(0)='1' AND  A( 7)='0' AND B( 1)='0' AND B( 2)='1' )then
          cVar2S23S57P005N035P033nsss(0) <='1';
          else
          cVar2S23S57P005N035P033nsss(0) <='0';
          end if;
        if(cVar1S24S57P056P052P027P050(0)='1' AND  A( 7)='1' AND A( 5)='0' AND E( 1)='1' )then
          cVar2S24S57P005P009P064nsss(0) <='1';
          else
          cVar2S24S57P005P009P064nsss(0) <='0';
          end if;
        if(cVar1S25S57P056P052P027P050(0)='1' AND  B( 1)='1' )then
          cVar2S25S57P035nsss(0) <='1';
          else
          cVar2S25S57P035nsss(0) <='0';
          end if;
        if(cVar1S28S57P056P052N009N008(0)='1' AND  A(13)='1' AND D( 4)='1' )then
          cVar2S28S57P012P050nsss(0) <='1';
          else
          cVar2S28S57P012P050nsss(0) <='0';
          end if;
        if(cVar1S0S58P017P065P041P062(0)='1' AND  A( 7)='1' )then
          cVar2S0S58P005nsss(0) <='1';
          else
          cVar2S0S58P005nsss(0) <='0';
          end if;
        if(cVar1S1S58P017P065P041P062(0)='1' AND  A( 7)='0' AND B( 7)='1' )then
          cVar2S1S58N005P023nsss(0) <='1';
          else
          cVar2S1S58N005P023nsss(0) <='0';
          end if;
        if(cVar1S2S58P017P065P041P062(0)='1' AND  A( 7)='0' AND B( 7)='0' AND A(17)='1' )then
          cVar2S2S58N005N023P004nsss(0) <='1';
          else
          cVar2S2S58N005N023P004nsss(0) <='0';
          end if;
        if(cVar1S3S58P017P065P041P062(0)='1' AND  D(15)='1' )then
          cVar2S3S58P039nsss(0) <='1';
          else
          cVar2S3S58P039nsss(0) <='0';
          end if;
        if(cVar1S4S58P017P065N041P038(0)='1' AND  A(18)='1' )then
          cVar2S4S58P002nsss(0) <='1';
          else
          cVar2S4S58P002nsss(0) <='0';
          end if;
        if(cVar1S5S58P017P065N041P038(0)='1' AND  A(18)='0' AND B( 8)='1' )then
          cVar2S5S58N002P021nsss(0) <='1';
          else
          cVar2S5S58N002P021nsss(0) <='0';
          end if;
        if(cVar1S6S58P017P065N041N038(0)='1' AND  A( 2)='1' AND B( 9)='0' )then
          cVar2S6S58P015P036nsss(0) <='1';
          else
          cVar2S6S58P015P036nsss(0) <='0';
          end if;
        if(cVar1S7S58P017P065N041N038(0)='1' AND  A( 2)='1' AND B( 9)='1' AND E(10)='1' )then
          cVar2S7S58P015P036P061nsss(0) <='1';
          else
          cVar2S7S58P015P036P061nsss(0) <='0';
          end if;
        if(cVar1S8S58P017P065N041N038(0)='1' AND  A( 2)='0' AND D( 2)='0' )then
          cVar2S8S58N015P058nsss(0) <='1';
          else
          cVar2S8S58N015P058nsss(0) <='0';
          end if;
        if(cVar1S9S58P017P065P063P056(0)='1' AND  B( 1)='1' AND B(10)='0' AND A( 3)='0' )then
          cVar2S9S58P035P034P013nsss(0) <='1';
          else
          cVar2S9S58P035P034P013nsss(0) <='0';
          end if;
        if(cVar1S10S58P017P065P063P056(0)='1' AND  B( 1)='1' AND B(10)='1' AND A(12)='0' )then
          cVar2S10S58P035P034P014nsss(0) <='1';
          else
          cVar2S10S58P035P034P014nsss(0) <='0';
          end if;
        if(cVar1S11S58P017P065P063P056(0)='1' AND  B( 1)='0' AND A( 3)='1' )then
          cVar2S11S58N035P013nsss(0) <='1';
          else
          cVar2S11S58N035P013nsss(0) <='0';
          end if;
        if(cVar1S12S58P017P065P063P056(0)='1' AND  B( 1)='0' AND A( 3)='0' AND A(12)='1' )then
          cVar2S12S58N035N013P014nsss(0) <='1';
          else
          cVar2S12S58N035N013P014nsss(0) <='0';
          end if;
        if(cVar1S13S58P017P065P063P056(0)='1' AND  E( 1)='1' AND A(11)='0' )then
          cVar2S13S58P064P016nsss(0) <='1';
          else
          cVar2S13S58P064P016nsss(0) <='0';
          end if;
        if(cVar1S14S58P017P065P063P056(0)='1' AND  E( 1)='1' AND A(11)='1' AND A( 3)='1' )then
          cVar2S14S58P064P016P013nsss(0) <='1';
          else
          cVar2S14S58P064P016P013nsss(0) <='0';
          end if;
        if(cVar1S15S58P017P065P063P056(0)='1' AND  E( 1)='0' AND B( 0)='1' )then
          cVar2S15S58N064P037nsss(0) <='1';
          else
          cVar2S15S58N064P037nsss(0) <='0';
          end if;
        if(cVar1S16S58P017P065N063P000(0)='1' AND  A(10)='0' )then
          cVar2S16S58P018nsss(0) <='1';
          else
          cVar2S16S58P018nsss(0) <='0';
          end if;
        if(cVar1S17S58P017P065N063N000(0)='1' AND  B(12)='1' AND D(10)='0' )then
          cVar2S17S58P030P059nsss(0) <='1';
          else
          cVar2S17S58P030P059nsss(0) <='0';
          end if;
        if(cVar1S18S58P017P065N063N000(0)='1' AND  B(12)='0' AND A( 2)='1' AND B( 9)='1' )then
          cVar2S18S58N030P015P036nsss(0) <='1';
          else
          cVar2S18S58N030P015P036nsss(0) <='0';
          end if;
        if(cVar1S19S58P017P065N063N000(0)='1' AND  B(12)='0' AND A( 2)='0' AND A( 5)='1' )then
          cVar2S19S58N030N015P009nsss(0) <='1';
          else
          cVar2S19S58N030N015P009nsss(0) <='0';
          end if;
        if(cVar1S20S58P017P064P037P026(0)='1' AND  B( 1)='1' AND A(12)='1' AND B( 2)='0' )then
          cVar2S20S58P035P014P033nsss(0) <='1';
          else
          cVar2S20S58P035P014P033nsss(0) <='0';
          end if;
        if(cVar1S21S58P017P064P037P026(0)='1' AND  B( 1)='1' AND A(12)='0' AND D( 9)='0' )then
          cVar2S21S58P035N014P063nsss(0) <='1';
          else
          cVar2S21S58P035N014P063nsss(0) <='0';
          end if;
        if(cVar1S22S58P017P064P037P026(0)='1' AND  B( 1)='0' AND A(12)='0' AND D( 3)='0' )then
          cVar2S22S58N035P014P054nsss(0) <='1';
          else
          cVar2S22S58N035P014P054nsss(0) <='0';
          end if;
        if(cVar1S23S58P017P064P037P026(0)='1' AND  B( 1)='0' AND A(12)='1' AND E( 0)='1' )then
          cVar2S23S58N035P014P068nsss(0) <='1';
          else
          cVar2S23S58N035P014P068nsss(0) <='0';
          end if;
        if(cVar1S24S58P017P064N037P003(0)='1' AND  A( 3)='0' AND E( 8)='0' AND D( 1)='1' )then
          cVar2S24S58P013P069P062nsss(0) <='1';
          else
          cVar2S24S58P013P069P062nsss(0) <='0';
          end if;
        if(cVar1S25S58P017P064N037P003(0)='1' AND  A( 3)='0' AND E( 8)='1' )then
          cVar2S25S58P013P069psss(0) <='1';
          else
          cVar2S25S58P013P069psss(0) <='0';
          end if;
        if(cVar1S26S58P017P064N037P003(0)='1' AND  A( 3)='1' AND A(11)='0' )then
          cVar2S26S58P013P016nsss(0) <='1';
          else
          cVar2S26S58P013P016nsss(0) <='0';
          end if;
        if(cVar1S27S58P017P064N037N003(0)='1' AND  D( 5)='1' )then
          cVar2S27S58P046nsss(0) <='1';
          else
          cVar2S27S58P046nsss(0) <='0';
          end if;
        if(cVar1S28S58P017N064P063P068(0)='1' AND  A( 0)='0' AND B( 2)='0' )then
          cVar2S28S58P019P033nsss(0) <='1';
          else
          cVar2S28S58P019P033nsss(0) <='0';
          end if;
        if(cVar1S29S58P017N064P063P068(0)='1' AND  A( 0)='0' AND B( 2)='1' AND E(10)='0' )then
          cVar2S29S58P019P033P061nsss(0) <='1';
          else
          cVar2S29S58P019P033P061nsss(0) <='0';
          end if;
        if(cVar1S30S58P017N064P063P068(0)='1' AND  A( 0)='1' AND E( 8)='0' AND A(10)='0' )then
          cVar2S30S58P019P069P018nsss(0) <='1';
          else
          cVar2S30S58P019P069P018nsss(0) <='0';
          end if;
        if(cVar1S31S58P017N064P063P068(0)='1' AND  A(10)='1' AND B( 9)='0' )then
          cVar2S31S58P018P036nsss(0) <='1';
          else
          cVar2S31S58P018P036nsss(0) <='0';
          end if;
        if(cVar1S32S58P017N064P063P068(0)='1' AND  A(10)='0' AND E( 8)='1' AND A(11)='1' )then
          cVar2S32S58N018P069P016nsss(0) <='1';
          else
          cVar2S32S58N018P069P016nsss(0) <='0';
          end if;
        if(cVar1S33S58P017N064N063P036(0)='1' AND  E(14)='0' )then
          cVar2S33S58P045nsss(0) <='1';
          else
          cVar2S33S58P045nsss(0) <='0';
          end if;
        if(cVar1S34S58P017N064N063P036(0)='1' AND  E(14)='1' AND A(10)='0' )then
          cVar2S34S58P045P018nsss(0) <='1';
          else
          cVar2S34S58P045P018nsss(0) <='0';
          end if;
        if(cVar1S35S58P017N064N063N036(0)='1' AND  B( 0)='1' AND A( 2)='1' AND A(17)='0' )then
          cVar2S35S58P037P015P004nsss(0) <='1';
          else
          cVar2S35S58P037P015P004nsss(0) <='0';
          end if;
        if(cVar1S36S58P017N064N063N036(0)='1' AND  B( 0)='0' AND D(13)='1' AND A(12)='0' )then
          cVar2S36S58N037P047P014nsss(0) <='1';
          else
          cVar2S36S58N037P047P014nsss(0) <='0';
          end if;
        if(cVar1S37S58P017N064N063N036(0)='1' AND  B( 0)='0' AND D(13)='0' AND B( 3)='1' )then
          cVar2S37S58N037N047P031nsss(0) <='1';
          else
          cVar2S37S58N037N047P031nsss(0) <='0';
          end if;
        if(cVar1S0S59P063P001P035P015(0)='1' AND  D( 0)='0' AND E( 0)='1' )then
          cVar2S0S59P066P068nsss(0) <='1';
          else
          cVar2S0S59P066P068nsss(0) <='0';
          end if;
        if(cVar1S1S59P063P001P035P015(0)='1' AND  D( 0)='0' AND E( 0)='0' AND E( 3)='0' )then
          cVar2S1S59P066N068P056nsss(0) <='1';
          else
          cVar2S1S59P066N068P056nsss(0) <='0';
          end if;
        if(cVar1S2S59P063P001P035P015(0)='1' AND  D( 0)='1' AND A( 0)='1' )then
          cVar2S2S59P066P019nsss(0) <='1';
          else
          cVar2S2S59P066P019nsss(0) <='0';
          end if;
        if(cVar1S3S59P063P001P035P015(0)='1' AND  B(10)='0' AND A( 1)='0' AND A(10)='0' )then
          cVar2S3S59P034P017P018nsss(0) <='1';
          else
          cVar2S3S59P034P017P018nsss(0) <='0';
          end if;
        if(cVar1S4S59P063P001P035P015(0)='1' AND  B(10)='0' AND A( 1)='1' AND D( 1)='0' )then
          cVar2S4S59P034P017P062nsss(0) <='1';
          else
          cVar2S4S59P034P017P062nsss(0) <='0';
          end if;
        if(cVar1S5S59P063P001N035P057(0)='1' AND  A(13)='1' AND D( 8)='0' AND A(14)='0' )then
          cVar2S5S59P012P067P010nsss(0) <='1';
          else
          cVar2S5S59P012P067P010nsss(0) <='0';
          end if;
        if(cVar1S6S59P063P001N035P057(0)='1' AND  A(13)='1' AND D( 8)='1' AND B(10)='1' )then
          cVar2S6S59P012P067P034nsss(0) <='1';
          else
          cVar2S6S59P012P067P034nsss(0) <='0';
          end if;
        if(cVar1S7S59P063P001N035P057(0)='1' AND  A(13)='0' AND B( 3)='0' AND D( 1)='0' )then
          cVar2S7S59N012P031P062nsss(0) <='1';
          else
          cVar2S7S59N012P031P062nsss(0) <='0';
          end if;
        if(cVar1S8S59P063P001N035P057(0)='1' AND  A(13)='0' AND B( 3)='1' AND E( 9)='0' )then
          cVar2S8S59N012P031P065nsss(0) <='1';
          else
          cVar2S8S59N012P031P065nsss(0) <='0';
          end if;
        if(cVar1S9S59P063P001N035P057(0)='1' AND  A(14)='0' AND D( 3)='0' AND A( 3)='1' )then
          cVar2S9S59P010P054P013nsss(0) <='1';
          else
          cVar2S9S59P010P054P013nsss(0) <='0';
          end if;
        if(cVar1S10S59P063P001P034P068(0)='1' AND  A( 1)='1' )then
          cVar2S10S59P017nsss(0) <='1';
          else
          cVar2S10S59P017nsss(0) <='0';
          end if;
        if(cVar1S11S59N063P060P054P064(0)='1' AND  A( 0)='0' AND B( 1)='0' )then
          cVar2S11S59P019P035nsss(0) <='1';
          else
          cVar2S11S59P019P035nsss(0) <='0';
          end if;
        if(cVar1S12S59N063P060P054P064(0)='1' AND  A( 0)='0' AND B( 1)='1' AND D( 0)='1' )then
          cVar2S12S59P019P035P066nsss(0) <='1';
          else
          cVar2S12S59P019P035P066nsss(0) <='0';
          end if;
        if(cVar1S13S59N063P060P054P064(0)='1' AND  A( 0)='1' AND B(10)='1' AND A(10)='0' )then
          cVar2S13S59P019P034P018nsss(0) <='1';
          else
          cVar2S13S59P019P034P018nsss(0) <='0';
          end if;
        if(cVar1S14S59N063P060P054P064(0)='1' AND  A( 0)='1' AND B(10)='0' AND B( 2)='1' )then
          cVar2S14S59P019N034P033nsss(0) <='1';
          else
          cVar2S14S59P019N034P033nsss(0) <='0';
          end if;
        if(cVar1S15S59N063P060P054P064(0)='1' AND  D(11)='0' AND E(10)='0' AND E( 8)='0' )then
          cVar2S15S59P055P061P069nsss(0) <='1';
          else
          cVar2S15S59P055P061P069nsss(0) <='0';
          end if;
        if(cVar1S16S59N063P060P054P056(0)='1' AND  D( 8)='0' AND B( 1)='1' )then
          cVar2S16S59P067P035nsss(0) <='1';
          else
          cVar2S16S59P067P035nsss(0) <='0';
          end if;
        if(cVar1S17S59N063N060P064P065(0)='1' AND  A(14)='0' AND B( 9)='0' )then
          cVar2S17S59P010P036nsss(0) <='1';
          else
          cVar2S17S59P010P036nsss(0) <='0';
          end if;
        if(cVar1S18S59N063N060P064N065(0)='1' AND  D(12)='0' AND D( 2)='0' AND B( 0)='0' )then
          cVar2S18S59P051P058P037nsss(0) <='1';
          else
          cVar2S18S59P051P058P037nsss(0) <='0';
          end if;
        if(cVar1S19S59N063N060N064P062(0)='1' AND  E(15)='1' AND A(11)='0' )then
          cVar2S19S59P041P016nsss(0) <='1';
          else
          cVar2S19S59P041P016nsss(0) <='0';
          end if;
        if(cVar1S20S59N063N060N064P062(0)='1' AND  E(15)='1' AND A(11)='1' AND A( 3)='1' )then
          cVar2S20S59P041P016P013nsss(0) <='1';
          else
          cVar2S20S59P041P016P013nsss(0) <='0';
          end if;
        if(cVar1S21S59N063N060N064P062(0)='1' AND  E(15)='0' AND D( 7)='1' )then
          cVar2S21S59N041P038nsss(0) <='1';
          else
          cVar2S21S59N041P038nsss(0) <='0';
          end if;
        if(cVar1S22S59N063N060N064P062(0)='1' AND  A(15)='1' AND A( 0)='1' AND A(10)='0' )then
          cVar2S22S59P008P019P018nsss(0) <='1';
          else
          cVar2S22S59P008P019P018nsss(0) <='0';
          end if;
        if(cVar1S23S59N063N060N064P062(0)='1' AND  A(15)='1' AND A( 0)='0' AND A( 3)='1' )then
          cVar2S23S59P008N019P013nsss(0) <='1';
          else
          cVar2S23S59P008N019P013nsss(0) <='0';
          end if;
        if(cVar1S24S59N063N060N064P062(0)='1' AND  A(15)='0' AND A( 4)='1' AND A( 1)='0' )then
          cVar2S24S59N008P011P017nsss(0) <='1';
          else
          cVar2S24S59N008P011P017nsss(0) <='0';
          end if;
        if(cVar1S0S60P037P063P033P017(0)='1' AND  A( 6)='0' AND B( 1)='1' AND B(17)='0' )then
          cVar2S0S60P007P035P020nsss(0) <='1';
          else
          cVar2S0S60P007P035P020nsss(0) <='0';
          end if;
        if(cVar1S1S60P037P063P033P017(0)='1' AND  A( 6)='0' AND B( 1)='0' AND D( 0)='1' )then
          cVar2S1S60P007N035P066nsss(0) <='1';
          else
          cVar2S1S60P007N035P066nsss(0) <='0';
          end if;
        if(cVar1S2S60P037P063P033P017(0)='1' AND  A( 6)='1' AND E(11)='0' AND E( 1)='1' )then
          cVar2S2S60P007P057P064nsss(0) <='1';
          else
          cVar2S2S60P007P057P064nsss(0) <='0';
          end if;
        if(cVar1S3S60P037P063P033N017(0)='1' AND  A(13)='1' AND E( 5)='0' AND D( 0)='1' )then
          cVar2S3S60P012P048P066nsss(0) <='1';
          else
          cVar2S3S60P012P048P066nsss(0) <='0';
          end if;
        if(cVar1S4S60P037P063P033N017(0)='1' AND  A(13)='0' AND A(17)='1' )then
          cVar2S4S60N012P004nsss(0) <='1';
          else
          cVar2S4S60N012P004nsss(0) <='0';
          end if;
        if(cVar1S5S60P037P063P033N017(0)='1' AND  A(13)='0' AND A(17)='0' AND B(14)='1' )then
          cVar2S5S60N012N004P026nsss(0) <='1';
          else
          cVar2S5S60N012N004P026nsss(0) <='0';
          end if;
        if(cVar1S6S60P037P063P033P059(0)='1' AND  A( 2)='1' AND A( 3)='0' )then
          cVar2S6S60P015P013nsss(0) <='1';
          else
          cVar2S6S60P015P013nsss(0) <='0';
          end if;
        if(cVar1S7S60P037P063P033P059(0)='1' AND  A( 2)='0' AND A( 3)='1' )then
          cVar2S7S60N015P013nsss(0) <='1';
          else
          cVar2S7S60N015P013nsss(0) <='0';
          end if;
        if(cVar1S8S60P037P063P033N059(0)='1' AND  D( 8)='1' AND D( 1)='1' AND E( 2)='0' )then
          cVar2S8S60P067P062P060nsss(0) <='1';
          else
          cVar2S8S60P067P062P060nsss(0) <='0';
          end if;
        if(cVar1S9S60P037P063P033N059(0)='1' AND  D( 8)='1' AND D( 1)='0' AND A( 4)='1' )then
          cVar2S9S60P067N062P011nsss(0) <='1';
          else
          cVar2S9S60P067N062P011nsss(0) <='0';
          end if;
        if(cVar1S10S60P037P063P033N059(0)='1' AND  D( 8)='0' AND D( 2)='1' AND A(13)='1' )then
          cVar2S10S60N067P058P012nsss(0) <='1';
          else
          cVar2S10S60N067P058P012nsss(0) <='0';
          end if;
        if(cVar1S11S60P037P063P068P013(0)='1' AND  A(12)='0' AND A(11)='1' )then
          cVar2S11S60P014P016nsss(0) <='1';
          else
          cVar2S11S60P014P016nsss(0) <='0';
          end if;
        if(cVar1S12S60P037P063P068P013(0)='1' AND  A(12)='0' AND A(11)='0' AND A( 1)='1' )then
          cVar2S12S60P014N016P017nsss(0) <='1';
          else
          cVar2S12S60P014N016P017nsss(0) <='0';
          end if;
        if(cVar1S13S60P037P063P068P013(0)='1' AND  A(12)='1' AND A( 4)='0' )then
          cVar2S13S60P014P011nsss(0) <='1';
          else
          cVar2S13S60P014P011nsss(0) <='0';
          end if;
        if(cVar1S14S60P037P063P068N013(0)='1' AND  D( 8)='0' AND E( 9)='0' AND A( 2)='0' )then
          cVar2S14S60P067P065P015nsss(0) <='1';
          else
          cVar2S14S60P067P065P015nsss(0) <='0';
          end if;
        if(cVar1S15S60P037P063P068N013(0)='1' AND  D( 8)='0' AND E( 9)='1' AND D( 0)='1' )then
          cVar2S15S60P067P065P066nsss(0) <='1';
          else
          cVar2S15S60P067P065P066nsss(0) <='0';
          end if;
        if(cVar1S16S60P037P063P068N013(0)='1' AND  D( 8)='1' AND E( 1)='0' AND A(11)='0' )then
          cVar2S16S60P067P064P016nsss(0) <='1';
          else
          cVar2S16S60P067P064P016nsss(0) <='0';
          end if;
        if(cVar1S18S60P037P063P068N052(0)='1' AND  A(13)='1' AND A( 3)='0' )then
          cVar2S18S60P012P013nsss(0) <='1';
          else
          cVar2S18S60P012P013nsss(0) <='0';
          end if;
        if(cVar1S19S60P037P063P068N052(0)='1' AND  A(13)='0' AND D(10)='0' AND B( 2)='1' )then
          cVar2S19S60N012P059P033nsss(0) <='1';
          else
          cVar2S19S60N012P059P033nsss(0) <='0';
          end if;
        if(cVar1S20S60N037P035P065P022(0)='1' AND  A( 6)='1' )then
          cVar2S20S60P007nsss(0) <='1';
          else
          cVar2S20S60P007nsss(0) <='0';
          end if;
        if(cVar1S21S60N037P035P065P022(0)='1' AND  A( 6)='0' AND E( 3)='0' )then
          cVar2S21S60N007P056nsss(0) <='1';
          else
          cVar2S21S60N007P056nsss(0) <='0';
          end if;
        if(cVar1S22S60N037P035P065N022(0)='1' AND  A(12)='0' AND B(15)='1' )then
          cVar2S22S60P014P024nsss(0) <='1';
          else
          cVar2S22S60P014P024nsss(0) <='0';
          end if;
        if(cVar1S23S60N037P035P065N022(0)='1' AND  A(12)='0' AND B(15)='0' AND A( 2)='1' )then
          cVar2S23S60P014N024P015nsss(0) <='1';
          else
          cVar2S23S60P014N024P015nsss(0) <='0';
          end if;
        if(cVar1S24S60N037P035P065N022(0)='1' AND  A(12)='1' AND B( 7)='1' AND E( 8)='0' )then
          cVar2S24S60P014P023P069nsss(0) <='1';
          else
          cVar2S24S60P014P023P069nsss(0) <='0';
          end if;
        if(cVar1S25S60N037P035P065P002(0)='1' AND  B( 9)='1' AND E( 1)='1' )then
          cVar2S25S60P036P064nsss(0) <='1';
          else
          cVar2S25S60P036P064nsss(0) <='0';
          end if;
        if(cVar1S26S60N037P035P065P002(0)='1' AND  B( 9)='1' AND E( 1)='0' AND A( 1)='0' )then
          cVar2S26S60P036N064P017nsss(0) <='1';
          else
          cVar2S26S60P036N064P017nsss(0) <='0';
          end if;
        if(cVar1S27S60N037P035P065P002(0)='1' AND  E( 8)='0' AND B(10)='1' AND A( 1)='1' )then
          cVar2S27S60P069P034P017nsss(0) <='1';
          else
          cVar2S27S60P069P034P017nsss(0) <='0';
          end if;
        if(cVar1S28S60N037P035P065P041(0)='1' AND  D( 8)='1' AND B( 9)='0' )then
          cVar2S28S60P067P036nsss(0) <='1';
          else
          cVar2S28S60P067P036nsss(0) <='0';
          end if;
        if(cVar1S29S60N037P035P065P041(0)='1' AND  D( 8)='1' AND B( 9)='1' AND B(10)='1' )then
          cVar2S29S60P067P036P034nsss(0) <='1';
          else
          cVar2S29S60P067P036P034nsss(0) <='0';
          end if;
        if(cVar1S30S60N037P035P065P041(0)='1' AND  D( 8)='0' AND D(12)='0' AND D( 0)='0' )then
          cVar2S30S60N067P051P066nsss(0) <='1';
          else
          cVar2S30S60N067P051P066nsss(0) <='0';
          end if;
        if(cVar1S31S60N037P035N065P054(0)='1' AND  A(14)='1' )then
          cVar2S31S60P010nsss(0) <='1';
          else
          cVar2S31S60P010nsss(0) <='0';
          end if;
        if(cVar1S32S60N037P035N065P054(0)='1' AND  A(14)='0' AND B( 3)='1' AND A( 2)='0' )then
          cVar2S32S60N010P031P015nsss(0) <='1';
          else
          cVar2S32S60N010P031P015nsss(0) <='0';
          end if;
        if(cVar1S33S60N037P035N065P054(0)='1' AND  A(14)='0' AND B( 3)='0' AND D( 1)='1' )then
          cVar2S33S60N010N031P062nsss(0) <='1';
          else
          cVar2S33S60N010N031P062nsss(0) <='0';
          end if;
        if(cVar1S34S60N037P035N065N054(0)='1' AND  B( 2)='1' AND E( 2)='1' AND A(13)='0' )then
          cVar2S34S60P033P060P012nsss(0) <='1';
          else
          cVar2S34S60P033P060P012nsss(0) <='0';
          end if;
        if(cVar1S35S60N037P035N065N054(0)='1' AND  B( 2)='1' AND E( 2)='0' AND D(11)='1' )then
          cVar2S35S60P033N060P055nsss(0) <='1';
          else
          cVar2S35S60P033N060P055nsss(0) <='0';
          end if;
        if(cVar1S36S60N037P035N065N054(0)='1' AND  B( 2)='0' AND D(11)='1' AND B( 3)='1' )then
          cVar2S36S60N033P055P031nsss(0) <='1';
          else
          cVar2S36S60N033P055P031nsss(0) <='0';
          end if;
        if(cVar1S0S61P063P035P015P017(0)='1' AND  E( 9)='0' AND D(11)='0' )then
          cVar2S0S61P065P055nsss(0) <='1';
          else
          cVar2S0S61P065P055nsss(0) <='0';
          end if;
        if(cVar1S1S61P063P035P015P017(0)='1' AND  E( 9)='0' AND D(11)='1' AND E( 3)='0' )then
          cVar2S1S61P065P055P056nsss(0) <='1';
          else
          cVar2S1S61P065P055P056nsss(0) <='0';
          end if;
        if(cVar1S2S61P063P035P015P017(0)='1' AND  E( 9)='1' AND B(12)='1' )then
          cVar2S2S61P065P030nsss(0) <='1';
          else
          cVar2S2S61P065P030nsss(0) <='0';
          end if;
        if(cVar1S3S61P063P035P015P017(0)='1' AND  E( 9)='1' AND B(12)='0' AND A( 5)='1' )then
          cVar2S3S61P065N030P009nsss(0) <='1';
          else
          cVar2S3S61P065N030P009nsss(0) <='0';
          end if;
        if(cVar1S4S61P063P035P015P017(0)='1' AND  D( 8)='1' AND E( 1)='1' AND E( 0)='0' )then
          cVar2S4S61P067P064P068nsss(0) <='1';
          else
          cVar2S4S61P067P064P068nsss(0) <='0';
          end if;
        if(cVar1S5S61P063P035P015P017(0)='1' AND  D( 8)='1' AND E( 1)='0' )then
          cVar2S5S61P067N064psss(0) <='1';
          else
          cVar2S5S61P067N064psss(0) <='0';
          end if;
        if(cVar1S6S61P063P035P015P017(0)='1' AND  D( 8)='0' AND B( 2)='0' AND E( 8)='0' )then
          cVar2S6S61N067P033P069nsss(0) <='1';
          else
          cVar2S6S61N067P033P069nsss(0) <='0';
          end if;
        if(cVar1S7S61P063P035P015P017(0)='1' AND  D( 8)='0' AND B( 2)='1' AND B(13)='1' )then
          cVar2S7S61N067P033P028nsss(0) <='1';
          else
          cVar2S7S61N067P033P028nsss(0) <='0';
          end if;
        if(cVar1S8S61P063P035P015P025(0)='1' AND  D( 5)='1' )then
          cVar2S8S61P046nsss(0) <='1';
          else
          cVar2S8S61P046nsss(0) <='0';
          end if;
        if(cVar1S9S61P063P035P015P025(0)='1' AND  D( 5)='0' AND E( 0)='1' AND A( 0)='1' )then
          cVar2S9S61N046P068P019nsss(0) <='1';
          else
          cVar2S9S61N046P068P019nsss(0) <='0';
          end if;
        if(cVar1S10S61P063P035P015N025(0)='1' AND  E( 1)='0' AND E(10)='1' )then
          cVar2S10S61P064P061nsss(0) <='1';
          else
          cVar2S10S61P064P061nsss(0) <='0';
          end if;
        if(cVar1S11S61P063P035P015N025(0)='1' AND  E( 1)='1' AND B( 0)='1' AND E( 8)='1' )then
          cVar2S11S61P064P037P069nsss(0) <='1';
          else
          cVar2S11S61P064P037P069nsss(0) <='0';
          end if;
        if(cVar1S12S61P063P035P015N025(0)='1' AND  E( 1)='1' AND B( 0)='0' AND E( 3)='1' )then
          cVar2S12S61P064N037P056nsss(0) <='1';
          else
          cVar2S12S61P064N037P056nsss(0) <='0';
          end if;
        if(cVar1S13S61P063P035P014P047(0)='1' AND  D(10)='0' AND D( 1)='1' AND D(11)='0' )then
          cVar2S13S61P059P062P055nsss(0) <='1';
          else
          cVar2S13S61P059P062P055nsss(0) <='0';
          end if;
        if(cVar1S14S61P063P035P014P047(0)='1' AND  D(10)='0' AND D( 1)='0' AND A( 2)='0' )then
          cVar2S14S61P059N062P015nsss(0) <='1';
          else
          cVar2S14S61P059N062P015nsss(0) <='0';
          end if;
        if(cVar1S15S61P063P035P014P047(0)='1' AND  D(10)='1' AND A(10)='1' AND B(11)='0' )then
          cVar2S15S61P059P018P032nsss(0) <='1';
          else
          cVar2S15S61P059P018P032nsss(0) <='0';
          end if;
        if(cVar1S16S61P063P035N014P061(0)='1' AND  A(13)='0' AND B(11)='0' )then
          cVar2S16S61P012P032nsss(0) <='1';
          else
          cVar2S16S61P012P032nsss(0) <='0';
          end if;
        if(cVar1S17S61P063P035N014P061(0)='1' AND  A(13)='0' AND B(11)='1' AND A(11)='0' )then
          cVar2S17S61P012P032P016nsss(0) <='1';
          else
          cVar2S17S61P012P032P016nsss(0) <='0';
          end if;
        if(cVar1S18S61P063P035N014P061(0)='1' AND  A(13)='1' AND A(10)='1' )then
          cVar2S18S61P012P018nsss(0) <='1';
          else
          cVar2S18S61P012P018nsss(0) <='0';
          end if;
        if(cVar1S19S61P063P035N014N061(0)='1' AND  D( 1)='1' AND E( 3)='1' )then
          cVar2S19S61P062P056nsss(0) <='1';
          else
          cVar2S19S61P062P056nsss(0) <='0';
          end if;
        if(cVar1S20S61P063P035N014N061(0)='1' AND  D( 1)='0' AND E(13)='1' AND D(13)='1' )then
          cVar2S20S61N062P049P047nsss(0) <='1';
          else
          cVar2S20S61N062P049P047nsss(0) <='0';
          end if;
        if(cVar1S21S61P063P035N014N061(0)='1' AND  D( 1)='0' AND E(13)='0' AND E( 4)='1' )then
          cVar2S21S61N062N049P052nsss(0) <='1';
          else
          cVar2S21S61N062N049P052nsss(0) <='0';
          end if;
        if(cVar1S23S61P063P062P068N060(0)='1' AND  D( 8)='1' AND A( 1)='1' )then
          cVar2S23S61P067P017nsss(0) <='1';
          else
          cVar2S23S61P067P017nsss(0) <='0';
          end if;
        if(cVar1S24S61P063P062P068N060(0)='1' AND  D( 8)='1' AND A( 1)='0' AND B(10)='1' )then
          cVar2S24S61P067N017P034nsss(0) <='1';
          else
          cVar2S24S61P067N017P034nsss(0) <='0';
          end if;
        if(cVar1S25S61P063P062P068N060(0)='1' AND  D( 8)='0' AND A(12)='1' AND A(10)='0' )then
          cVar2S25S61N067P014P018nsss(0) <='1';
          else
          cVar2S25S61N067P014P018nsss(0) <='0';
          end if;
        if(cVar1S26S61P063P062N068P022(0)='1' AND  B( 0)='1' AND B(10)='1' AND A(12)='0' )then
          cVar2S26S61P037P034P014nsss(0) <='1';
          else
          cVar2S26S61P037P034P014nsss(0) <='0';
          end if;
        if(cVar1S27S61P063P062N068P022(0)='1' AND  B( 0)='1' AND B(10)='0' AND A(12)='1' )then
          cVar2S27S61P037N034P014nsss(0) <='1';
          else
          cVar2S27S61P037N034P014nsss(0) <='0';
          end if;
        if(cVar1S28S61P063P062N068P022(0)='1' AND  B( 0)='0' AND E( 8)='1' AND D( 8)='0' )then
          cVar2S28S61N037P069P067nsss(0) <='1';
          else
          cVar2S28S61N037P069P067nsss(0) <='0';
          end if;
        if(cVar1S29S61P063P062N068P022(0)='1' AND  B( 0)='0' AND E( 8)='0' AND A(13)='1' )then
          cVar2S29S61N037N069P012nsss(0) <='1';
          else
          cVar2S29S61N037N069P012nsss(0) <='0';
          end if;
        if(cVar1S30S61P063N062P002P035(0)='1' AND  A( 6)='0' AND E(12)='0' AND B( 9)='0' )then
          cVar2S30S61P007P053P036nsss(0) <='1';
          else
          cVar2S30S61P007P053P036nsss(0) <='0';
          end if;
        if(cVar1S31S61P063N062P002N035(0)='1' AND  D( 0)='0' AND E(14)='0' AND B( 6)='0' )then
          cVar2S31S61P066P045P025nsss(0) <='1';
          else
          cVar2S31S61P066P045P025nsss(0) <='0';
          end if;
        if(cVar1S32S61P063N062P002N035(0)='1' AND  D( 0)='1' AND E( 4)='0' AND D( 3)='1' )then
          cVar2S32S61P066P052P054nsss(0) <='1';
          else
          cVar2S32S61P066P052P054nsss(0) <='0';
          end if;
        if(cVar1S33S61P063N062P002P037(0)='1' AND  A( 0)='1' )then
          cVar2S33S61P019nsss(0) <='1';
          else
          cVar2S33S61P019nsss(0) <='0';
          end if;
        if(cVar1S34S61P063N062P002N037(0)='1' AND  D( 8)='0' AND D( 0)='0' AND A( 2)='0' )then
          cVar2S34S61P067P066P015nsss(0) <='1';
          else
          cVar2S34S61P067P066P015nsss(0) <='0';
          end if;
        if(cVar1S0S62P062P017P048P022(0)='1' AND  A(11)='1' AND E( 9)='1' )then
          cVar2S0S62P016P065nsss(0) <='1';
          else
          cVar2S0S62P016P065nsss(0) <='0';
          end if;
        if(cVar1S1S62P062P017P048P022(0)='1' AND  A(11)='1' AND E( 9)='0' AND A( 6)='0' )then
          cVar2S1S62P016N065P007nsss(0) <='1';
          else
          cVar2S1S62P016N065P007nsss(0) <='0';
          end if;
        if(cVar1S2S62P062P017P048P022(0)='1' AND  A(11)='0' AND B( 6)='1' )then
          cVar2S2S62N016P025nsss(0) <='1';
          else
          cVar2S2S62N016P025nsss(0) <='0';
          end if;
        if(cVar1S3S62P062P017P048P022(0)='1' AND  A(11)='0' AND B( 6)='0' AND A(14)='0' )then
          cVar2S3S62N016N025P010nsss(0) <='1';
          else
          cVar2S3S62N016N025P010nsss(0) <='0';
          end if;
        if(cVar1S5S62P062P017P048N046(0)='1' AND  A(11)='1' AND B( 1)='1' )then
          cVar2S5S62P016P035nsss(0) <='1';
          else
          cVar2S5S62P016P035nsss(0) <='0';
          end if;
        if(cVar1S6S62P062N017P047P005(0)='1' AND  E(14)='1' AND A(13)='0' )then
          cVar2S6S62P045P012nsss(0) <='1';
          else
          cVar2S6S62P045P012nsss(0) <='0';
          end if;
        if(cVar1S7S62P062N017P047P005(0)='1' AND  E(14)='0' AND A( 2)='1' AND E(13)='0' )then
          cVar2S7S62N045P015P049nsss(0) <='1';
          else
          cVar2S7S62N045P015P049nsss(0) <='0';
          end if;
        if(cVar1S8S62P062N017P047P005(0)='1' AND  E(14)='0' AND A( 2)='0' AND D( 0)='0' )then
          cVar2S8S62N045N015P066nsss(0) <='1';
          else
          cVar2S8S62N045N015P066nsss(0) <='0';
          end if;
        if(cVar1S9S62P062N017P047P005(0)='1' AND  D(15)='1' )then
          cVar2S9S62P039nsss(0) <='1';
          else
          cVar2S9S62P039nsss(0) <='0';
          end if;
        if(cVar1S10S62P062N017P047P005(0)='1' AND  D(15)='0' AND A(12)='1' AND E( 2)='0' )then
          cVar2S10S62N039P014P060nsss(0) <='1';
          else
          cVar2S10S62N039P014P060nsss(0) <='0';
          end if;
        if(cVar1S12S62P062N017P047N026(0)='1' AND  A( 6)='1' )then
          cVar2S12S62P007nsss(0) <='1';
          else
          cVar2S12S62P007nsss(0) <='0';
          end if;
        if(cVar1S13S62N062P066P067P059(0)='1' AND  B( 2)='0' AND A( 2)='0' )then
          cVar2S13S62P033P015nsss(0) <='1';
          else
          cVar2S13S62P033P015nsss(0) <='0';
          end if;
        if(cVar1S14S62N062P066P067P059(0)='1' AND  B( 2)='0' AND A( 2)='1' AND B( 1)='0' )then
          cVar2S14S62P033P015P035nsss(0) <='1';
          else
          cVar2S14S62P033P015P035nsss(0) <='0';
          end if;
        if(cVar1S15S62N062P066P067P059(0)='1' AND  B( 2)='1' AND D( 2)='1' AND A( 6)='0' )then
          cVar2S15S62P033P058P007nsss(0) <='1';
          else
          cVar2S15S62P033P058P007nsss(0) <='0';
          end if;
        if(cVar1S16S62N062P066P067P059(0)='1' AND  A( 2)='1' AND B(11)='0' AND D( 2)='0' )then
          cVar2S16S62P015P032P058nsss(0) <='1';
          else
          cVar2S16S62P015P032P058nsss(0) <='0';
          end if;
        if(cVar1S17S62N062P066P067P059(0)='1' AND  A( 2)='1' AND B(11)='1' AND A(13)='1' )then
          cVar2S17S62P015P032P012nsss(0) <='1';
          else
          cVar2S17S62P015P032P012nsss(0) <='0';
          end if;
        if(cVar1S18S62N062P066P067P059(0)='1' AND  A( 2)='0' AND B(11)='1' AND E( 2)='0' )then
          cVar2S18S62N015P032P060nsss(0) <='1';
          else
          cVar2S18S62N015P032P060nsss(0) <='0';
          end if;
        if(cVar1S19S62N062P066P067P059(0)='1' AND  A( 2)='0' AND B(11)='0' AND B(12)='1' )then
          cVar2S19S62N015N032P030nsss(0) <='1';
          else
          cVar2S19S62N015N032P030nsss(0) <='0';
          end if;
        if(cVar1S20S62N062P066P067P016(0)='1' AND  B( 9)='0' AND B(10)='0' AND A( 2)='0' )then
          cVar2S20S62P036P034P015nsss(0) <='1';
          else
          cVar2S20S62P036P034P015nsss(0) <='0';
          end if;
        if(cVar1S21S62N062P066P067P016(0)='1' AND  B( 9)='0' AND B(10)='1' AND A(10)='1' )then
          cVar2S21S62P036P034P018nsss(0) <='1';
          else
          cVar2S21S62P036P034P018nsss(0) <='0';
          end if;
        if(cVar1S22S62N062P066P067P016(0)='1' AND  B( 9)='1' AND D(12)='1' )then
          cVar2S22S62P036P051nsss(0) <='1';
          else
          cVar2S22S62P036P051nsss(0) <='0';
          end if;
        if(cVar1S23S62N062P066P067N016(0)='1' AND  D( 2)='1' AND E(10)='0' AND E( 0)='1' )then
          cVar2S23S62P058P061P068nsss(0) <='1';
          else
          cVar2S23S62P058P061P068nsss(0) <='0';
          end if;
        if(cVar1S24S62N062P066P067N016(0)='1' AND  D( 2)='1' AND E(10)='1' AND B(11)='1' )then
          cVar2S24S62P058P061P032nsss(0) <='1';
          else
          cVar2S24S62P058P061P032nsss(0) <='0';
          end if;
        if(cVar1S25S62N062P066P067N016(0)='1' AND  D( 2)='0' AND D(11)='1' AND A( 1)='1' )then
          cVar2S25S62N058P055P017nsss(0) <='1';
          else
          cVar2S25S62N058P055P017nsss(0) <='0';
          end if;
        if(cVar1S26S62N062N066P034P010(0)='1' AND  D( 9)='0' AND E( 1)='0' AND E( 2)='0' )then
          cVar2S26S62P063P064P060nsss(0) <='1';
          else
          cVar2S26S62P063P064P060nsss(0) <='0';
          end if;
        if(cVar1S27S62N062N066P034P010(0)='1' AND  D( 9)='1' AND B( 4)='1' )then
          cVar2S27S62P063P029nsss(0) <='1';
          else
          cVar2S27S62P063P029nsss(0) <='0';
          end if;
        if(cVar1S28S62N062N066P034P010(0)='1' AND  D( 9)='1' AND B( 4)='0' AND E(12)='1' )then
          cVar2S28S62P063N029P053nsss(0) <='1';
          else
          cVar2S28S62P063N029P053nsss(0) <='0';
          end if;
        if(cVar1S29S62N062N066P034N010(0)='1' AND  A(13)='1' AND E( 5)='0' )then
          cVar2S29S62P012P048nsss(0) <='1';
          else
          cVar2S29S62P012P048nsss(0) <='0';
          end if;
        if(cVar1S30S62N062N066P034N010(0)='1' AND  A(13)='1' AND E( 5)='1' AND A( 2)='1' )then
          cVar2S30S62P012P048P015nsss(0) <='1';
          else
          cVar2S30S62P012P048P015nsss(0) <='0';
          end if;
        if(cVar1S31S62N062N066P034N010(0)='1' AND  A(13)='0' AND A(15)='1' AND B(11)='0' )then
          cVar2S31S62N012P008P032nsss(0) <='1';
          else
          cVar2S31S62N012P008P032nsss(0) <='0';
          end if;
        if(cVar1S32S62N062N066P034P016(0)='1' AND  E( 2)='0' AND E( 8)='0' AND D( 6)='0' )then
          cVar2S32S62P060P069P042nsss(0) <='1';
          else
          cVar2S32S62P060P069P042nsss(0) <='0';
          end if;
        if(cVar1S33S62N062N066P034P016(0)='1' AND  E( 2)='1' AND A( 4)='1' )then
          cVar2S33S62P060P011nsss(0) <='1';
          else
          cVar2S33S62P060P011nsss(0) <='0';
          end if;
        if(cVar1S34S62N062N066P034P016(0)='1' AND  E( 2)='1' AND A( 4)='0' AND B(11)='1' )then
          cVar2S34S62P060N011P032nsss(0) <='1';
          else
          cVar2S34S62P060N011P032nsss(0) <='0';
          end if;
        if(cVar1S35S62N062N066P034N016(0)='1' AND  D( 8)='1' AND E( 9)='1' )then
          cVar2S35S62P067P065nsss(0) <='1';
          else
          cVar2S35S62P067P065nsss(0) <='0';
          end if;
        if(cVar1S36S62N062N066P034N016(0)='1' AND  D( 8)='1' AND E( 9)='0' AND E(10)='1' )then
          cVar2S36S62P067N065P061nsss(0) <='1';
          else
          cVar2S36S62P067N065P061nsss(0) <='0';
          end if;
        if(cVar1S37S62N062N066P034N016(0)='1' AND  D( 8)='0' AND E( 0)='1' AND A( 0)='1' )then
          cVar2S37S62N067P068P019nsss(0) <='1';
          else
          cVar2S37S62N067P068P019nsss(0) <='0';
          end if;
        if(cVar1S0S63P067P018P050P062(0)='1' AND  B(13)='0' AND A( 1)='0' )then
          cVar2S0S63P028P017nsss(0) <='1';
          else
          cVar2S0S63P028P017nsss(0) <='0';
          end if;
        if(cVar1S1S63P067P018P050P062(0)='1' AND  B(13)='0' AND A( 1)='1' AND E( 2)='0' )then
          cVar2S1S63P028P017P060nsss(0) <='1';
          else
          cVar2S1S63P028P017P060nsss(0) <='0';
          end if;
        if(cVar1S2S63P067P018P050P062(0)='1' AND  B(13)='1' AND A( 4)='1' AND D( 0)='0' )then
          cVar2S2S63P028P011P066nsss(0) <='1';
          else
          cVar2S2S63P028P011P066nsss(0) <='0';
          end if;
        if(cVar1S3S63P067P018P050P062(0)='1' AND  A( 0)='1' AND A(13)='0' AND A(14)='0' )then
          cVar2S3S63P019P012P010nsss(0) <='1';
          else
          cVar2S3S63P019P012P010nsss(0) <='0';
          end if;
        if(cVar1S4S63P067P018P050P062(0)='1' AND  A( 0)='0' AND A( 3)='1' AND E( 1)='1' )then
          cVar2S4S63N019P013P064nsss(0) <='1';
          else
          cVar2S4S63N019P013P064nsss(0) <='0';
          end if;
        if(cVar1S5S63P067P018P050P010(0)='1' AND  A( 1)='1' )then
          cVar2S5S63P017nsss(0) <='1';
          else
          cVar2S5S63P017nsss(0) <='0';
          end if;
        if(cVar1S6S63P067P018P050N010(0)='1' AND  E( 0)='1' AND B( 4)='1' )then
          cVar2S6S63P068P029nsss(0) <='1';
          else
          cVar2S6S63P068P029nsss(0) <='0';
          end if;
        if(cVar1S7S63P067P018P050N010(0)='1' AND  E( 0)='1' AND B( 4)='0' AND E( 4)='0' )then
          cVar2S7S63P068N029P052nsss(0) <='1';
          else
          cVar2S7S63P068N029P052nsss(0) <='0';
          end if;
        if(cVar1S8S63P067N018P068P049(0)='1' AND  E( 7)='0' AND B(12)='0' AND B( 8)='0' )then
          cVar2S8S63P040P030P021nsss(0) <='1';
          else
          cVar2S8S63P040P030P021nsss(0) <='0';
          end if;
        if(cVar1S9S63P067N018P068P049(0)='1' AND  E( 7)='0' AND B(12)='1' AND A( 2)='1' )then
          cVar2S9S63P040P030P015nsss(0) <='1';
          else
          cVar2S9S63P040P030P015nsss(0) <='0';
          end if;
        if(cVar1S10S63P067N018N068P015(0)='1' AND  B(10)='0' AND E( 1)='0' )then
          cVar2S10S63P034P064nsss(0) <='1';
          else
          cVar2S10S63P034P064nsss(0) <='0';
          end if;
        if(cVar1S11S63P067N018N068P015(0)='1' AND  B(10)='0' AND E( 1)='1' AND A( 1)='0' )then
          cVar2S11S63P034P064P017nsss(0) <='1';
          else
          cVar2S11S63P034P064P017nsss(0) <='0';
          end if;
        if(cVar1S12S63P067N018N068P015(0)='1' AND  B(10)='1' AND E( 8)='1' AND D( 1)='1' )then
          cVar2S12S63P034P069P062nsss(0) <='1';
          else
          cVar2S12S63P034P069P062nsss(0) <='0';
          end if;
        if(cVar1S13S63P067N018N068N015(0)='1' AND  A( 1)='1' AND E( 8)='1' AND A( 8)='0' )then
          cVar2S13S63P017P069P003nsss(0) <='1';
          else
          cVar2S13S63P017P069P003nsss(0) <='0';
          end if;
        if(cVar1S14S63P067N018N068N015(0)='1' AND  A( 1)='0' AND E(14)='1' )then
          cVar2S14S63N017P045nsss(0) <='1';
          else
          cVar2S14S63N017P045nsss(0) <='0';
          end if;
        if(cVar1S15S63P067N018N068N015(0)='1' AND  A( 1)='0' AND E(14)='0' AND D( 7)='1' )then
          cVar2S15S63N017N045P038nsss(0) <='1';
          else
          cVar2S15S63N017N045P038nsss(0) <='0';
          end if;
        if(cVar1S17S63N067P044N028P023(0)='1' AND  A(13)='0' )then
          cVar2S17S63P012nsss(0) <='1';
          else
          cVar2S17S63P012nsss(0) <='0';
          end if;
        if(cVar1S18S63N067P044N028N023(0)='1' AND  B( 6)='1' AND D( 1)='1' )then
          cVar2S18S63P025P062nsss(0) <='1';
          else
          cVar2S18S63P025P062nsss(0) <='0';
          end if;
        if(cVar1S19S63N067P044N028N023(0)='1' AND  B( 6)='1' AND D( 1)='0' AND D( 6)='0' )then
          cVar2S19S63P025N062P042nsss(0) <='1';
          else
          cVar2S19S63P025N062P042nsss(0) <='0';
          end if;
        if(cVar1S20S63N067P044N028N023(0)='1' AND  B( 6)='0' AND E( 9)='1' AND A( 1)='1' )then
          cVar2S20S63N025P065P017nsss(0) <='1';
          else
          cVar2S20S63N025P065P017nsss(0) <='0';
          end if;
        if(cVar1S21S63N067P044N028N023(0)='1' AND  B( 6)='0' AND E( 9)='0' AND A(16)='1' )then
          cVar2S21S63N025N065P006nsss(0) <='1';
          else
          cVar2S21S63N025N065P006nsss(0) <='0';
          end if;
        if(cVar1S22S63N067N044P059P049(0)='1' AND  A(14)='0' AND D(11)='0' AND D( 3)='0' )then
          cVar2S22S63P010P055P054nsss(0) <='1';
          else
          cVar2S22S63P010P055P054nsss(0) <='0';
          end if;
        if(cVar1S23S63N067N044P059P049(0)='1' AND  A(14)='0' AND D(11)='1' AND B(10)='1' )then
          cVar2S23S63P010P055P034nsss(0) <='1';
          else
          cVar2S23S63P010P055P034nsss(0) <='0';
          end if;
        if(cVar1S24S63N067N044P059P049(0)='1' AND  A(14)='1' AND B(15)='0' AND A( 2)='1' )then
          cVar2S24S63P010P024P015nsss(0) <='1';
          else
          cVar2S24S63P010P024P015nsss(0) <='0';
          end if;
        if(cVar1S25S63N067N044P059P049(0)='1' AND  D(12)='1' )then
          cVar2S25S63P051nsss(0) <='1';
          else
          cVar2S25S63P051nsss(0) <='0';
          end if;
        if(cVar1S26S63N067N044N059P031(0)='1' AND  B(12)='0' AND A( 3)='1' )then
          cVar2S26S63P030P013nsss(0) <='1';
          else
          cVar2S26S63P030P013nsss(0) <='0';
          end if;
        if(cVar1S27S63N067N044N059P031(0)='1' AND  B(12)='0' AND A( 3)='0' AND D( 2)='1' )then
          cVar2S27S63P030N013P058nsss(0) <='1';
          else
          cVar2S27S63P030N013P058nsss(0) <='0';
          end if;
        if(cVar1S28S63N067N044N059P031(0)='1' AND  B(12)='1' AND A( 5)='0' AND E( 9)='1' )then
          cVar2S28S63P030P009P065nsss(0) <='1';
          else
          cVar2S28S63P030P009P065nsss(0) <='0';
          end if;
        if(cVar1S29S63N067N044N059N031(0)='1' AND  B(10)='1' AND A(15)='0' AND D( 1)='1' )then
          cVar2S29S63P034P008P062nsss(0) <='1';
          else
          cVar2S29S63P034P008P062nsss(0) <='0';
          end if;
        if(cVar1S30S63N067N044N059N031(0)='1' AND  B(10)='1' AND A(15)='1' AND E(12)='1' )then
          cVar2S30S63P034P008P053nsss(0) <='1';
          else
          cVar2S30S63P034P008P053nsss(0) <='0';
          end if;
        if(cVar1S31S63N067N044N059N031(0)='1' AND  B(10)='0' AND B( 6)='1' AND D(12)='0' )then
          cVar2S31S63N034P025P051nsss(0) <='1';
          else
          cVar2S31S63N034P025P051nsss(0) <='0';
          end if;
        if(cVar1S0S64P059P061P058P032(0)='1' AND  B(12)='0' AND D( 8)='0' AND A(10)='0' )then
          cVar2S0S64P030P067P018nsss(0) <='1';
          else
          cVar2S0S64P030P067P018nsss(0) <='0';
          end if;
        if(cVar1S1S64P059P061P058P032(0)='1' AND  B(12)='0' AND D( 8)='1' AND A( 1)='0' )then
          cVar2S1S64P030P067P017nsss(0) <='1';
          else
          cVar2S1S64P030P067P017nsss(0) <='0';
          end if;
        if(cVar1S2S64P059P061P058N032(0)='1' AND  D( 1)='0' AND D(13)='1' AND D( 0)='0' )then
          cVar2S2S64P062P047P066nsss(0) <='1';
          else
          cVar2S2S64P062P047P066nsss(0) <='0';
          end if;
        if(cVar1S3S64P059P061P058N032(0)='1' AND  D( 1)='0' AND D(13)='0' AND B(14)='0' )then
          cVar2S3S64P062N047P026nsss(0) <='1';
          else
          cVar2S3S64P062N047P026nsss(0) <='0';
          end if;
        if(cVar1S4S64P059P061P058N032(0)='1' AND  D( 1)='1' AND A(16)='0' AND B(12)='1' )then
          cVar2S4S64P062P006P030nsss(0) <='1';
          else
          cVar2S4S64P062P006P030nsss(0) <='0';
          end if;
        if(cVar1S5S64P059P061N058P033(0)='1' AND  E( 2)='0' )then
          cVar2S5S64P060nsss(0) <='1';
          else
          cVar2S5S64P060nsss(0) <='0';
          end if;
        if(cVar1S6S64P059P061N058P033(0)='1' AND  E( 2)='1' AND D( 1)='1' AND E( 1)='0' )then
          cVar2S6S64P060P062P064nsss(0) <='1';
          else
          cVar2S6S64P060P062P064nsss(0) <='0';
          end if;
        if(cVar1S7S64P059P061N058P033(0)='1' AND  B(11)='0' AND E( 2)='1' AND D( 1)='1' )then
          cVar2S7S64P032P060P062nsss(0) <='1';
          else
          cVar2S7S64P032P060P062nsss(0) <='0';
          end if;
        if(cVar1S8S64P059P061N058P033(0)='1' AND  B(11)='0' AND E( 2)='0' AND D(11)='1' )then
          cVar2S8S64P032N060P055nsss(0) <='1';
          else
          cVar2S8S64P032N060P055nsss(0) <='0';
          end if;
        if(cVar1S10S64P059P061P067N069(0)='1' AND  E( 9)='0' AND A( 6)='0' )then
          cVar2S10S64P065P007nsss(0) <='1';
          else
          cVar2S10S64P065P007nsss(0) <='0';
          end if;
        if(cVar1S11S64P059P061P067P037(0)='1' AND  A( 0)='1' )then
          cVar2S11S64P019nsss(0) <='1';
          else
          cVar2S11S64P019nsss(0) <='0';
          end if;
        if(cVar1S12S64P059P049P030P004(0)='1' AND  A( 3)='1' AND B( 1)='0' )then
          cVar2S12S64P013P035nsss(0) <='1';
          else
          cVar2S12S64P013P035nsss(0) <='0';
          end if;
        if(cVar1S13S64P059P049P030P004(0)='1' AND  A( 3)='0' AND E( 3)='1' )then
          cVar2S13S64N013P056nsss(0) <='1';
          else
          cVar2S13S64N013P056nsss(0) <='0';
          end if;
        if(cVar1S14S64P059P049P030P004(0)='1' AND  A( 3)='0' AND E( 3)='0' AND E( 2)='1' )then
          cVar2S14S64N013N056P060nsss(0) <='1';
          else
          cVar2S14S64N013N056P060nsss(0) <='0';
          end if;
        if(cVar1S15S64P059P049N030P005(0)='1' AND  A( 4)='1' AND E( 2)='1' AND E(10)='1' )then
          cVar2S15S64P011P060P061nsss(0) <='1';
          else
          cVar2S15S64P011P060P061nsss(0) <='0';
          end if;
        if(cVar1S16S64P059P049N030P005(0)='1' AND  A( 4)='1' AND E( 2)='0' AND B( 9)='0' )then
          cVar2S16S64P011N060P036nsss(0) <='1';
          else
          cVar2S16S64P011N060P036nsss(0) <='0';
          end if;
        if(cVar1S17S64P059P049N030P005(0)='1' AND  A( 4)='0' AND A(12)='0' AND B( 3)='1' )then
          cVar2S17S64N011N014P031nsss(0) <='1';
          else
          cVar2S17S64N011N014P031nsss(0) <='0';
          end if;
        if(cVar1S18S64P059P049N030P005(0)='1' AND  E( 2)='1' )then
          cVar2S18S64P060nsss(0) <='1';
          else
          cVar2S18S64P060nsss(0) <='0';
          end if;
        if(cVar1S19S64P059P049N030P005(0)='1' AND  E( 2)='0' AND A( 8)='1' )then
          cVar2S19S64N060P003nsss(0) <='1';
          else
          cVar2S19S64N060P003nsss(0) <='0';
          end if;
        if(cVar1S21S64P059P049P055N051(0)='1' AND  B( 2)='1' )then
          cVar2S21S64P033nsss(0) <='1';
          else
          cVar2S21S64P033nsss(0) <='0';
          end if;
        if(cVar1S1S65P058P054P047N026(0)='1' AND  B( 0)='0' AND B(15)='0' AND A(11)='0' )then
          cVar2S1S65P037P024P016nsss(0) <='1';
          else
          cVar2S1S65P037P024P016nsss(0) <='0';
          end if;
        if(cVar1S2S65P058P054N047P013(0)='1' AND  A( 0)='1' AND B( 0)='0' AND B( 1)='0' )then
          cVar2S2S65P019P037P035nsss(0) <='1';
          else
          cVar2S2S65P019P037P035nsss(0) <='0';
          end if;
        if(cVar1S3S65P058P054N047P013(0)='1' AND  A( 0)='1' AND B( 0)='1' AND B( 9)='1' )then
          cVar2S3S65P019P037P036nsss(0) <='1';
          else
          cVar2S3S65P019P037P036nsss(0) <='0';
          end if;
        if(cVar1S4S65P058P054N047P013(0)='1' AND  A( 0)='0' AND A( 6)='0' AND B(13)='0' )then
          cVar2S4S65N019P007P028nsss(0) <='1';
          else
          cVar2S4S65N019P007P028nsss(0) <='0';
          end if;
        if(cVar1S5S65P058P054N047N013(0)='1' AND  A( 8)='1' AND E( 9)='1' )then
          cVar2S5S65P003P065nsss(0) <='1';
          else
          cVar2S5S65P003P065nsss(0) <='0';
          end if;
        if(cVar1S6S65P058P054N047N013(0)='1' AND  A( 8)='1' AND E( 9)='0' AND A( 5)='0' )then
          cVar2S6S65P003N065P009nsss(0) <='1';
          else
          cVar2S6S65P003N065P009nsss(0) <='0';
          end if;
        if(cVar1S7S65P058P054N047N013(0)='1' AND  A( 8)='0' AND A( 5)='1' )then
          cVar2S7S65N003P009nsss(0) <='1';
          else
          cVar2S7S65N003P009nsss(0) <='0';
          end if;
        if(cVar1S9S65P058P054P015N013(0)='1' AND  A(13)='0' AND E( 3)='1' AND B( 2)='1' )then
          cVar2S9S65P012P056P033nsss(0) <='1';
          else
          cVar2S9S65P012P056P033nsss(0) <='0';
          end if;
        if(cVar1S10S65P058P054N015P033(0)='1' AND  A( 4)='1' )then
          cVar2S10S65P011nsss(0) <='1';
          else
          cVar2S10S65P011nsss(0) <='0';
          end if;
        if(cVar1S11S65P058P054N015P033(0)='1' AND  A( 4)='0' AND B( 3)='0' AND A( 3)='1' )then
          cVar2S11S65N011P031P013nsss(0) <='1';
          else
          cVar2S11S65N011P031P013nsss(0) <='0';
          end if;
        if(cVar1S12S65P058P054N015N033(0)='1' AND  B( 9)='0' AND E( 0)='0' AND A( 3)='1' )then
          cVar2S12S65P036P068P013nsss(0) <='1';
          else
          cVar2S12S65P036P068P013nsss(0) <='0';
          end if;
        if(cVar1S14S65N058P043P022N003(0)='1' AND  B(10)='1' )then
          cVar2S14S65P034nsss(0) <='1';
          else
          cVar2S14S65P034nsss(0) <='0';
          end if;
        if(cVar1S15S65N058P043P022N003(0)='1' AND  B(10)='0' AND E( 8)='0' AND E( 1)='0' )then
          cVar2S15S65N034P069P064nsss(0) <='1';
          else
          cVar2S15S65N034P069P064nsss(0) <='0';
          end if;
        if(cVar1S16S65N058P043N022P047(0)='1' AND  A( 6)='1' AND A(11)='1' )then
          cVar2S16S65P007P016nsss(0) <='1';
          else
          cVar2S16S65P007P016nsss(0) <='0';
          end if;
        if(cVar1S17S65N058P043N022P047(0)='1' AND  A( 6)='1' AND A(11)='0' AND E(14)='1' )then
          cVar2S17S65P007N016P045nsss(0) <='1';
          else
          cVar2S17S65P007N016P045nsss(0) <='0';
          end if;
        if(cVar1S18S65N058P043N022P047(0)='1' AND  A( 6)='0' AND B( 8)='1' )then
          cVar2S18S65N007P021nsss(0) <='1';
          else
          cVar2S18S65N007P021nsss(0) <='0';
          end if;
        if(cVar1S19S65N058N043P040P002(0)='1' AND  B( 9)='0' AND B( 8)='1' )then
          cVar2S19S65P036P021nsss(0) <='1';
          else
          cVar2S19S65P036P021nsss(0) <='0';
          end if;
        if(cVar1S20S65N058N043P040P002(0)='1' AND  B( 9)='0' AND B( 8)='0' AND B(17)='1' )then
          cVar2S20S65P036N021P020nsss(0) <='1';
          else
          cVar2S20S65P036N021P020nsss(0) <='0';
          end if;
        if(cVar1S21S65N058N043P040P002(0)='1' AND  B( 9)='1' )then
          cVar2S21S65P036psss(0) <='1';
          else
          cVar2S21S65P036psss(0) <='0';
          end if;
        if(cVar1S22S65N058N043P040N002(0)='1' AND  A(17)='1' AND E( 0)='0' )then
          cVar2S22S65P004P068nsss(0) <='1';
          else
          cVar2S22S65P004P068nsss(0) <='0';
          end if;
        if(cVar1S23S65N058N043P040N002(0)='1' AND  A(17)='0' AND B( 0)='1' AND D( 1)='1' )then
          cVar2S23S65N004P037P062nsss(0) <='1';
          else
          cVar2S23S65N004P037P062nsss(0) <='0';
          end if;
        if(cVar1S24S65N058N043N040P038(0)='1' AND  D(15)='1' AND B(17)='1' )then
          cVar2S24S65P039P020nsss(0) <='1';
          else
          cVar2S24S65P039P020nsss(0) <='0';
          end if;
        if(cVar1S25S65N058N043N040P038(0)='1' AND  D(15)='1' AND B(17)='0' AND B( 8)='1' )then
          cVar2S25S65P039N020P021nsss(0) <='1';
          else
          cVar2S25S65P039N020P021nsss(0) <='0';
          end if;
        if(cVar1S26S65N058N043N040P038(0)='1' AND  D(15)='0' AND B( 8)='1' AND D(13)='1' )then
          cVar2S26S65N039P021P047nsss(0) <='1';
          else
          cVar2S26S65N039P021P047nsss(0) <='0';
          end if;
        if(cVar1S27S65N058N043N040P038(0)='1' AND  B( 0)='1' AND E( 8)='0' AND D( 0)='1' )then
          cVar2S27S65P037P069P066nsss(0) <='1';
          else
          cVar2S27S65P037P069P066nsss(0) <='0';
          end if;
        if(cVar1S2S66P015P044N025N023(0)='1' AND  D( 2)='0' AND B(16)='1' )then
          cVar2S2S66P058P022nsss(0) <='1';
          else
          cVar2S2S66P058P022nsss(0) <='0';
          end if;
        if(cVar1S3S66P015P044N025N023(0)='1' AND  D( 2)='0' AND B(16)='0' AND E( 0)='1' )then
          cVar2S3S66P058N022P068nsss(0) <='1';
          else
          cVar2S3S66P058N022P068nsss(0) <='0';
          end if;
        if(cVar1S4S66P015N044P003P055(0)='1' AND  B( 1)='0' )then
          cVar2S4S66P035nsss(0) <='1';
          else
          cVar2S4S66P035nsss(0) <='0';
          end if;
        if(cVar1S5S66P015N044P003N055(0)='1' AND  A( 6)='0' AND A( 7)='1' )then
          cVar2S5S66P007P005nsss(0) <='1';
          else
          cVar2S5S66P007P005nsss(0) <='0';
          end if;
        if(cVar1S6S66P015N044P003N055(0)='1' AND  A( 6)='0' AND A( 7)='0' AND A( 4)='0' )then
          cVar2S6S66P007N005P011nsss(0) <='1';
          else
          cVar2S6S66P007N005P011nsss(0) <='0';
          end if;
        if(cVar1S7S66P015N044P003N055(0)='1' AND  A( 6)='1' AND A( 3)='0' AND D( 0)='1' )then
          cVar2S7S66P007P013P066nsss(0) <='1';
          else
          cVar2S7S66P007P013P066nsss(0) <='0';
          end if;
        if(cVar1S8S66P015N044N003P027(0)='1' AND  B(14)='0' AND B( 6)='0' )then
          cVar2S8S66P026P025nsss(0) <='1';
          else
          cVar2S8S66P026P025nsss(0) <='0';
          end if;
        if(cVar1S9S66P015N044N003N027(0)='1' AND  D(15)='0' AND E( 5)='0' AND A(16)='0' )then
          cVar2S9S66P039P048P006nsss(0) <='1';
          else
          cVar2S9S66P039P048P006nsss(0) <='0';
          end if;
        if(cVar1S10S66P015N044N003N027(0)='1' AND  D(15)='0' AND E( 5)='1' AND E(10)='1' )then
          cVar2S10S66P039P048P061nsss(0) <='1';
          else
          cVar2S10S66P039P048P061nsss(0) <='0';
          end if;
        if(cVar1S11S66P015N044N003N027(0)='1' AND  D(15)='1' AND D( 8)='1' )then
          cVar2S11S66P039P067nsss(0) <='1';
          else
          cVar2S11S66P039P067nsss(0) <='0';
          end if;
        if(cVar1S12S66N015P063P037P067(0)='1' AND  B(11)='1' AND A( 0)='1' )then
          cVar2S12S66P032P019nsss(0) <='1';
          else
          cVar2S12S66P032P019nsss(0) <='0';
          end if;
        if(cVar1S13S66N015P063P037P067(0)='1' AND  B(11)='1' AND A( 0)='0' AND A(12)='1' )then
          cVar2S13S66P032N019P014nsss(0) <='1';
          else
          cVar2S13S66P032N019P014nsss(0) <='0';
          end if;
        if(cVar1S14S66N015P063P037P067(0)='1' AND  B(11)='0' )then
          cVar2S14S66N032psss(0) <='1';
          else
          cVar2S14S66N032psss(0) <='0';
          end if;
        if(cVar1S15S66N015P063P037P067(0)='1' AND  A( 4)='1' AND D( 0)='1' )then
          cVar2S15S66P011P066nsss(0) <='1';
          else
          cVar2S15S66P011P066nsss(0) <='0';
          end if;
        if(cVar1S16S66N015P063P037P067(0)='1' AND  A( 4)='0' AND A(10)='1' AND B( 1)='0' )then
          cVar2S16S66N011P018P035nsss(0) <='1';
          else
          cVar2S16S66N011P018P035nsss(0) <='0';
          end if;
        if(cVar1S17S66N015P063N037P017(0)='1' AND  E( 4)='0' AND D(10)='0' AND A( 0)='0' )then
          cVar2S17S66P052P059P019nsss(0) <='1';
          else
          cVar2S17S66P052P059P019nsss(0) <='0';
          end if;
        if(cVar1S18S66N015P063N037P017(0)='1' AND  E( 4)='0' AND D(10)='1' AND A( 0)='1' )then
          cVar2S18S66P052P059P019nsss(0) <='1';
          else
          cVar2S18S66P052P059P019nsss(0) <='0';
          end if;
        if(cVar1S19S66N015P063N037P017(0)='1' AND  E( 4)='1' AND B( 4)='0' AND D( 4)='1' )then
          cVar2S19S66P052P029P050nsss(0) <='1';
          else
          cVar2S19S66P052P029P050nsss(0) <='0';
          end if;
        if(cVar1S20S66N015P063N037N017(0)='1' AND  E( 0)='1' AND A(10)='0' )then
          cVar2S20S66P068P018nsss(0) <='1';
          else
          cVar2S20S66P068P018nsss(0) <='0';
          end if;
        if(cVar1S21S66N015P063N037N017(0)='1' AND  E( 0)='1' AND A(10)='1' AND A( 3)='1' )then
          cVar2S21S66P068P018P013nsss(0) <='1';
          else
          cVar2S21S66P068P018P013nsss(0) <='0';
          end if;
        if(cVar1S22S66N015P063N037N017(0)='1' AND  E( 0)='0' AND B( 9)='1' AND E(12)='1' )then
          cVar2S22S66N068P036P053nsss(0) <='1';
          else
          cVar2S22S66N068P036P053nsss(0) <='0';
          end if;
        if(cVar1S23S66N015N063P029P058(0)='1' AND  B( 9)='0' AND B( 0)='0' AND D(11)='0' )then
          cVar2S23S66P036P037P055nsss(0) <='1';
          else
          cVar2S23S66P036P037P055nsss(0) <='0';
          end if;
        if(cVar1S24S66N015N063P029P058(0)='1' AND  B( 9)='0' AND B( 0)='1' AND A( 5)='0' )then
          cVar2S24S66P036P037P009nsss(0) <='1';
          else
          cVar2S24S66P036P037P009nsss(0) <='0';
          end if;
        if(cVar1S25S66N015N063P029P058(0)='1' AND  B( 9)='1' AND A( 4)='1' )then
          cVar2S25S66P036P011nsss(0) <='1';
          else
          cVar2S25S66P036P011nsss(0) <='0';
          end if;
        if(cVar1S26S66N015N063P029P058(0)='1' AND  B( 9)='1' AND A( 4)='0' AND A( 5)='1' )then
          cVar2S26S66P036N011P009nsss(0) <='1';
          else
          cVar2S26S66P036N011P009nsss(0) <='0';
          end if;
        if(cVar1S27S66N015N063P029P058(0)='1' AND  A( 1)='0' AND D(12)='0' AND B( 2)='1' )then
          cVar2S27S66P017P051P033nsss(0) <='1';
          else
          cVar2S27S66P017P051P033nsss(0) <='0';
          end if;
        if(cVar1S28S66N015N063N029P028(0)='1' AND  D(14)='1' )then
          cVar2S28S66P043nsss(0) <='1';
          else
          cVar2S28S66P043nsss(0) <='0';
          end if;
        if(cVar1S29S66N015N063N029P028(0)='1' AND  D(14)='0' AND D(15)='0' )then
          cVar2S29S66N043P039nsss(0) <='1';
          else
          cVar2S29S66N043P039nsss(0) <='0';
          end if;
        if(cVar1S30S66N015N063N029N028(0)='1' AND  D( 4)='0' AND A( 4)='0' AND A(12)='1' )then
          cVar2S30S66P050P011P014nsss(0) <='1';
          else
          cVar2S30S66P050P011P014nsss(0) <='0';
          end if;
        if(cVar1S31S66N015N063N029N028(0)='1' AND  D( 4)='0' AND A( 4)='1' AND B( 3)='1' )then
          cVar2S31S66P050P011P031nsss(0) <='1';
          else
          cVar2S31S66P050P011P031nsss(0) <='0';
          end if;
        if(cVar1S32S66N015N063N029N028(0)='1' AND  D( 4)='1' AND B( 5)='1' AND A( 1)='1' )then
          cVar2S32S66P050P027P017nsss(0) <='1';
          else
          cVar2S32S66P050P027P017nsss(0) <='0';
          end if;
        if(cVar1S33S66N015N063N029N028(0)='1' AND  D( 4)='1' AND B( 5)='0' AND B(14)='1' )then
          cVar2S33S66P050N027P026nsss(0) <='1';
          else
          cVar2S33S66P050N027P026nsss(0) <='0';
          end if;
        if(cVar1S0S67P015P014P050P061(0)='1' AND  B(13)='0' AND B(10)='0' )then
          cVar2S0S67P028P034nsss(0) <='1';
          else
          cVar2S0S67P028P034nsss(0) <='0';
          end if;
        if(cVar1S1S67P015P014P050P061(0)='1' AND  B(13)='0' AND B(10)='1' AND E( 8)='0' )then
          cVar2S1S67P028P034P069nsss(0) <='1';
          else
          cVar2S1S67P028P034P069nsss(0) <='0';
          end if;
        if(cVar1S2S67P015P014P050P061(0)='1' AND  B(13)='1' AND A(10)='0' )then
          cVar2S2S67P028P018nsss(0) <='1';
          else
          cVar2S2S67P028P018nsss(0) <='0';
          end if;
        if(cVar1S3S67P015P014P050P061(0)='1' AND  B(13)='1' AND A(10)='1' AND B( 1)='1' )then
          cVar2S3S67P028P018P035nsss(0) <='1';
          else
          cVar2S3S67P028P018P035nsss(0) <='0';
          end if;
        if(cVar1S4S67P015P014P050P061(0)='1' AND  B( 1)='1' AND A( 5)='0' AND A(14)='0' )then
          cVar2S4S67P035P009P010nsss(0) <='1';
          else
          cVar2S4S67P035P009P010nsss(0) <='0';
          end if;
        if(cVar1S5S67P015P014P050P061(0)='1' AND  B( 1)='0' AND B(17)='1' )then
          cVar2S5S67N035P020nsss(0) <='1';
          else
          cVar2S5S67N035P020nsss(0) <='0';
          end if;
        if(cVar1S6S67P015P014P050P061(0)='1' AND  B( 1)='0' AND B(17)='0' AND B( 3)='1' )then
          cVar2S6S67N035N020P031nsss(0) <='1';
          else
          cVar2S6S67N035N020P031nsss(0) <='0';
          end if;
        if(cVar1S7S67P015P014P050P011(0)='1' AND  B( 1)='0' AND A(13)='1' )then
          cVar2S7S67P035P012nsss(0) <='1';
          else
          cVar2S7S67P035P012nsss(0) <='0';
          end if;
        if(cVar1S8S67P015P014P050P011(0)='1' AND  B( 1)='0' AND A(13)='0' AND D( 3)='0' )then
          cVar2S8S67P035N012P054nsss(0) <='1';
          else
          cVar2S8S67P035N012P054nsss(0) <='0';
          end if;
        if(cVar1S9S67P015P014P050N011(0)='1' AND  A(14)='1' AND A( 0)='1' )then
          cVar2S9S67P010P019nsss(0) <='1';
          else
          cVar2S9S67P010P019nsss(0) <='0';
          end if;
        if(cVar1S10S67P015P014P050N011(0)='1' AND  A(14)='1' AND A( 0)='0' AND D( 3)='0' )then
          cVar2S10S67P010N019P054nsss(0) <='1';
          else
          cVar2S10S67P010N019P054nsss(0) <='0';
          end if;
        if(cVar1S11S67P015P014P050N011(0)='1' AND  A(14)='0' AND B( 5)='1' AND A( 6)='1' )then
          cVar2S11S67N010P027P007nsss(0) <='1';
          else
          cVar2S11S67N010P027P007nsss(0) <='0';
          end if;
        if(cVar1S12S67P015P014P021P012(0)='1' AND  B( 2)='1' AND A( 0)='0' AND D(12)='0' )then
          cVar2S12S67P033P019P051nsss(0) <='1';
          else
          cVar2S12S67P033P019P051nsss(0) <='0';
          end if;
        if(cVar1S13S67P015P014P021P012(0)='1' AND  B( 2)='1' AND A( 0)='1' AND E( 3)='1' )then
          cVar2S13S67P033P019P056nsss(0) <='1';
          else
          cVar2S13S67P033P019P056nsss(0) <='0';
          end if;
        if(cVar1S14S67P015P014P021P012(0)='1' AND  B( 2)='0' AND E(11)='1' )then
          cVar2S14S67N033P057nsss(0) <='1';
          else
          cVar2S14S67N033P057nsss(0) <='0';
          end if;
        if(cVar1S15S67P015P014P021P012(0)='1' AND  B( 2)='0' AND E(11)='0' AND D( 4)='1' )then
          cVar2S15S67N033N057P050nsss(0) <='1';
          else
          cVar2S15S67N033N057P050nsss(0) <='0';
          end if;
        if(cVar1S16S67P015P014P021P012(0)='1' AND  A( 5)='0' AND E( 0)='1' )then
          cVar2S16S67P009P068nsss(0) <='1';
          else
          cVar2S16S67P009P068nsss(0) <='0';
          end if;
        if(cVar1S17S67P015P014P021P012(0)='1' AND  A( 5)='0' AND E( 0)='0' AND D( 1)='1' )then
          cVar2S17S67P009N068P062nsss(0) <='1';
          else
          cVar2S17S67P009N068P062nsss(0) <='0';
          end if;
        if(cVar1S18S67P015P014P021P012(0)='1' AND  A(14)='0' AND B(11)='1' )then
          cVar2S18S67P010P032nsss(0) <='1';
          else
          cVar2S18S67P010P032nsss(0) <='0';
          end if;
        if(cVar1S19S67P015P014P021P012(0)='1' AND  A(14)='0' AND B(11)='0' AND A(15)='1' )then
          cVar2S19S67P010N032P008nsss(0) <='1';
          else
          cVar2S19S67P010N032P008nsss(0) <='0';
          end if;
        if(cVar1S21S67P015P044P031N006(0)='1' AND  E( 0)='1' )then
          cVar2S21S67P068nsss(0) <='1';
          else
          cVar2S21S67P068nsss(0) <='0';
          end if;
        if(cVar1S22S67P015P044P031N006(0)='1' AND  E( 0)='0' AND A(17)='1' )then
          cVar2S22S67N068P004nsss(0) <='1';
          else
          cVar2S22S67N068P004nsss(0) <='0';
          end if;
        if(cVar1S24S67P015N044P003N055(0)='1' AND  A( 6)='0' AND A( 7)='1' )then
          cVar2S24S67P007P005nsss(0) <='1';
          else
          cVar2S24S67P007P005nsss(0) <='0';
          end if;
        if(cVar1S25S67P015N044P003N055(0)='1' AND  A( 6)='0' AND A( 7)='0' AND E( 0)='1' )then
          cVar2S25S67P007N005P068nsss(0) <='1';
          else
          cVar2S25S67P007N005P068nsss(0) <='0';
          end if;
        if(cVar1S26S67P015N044P003N055(0)='1' AND  A( 6)='1' AND A( 3)='0' AND D( 0)='1' )then
          cVar2S26S67P007P013P066nsss(0) <='1';
          else
          cVar2S26S67P007P013P066nsss(0) <='0';
          end if;
        if(cVar1S27S67P015N044N003P027(0)='1' AND  B(14)='0' AND B( 6)='0' )then
          cVar2S27S67P026P025nsss(0) <='1';
          else
          cVar2S27S67P026P025nsss(0) <='0';
          end if;
        if(cVar1S28S67P015N044N003P027(0)='1' AND  B(14)='1' AND A( 0)='1' )then
          cVar2S28S67P026P019nsss(0) <='1';
          else
          cVar2S28S67P026P019nsss(0) <='0';
          end if;
        if(cVar1S29S67P015N044N003N027(0)='1' AND  D(15)='0' AND B( 7)='0' AND A(10)='1' )then
          cVar2S29S67P039P023P018nsss(0) <='1';
          else
          cVar2S29S67P039P023P018nsss(0) <='0';
          end if;
        if(cVar1S30S67P015N044N003N027(0)='1' AND  D(15)='0' AND B( 7)='1' AND A(12)='1' )then
          cVar2S30S67P039P023P014nsss(0) <='1';
          else
          cVar2S30S67P039P023P014nsss(0) <='0';
          end if;
        if(cVar1S31S67P015N044N003N027(0)='1' AND  D(15)='1' AND D( 8)='1' )then
          cVar2S31S67P039P067nsss(0) <='1';
          else
          cVar2S31S67P039P067nsss(0) <='0';
          end if;
        if(cVar1S0S68P014P012P021P032(0)='1' AND  D( 1)='0' AND D(12)='0' )then
          cVar2S0S68P062P051nsss(0) <='1';
          else
          cVar2S0S68P062P051nsss(0) <='0';
          end if;
        if(cVar1S1S68P014P012P021P032(0)='1' AND  D( 1)='1' AND A( 0)='1' )then
          cVar2S1S68P062P019nsss(0) <='1';
          else
          cVar2S1S68P062P019nsss(0) <='0';
          end if;
        if(cVar1S2S68P014P012P021P032(0)='1' AND  D( 1)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar2S2S68P062N019P066nsss(0) <='1';
          else
          cVar2S2S68P062N019P066nsss(0) <='0';
          end if;
        if(cVar1S3S68P014P012P021N032(0)='1' AND  A(10)='0' AND E( 2)='1' )then
          cVar2S3S68P018P060nsss(0) <='1';
          else
          cVar2S3S68P018P060nsss(0) <='0';
          end if;
        if(cVar1S4S68P014P012P021N032(0)='1' AND  A(10)='0' AND E( 2)='0' AND A( 5)='0' )then
          cVar2S4S68P018N060P009nsss(0) <='1';
          else
          cVar2S4S68P018N060P009nsss(0) <='0';
          end if;
        if(cVar1S5S68P014P012P021N032(0)='1' AND  A(10)='1' AND B( 7)='1' AND A( 3)='0' )then
          cVar2S5S68P018P023P013nsss(0) <='1';
          else
          cVar2S5S68P018P023P013nsss(0) <='0';
          end if;
        if(cVar1S6S68P014P012P021N032(0)='1' AND  A(10)='1' AND B( 7)='0' AND A( 0)='0' )then
          cVar2S6S68P018N023P019nsss(0) <='1';
          else
          cVar2S6S68P018N023P019nsss(0) <='0';
          end if;
        if(cVar1S7S68P014P012P021P026(0)='1' AND  D( 0)='1' AND A( 1)='0' )then
          cVar2S7S68P066P017nsss(0) <='1';
          else
          cVar2S7S68P066P017nsss(0) <='0';
          end if;
        if(cVar1S9S68P014P012P001N010(0)='1' AND  B(10)='1' )then
          cVar2S9S68P034nsss(0) <='1';
          else
          cVar2S9S68P034nsss(0) <='0';
          end if;
        if(cVar1S10S68P014P012P001N010(0)='1' AND  B(10)='0' AND A( 5)='1' )then
          cVar2S10S68N034P009nsss(0) <='1';
          else
          cVar2S10S68N034P009nsss(0) <='0';
          end if;
        if(cVar1S11S68P014P012N001P009(0)='1' AND  D(12)='0' AND D( 0)='1' )then
          cVar2S11S68P051P066nsss(0) <='1';
          else
          cVar2S11S68P051P066nsss(0) <='0';
          end if;
        if(cVar1S12S68P014P012N001P009(0)='1' AND  D(12)='0' AND D( 0)='0' AND E( 3)='1' )then
          cVar2S12S68P051N066P056nsss(0) <='1';
          else
          cVar2S12S68P051N066P056nsss(0) <='0';
          end if;
        if(cVar1S13S68P014P012N001P009(0)='1' AND  D(12)='1' AND D( 0)='0' AND A(10)='1' )then
          cVar2S13S68P051P066P018nsss(0) <='1';
          else
          cVar2S13S68P051P066P018nsss(0) <='0';
          end if;
        if(cVar1S14S68P014P012N001P009(0)='1' AND  A(17)='1' AND A( 4)='0' )then
          cVar2S14S68P004P011nsss(0) <='1';
          else
          cVar2S14S68P004P011nsss(0) <='0';
          end if;
        if(cVar1S15S68N014P027P009P063(0)='1' AND  D( 8)='1' AND E(13)='1' )then
          cVar2S15S68P067P049nsss(0) <='1';
          else
          cVar2S15S68P067P049nsss(0) <='0';
          end if;
        if(cVar1S16S68N014P027P009P063(0)='1' AND  D( 8)='1' AND E(13)='0' AND A(10)='0' )then
          cVar2S16S68P067N049P018nsss(0) <='1';
          else
          cVar2S16S68P067N049P018nsss(0) <='0';
          end if;
        if(cVar1S17S68N014P027P009P063(0)='1' AND  D( 8)='0' )then
          cVar2S17S68N067psss(0) <='1';
          else
          cVar2S17S68N067psss(0) <='0';
          end if;
        if(cVar1S18S68N014P027P009P063(0)='1' AND  B(10)='0' )then
          cVar2S18S68P034nsss(0) <='1';
          else
          cVar2S18S68P034nsss(0) <='0';
          end if;
        if(cVar1S19S68N014P027N009P026(0)='1' AND  B( 7)='0' AND A( 7)='1' )then
          cVar2S19S68P023P005nsss(0) <='1';
          else
          cVar2S19S68P023P005nsss(0) <='0';
          end if;
        if(cVar1S20S68N014P027N009P026(0)='1' AND  B( 7)='0' AND A( 7)='0' AND A(15)='1' )then
          cVar2S20S68P023N005P008nsss(0) <='1';
          else
          cVar2S20S68P023N005P008nsss(0) <='0';
          end if;
        if(cVar1S21S68N014P027N009P026(0)='1' AND  A(14)='0' AND A( 2)='0' AND E( 0)='1' )then
          cVar2S21S68P010P015P068nsss(0) <='1';
          else
          cVar2S21S68P010P015P068nsss(0) <='0';
          end if;
        if(cVar1S22S68N014N027P017P069(0)='1' AND  A( 9)='1' AND E( 0)='1' )then
          cVar2S22S68P001P068nsss(0) <='1';
          else
          cVar2S22S68P001P068nsss(0) <='0';
          end if;
        if(cVar1S23S68N014N027P017P069(0)='1' AND  A( 9)='1' AND E( 0)='0' AND A( 0)='1' )then
          cVar2S23S68P001N068P019nsss(0) <='1';
          else
          cVar2S23S68P001N068P019nsss(0) <='0';
          end if;
        if(cVar1S24S68N014N027P017P069(0)='1' AND  A( 9)='0' AND D( 0)='0' AND A( 3)='0' )then
          cVar2S24S68N001P066P013nsss(0) <='1';
          else
          cVar2S24S68N001P066P013nsss(0) <='0';
          end if;
        if(cVar1S25S68N014N027P017P069(0)='1' AND  A( 9)='0' AND D( 0)='1' AND E( 1)='1' )then
          cVar2S25S68N001P066P064nsss(0) <='1';
          else
          cVar2S25S68N001P066P064nsss(0) <='0';
          end if;
        if(cVar1S26S68N014N027P017N069(0)='1' AND  D( 1)='0' AND D( 8)='0' AND A(10)='0' )then
          cVar2S26S68P062P067P018nsss(0) <='1';
          else
          cVar2S26S68P062P067P018nsss(0) <='0';
          end if;
        if(cVar1S27S68N014N027P017N069(0)='1' AND  D( 1)='1' AND A( 2)='1' AND A( 3)='0' )then
          cVar2S27S68P062P015P013nsss(0) <='1';
          else
          cVar2S27S68P062P015P013nsss(0) <='0';
          end if;
        if(cVar1S28S68N014N027P017N069(0)='1' AND  D( 1)='1' AND A( 2)='0' AND A( 3)='1' )then
          cVar2S28S68P062N015P013nsss(0) <='1';
          else
          cVar2S28S68P062N015P013nsss(0) <='0';
          end if;
        if(cVar1S29S68N014N027P017P061(0)='1' AND  A( 7)='0' AND D( 6)='0' AND A(16)='0' )then
          cVar2S29S68P005P042P006nsss(0) <='1';
          else
          cVar2S29S68P005P042P006nsss(0) <='0';
          end if;
        if(cVar1S30S68N014N027P017P061(0)='1' AND  A( 7)='1' AND A(10)='0' )then
          cVar2S30S68P005P018nsss(0) <='1';
          else
          cVar2S30S68P005P018nsss(0) <='0';
          end if;
        if(cVar1S31S68N014N027P017N061(0)='1' AND  E( 6)='1' AND B( 2)='0' )then
          cVar2S31S68P044P033nsss(0) <='1';
          else
          cVar2S31S68P044P033nsss(0) <='0';
          end if;
        if(cVar1S32S68N014N027P017N061(0)='1' AND  E( 6)='0' AND B( 7)='0' AND E(14)='1' )then
          cVar2S32S68N044P023P045nsss(0) <='1';
          else
          cVar2S32S68N044P023P045nsss(0) <='0';
          end if;
        if(cVar1S33S68N014N027P017N061(0)='1' AND  E( 6)='0' AND B( 7)='1' AND E( 9)='1' )then
          cVar2S33S68N044P023P065nsss(0) <='1';
          else
          cVar2S33S68N044P023P065nsss(0) <='0';
          end if;
        if(cVar1S0S69P017P062P034P064(0)='1' AND  D( 9)='0' AND E( 9)='1' )then
          cVar2S0S69P063P065nsss(0) <='1';
          else
          cVar2S0S69P063P065nsss(0) <='0';
          end if;
        if(cVar1S1S69P017P062P034P064(0)='1' AND  D( 9)='0' AND E( 9)='0' AND D(11)='0' )then
          cVar2S1S69P063N065P055nsss(0) <='1';
          else
          cVar2S1S69P063N065P055nsss(0) <='0';
          end if;
        if(cVar1S2S69P017P062P034P064(0)='1' AND  D( 9)='1' AND A( 7)='1' )then
          cVar2S2S69P063P005nsss(0) <='1';
          else
          cVar2S2S69P063P005nsss(0) <='0';
          end if;
        if(cVar1S3S69P017P062P034P064(0)='1' AND  D( 9)='1' AND A( 7)='0' AND E( 5)='0' )then
          cVar2S3S69P063N005P048nsss(0) <='1';
          else
          cVar2S3S69P063N005P048nsss(0) <='0';
          end if;
        if(cVar1S4S69P017P062P034N064(0)='1' AND  E( 9)='1' AND A( 0)='0' AND D( 8)='0' )then
          cVar2S4S69P065P019P067nsss(0) <='1';
          else
          cVar2S4S69P065P019P067nsss(0) <='0';
          end if;
        if(cVar1S5S69P017P062P034N064(0)='1' AND  E( 9)='0' AND B( 1)='1' AND B(11)='0' )then
          cVar2S5S69N065P035P032nsss(0) <='1';
          else
          cVar2S5S69N065P035P032nsss(0) <='0';
          end if;
        if(cVar1S6S69P017P062P034N064(0)='1' AND  E( 9)='0' AND B( 1)='0' AND B(12)='1' )then
          cVar2S6S69N065N035P030nsss(0) <='1';
          else
          cVar2S6S69N065N035P030nsss(0) <='0';
          end if;
        if(cVar1S7S69P017P062P034P060(0)='1' AND  D(10)='1' )then
          cVar2S7S69P059nsss(0) <='1';
          else
          cVar2S7S69P059nsss(0) <='0';
          end if;
        if(cVar1S8S69P017P062P034P060(0)='1' AND  D(10)='0' AND A( 2)='0' )then
          cVar2S8S69N059P015nsss(0) <='1';
          else
          cVar2S8S69N059P015nsss(0) <='0';
          end if;
        if(cVar1S9S69P017P062P034N060(0)='1' AND  A( 5)='1' AND A(12)='0' )then
          cVar2S9S69P009P014nsss(0) <='1';
          else
          cVar2S9S69P009P014nsss(0) <='0';
          end if;
        if(cVar1S10S69P017P062P034N060(0)='1' AND  A( 5)='1' AND A(12)='1' AND A(11)='1' )then
          cVar2S10S69P009P014P016nsss(0) <='1';
          else
          cVar2S10S69P009P014P016nsss(0) <='0';
          end if;
        if(cVar1S11S69P017P062P034N060(0)='1' AND  A( 5)='0' AND B( 9)='1' AND E( 8)='0' )then
          cVar2S11S69N009P036P069nsss(0) <='1';
          else
          cVar2S11S69N009P036P069nsss(0) <='0';
          end if;
        if(cVar1S12S69P017P062P034N060(0)='1' AND  A( 5)='0' AND B( 9)='0' AND E( 8)='1' )then
          cVar2S12S69N009N036P069nsss(0) <='1';
          else
          cVar2S12S69N009N036P069nsss(0) <='0';
          end if;
        if(cVar1S13S69P017N062P014P054(0)='1' AND  A(13)='1' AND B( 3)='1' )then
          cVar2S13S69P012P031nsss(0) <='1';
          else
          cVar2S13S69P012P031nsss(0) <='0';
          end if;
        if(cVar1S14S69P017N062P014P054(0)='1' AND  A(13)='1' AND B( 3)='0' AND B( 4)='1' )then
          cVar2S14S69P012N031P029nsss(0) <='1';
          else
          cVar2S14S69P012N031P029nsss(0) <='0';
          end if;
        if(cVar1S15S69P017N062P014P054(0)='1' AND  A(13)='0' AND B(14)='0' AND B( 4)='1' )then
          cVar2S15S69N012P026P029nsss(0) <='1';
          else
          cVar2S15S69N012P026P029nsss(0) <='0';
          end if;
        if(cVar1S16S69P017N062P014N054(0)='1' AND  E( 7)='1' AND A(18)='1' )then
          cVar2S16S69P040P002nsss(0) <='1';
          else
          cVar2S16S69P040P002nsss(0) <='0';
          end if;
        if(cVar1S17S69P017N062P014N054(0)='1' AND  E( 7)='1' AND A(18)='0' AND E( 8)='1' )then
          cVar2S17S69P040N002P069nsss(0) <='1';
          else
          cVar2S17S69P040N002P069nsss(0) <='0';
          end if;
        if(cVar1S18S69P017N062P014N054(0)='1' AND  E( 7)='0' AND D( 7)='0' AND D(13)='1' )then
          cVar2S18S69N040P038P047nsss(0) <='1';
          else
          cVar2S18S69N040P038P047nsss(0) <='0';
          end if;
        if(cVar1S19S69P017N062P014P035(0)='1' AND  B( 6)='1' AND E( 0)='1' )then
          cVar2S19S69P025P068nsss(0) <='1';
          else
          cVar2S19S69P025P068nsss(0) <='0';
          end if;
        if(cVar1S20S69P017N062P014P035(0)='1' AND  B( 6)='1' AND E( 0)='0' AND A(10)='0' )then
          cVar2S20S69P025N068P018nsss(0) <='1';
          else
          cVar2S20S69P025N068P018nsss(0) <='0';
          end if;
        if(cVar1S21S69P017N062P014P035(0)='1' AND  B( 6)='0' AND D(15)='0' AND D( 2)='1' )then
          cVar2S21S69N025P039P058nsss(0) <='1';
          else
          cVar2S21S69N025P039P058nsss(0) <='0';
          end if;
        if(cVar1S22S69P017N062P014P035(0)='1' AND  E( 0)='0' AND D( 0)='0' AND A( 6)='0' )then
          cVar2S22S69P068P066P007nsss(0) <='1';
          else
          cVar2S22S69P068P066P007nsss(0) <='0';
          end if;
        if(cVar1S23S69P017N062P014P035(0)='1' AND  E( 0)='1' AND A(11)='0' AND A( 2)='1' )then
          cVar2S23S69P068P016P015nsss(0) <='1';
          else
          cVar2S23S69P068P016P015nsss(0) <='0';
          end if;
        if(cVar1S24S69N017P066P028P055(0)='1' AND  D(12)='1' AND E( 1)='0' )then
          cVar2S24S69P051P064nsss(0) <='1';
          else
          cVar2S24S69P051P064nsss(0) <='0';
          end if;
        if(cVar1S25S69N017P066P028P055(0)='1' AND  D(12)='1' AND E( 1)='1' AND E( 0)='0' )then
          cVar2S25S69P051P064P068nsss(0) <='1';
          else
          cVar2S25S69P051P064P068nsss(0) <='0';
          end if;
        if(cVar1S26S69N017P066P028P055(0)='1' AND  D(12)='0' AND B(14)='0' )then
          cVar2S26S69N051P026nsss(0) <='1';
          else
          cVar2S26S69N051P026nsss(0) <='0';
          end if;
        if(cVar1S27S69N017P066P028P055(0)='1' AND  B(12)='1' AND A( 3)='1' AND A(10)='1' )then
          cVar2S27S69P030P013P018nsss(0) <='1';
          else
          cVar2S27S69P030P013P018nsss(0) <='0';
          end if;
        if(cVar1S28S69N017P066P028P055(0)='1' AND  B(12)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar2S28S69P030N013P011nsss(0) <='1';
          else
          cVar2S28S69P030N013P011nsss(0) <='0';
          end if;
        if(cVar1S29S69N017P066P028P055(0)='1' AND  B(12)='0' AND B(11)='1' )then
          cVar2S29S69N030P032nsss(0) <='1';
          else
          cVar2S29S69N030P032nsss(0) <='0';
          end if;
        if(cVar1S30S69N017P066P028P055(0)='1' AND  B(12)='0' AND B(11)='0' AND A( 6)='1' )then
          cVar2S30S69N030N032P007nsss(0) <='1';
          else
          cVar2S30S69N030N032P007nsss(0) <='0';
          end if;
        if(cVar1S31S69N017P066P028P030(0)='1' AND  E( 0)='1' AND D(12)='0' AND D(11)='1' )then
          cVar2S31S69P068P051P055nsss(0) <='1';
          else
          cVar2S31S69P068P051P055nsss(0) <='0';
          end if;
        if(cVar1S32S69N017N066P047P049(0)='1' AND  D(12)='0' AND B(14)='1' )then
          cVar2S32S69P051P026nsss(0) <='1';
          else
          cVar2S32S69P051P026nsss(0) <='0';
          end if;
        if(cVar1S33S69N017N066P047P049(0)='1' AND  D(12)='0' AND B(14)='0' AND A(10)='1' )then
          cVar2S33S69P051N026P018nsss(0) <='1';
          else
          cVar2S33S69P051N026P018nsss(0) <='0';
          end if;
        if(cVar1S34S69N017N066P047P049(0)='1' AND  D(12)='1' AND A(15)='1' )then
          cVar2S34S69P051P008nsss(0) <='1';
          else
          cVar2S34S69P051P008nsss(0) <='0';
          end if;
        if(cVar1S35S69N017N066P047N049(0)='1' AND  B(15)='1' AND E(14)='1' )then
          cVar2S35S69P024P045nsss(0) <='1';
          else
          cVar2S35S69P024P045nsss(0) <='0';
          end if;
        if(cVar1S36S69N017N066P047N049(0)='1' AND  B(15)='0' AND B( 6)='1' )then
          cVar2S36S69N024P025nsss(0) <='1';
          else
          cVar2S36S69N024P025nsss(0) <='0';
          end if;
        if(cVar1S37S69N017N066P047N049(0)='1' AND  B(15)='0' AND B( 6)='0' AND D(12)='1' )then
          cVar2S37S69N024N025P051nsss(0) <='1';
          else
          cVar2S37S69N024N025P051nsss(0) <='0';
          end if;
        if(cVar1S38S69N017N066N047P023(0)='1' AND  A(11)='1' )then
          cVar2S38S69P016nsss(0) <='1';
          else
          cVar2S38S69P016nsss(0) <='0';
          end if;
        if(cVar1S39S69N017N066N047P023(0)='1' AND  A(11)='0' AND E( 2)='0' )then
          cVar2S39S69N016P060nsss(0) <='1';
          else
          cVar2S39S69N016P060nsss(0) <='0';
          end if;
        if(cVar1S40S69N017N066N047N023(0)='1' AND  D( 6)='0' AND D( 8)='1' AND B(12)='1' )then
          cVar2S40S69P042P067P030nsss(0) <='1';
          else
          cVar2S40S69P042P067P030nsss(0) <='0';
          end if;
        if(cVar1S41S69N017N066N047N023(0)='1' AND  D( 6)='0' AND D( 8)='0' AND D( 5)='1' )then
          cVar2S41S69P042N067P046nsss(0) <='1';
          else
          cVar2S41S69P042N067P046nsss(0) <='0';
          end if;
        if(cVar1S42S69N017N066N047N023(0)='1' AND  D( 6)='1' AND B( 8)='1' AND E( 7)='0' )then
          cVar2S42S69P042P021P040nsss(0) <='1';
          else
          cVar2S42S69P042P021P040nsss(0) <='0';
          end if;
        if(cVar1S43S69N017N066N047N023(0)='1' AND  D( 6)='1' AND B( 8)='0' AND A(16)='1' )then
          cVar2S43S69P042N021P006nsss(0) <='1';
          else
          cVar2S43S69P042N021P006nsss(0) <='0';
          end if;
        if(cVar1S0S70P017P014P062P010(0)='1' AND  B(17)='0' AND D(13)='1' )then
          cVar2S0S70P020P047nsss(0) <='1';
          else
          cVar2S0S70P020P047nsss(0) <='0';
          end if;
        if(cVar1S1S70P017P014P062P010(0)='1' AND  B(17)='0' AND D(13)='0' AND A(13)='0' )then
          cVar2S1S70P020N047P012nsss(0) <='1';
          else
          cVar2S1S70P020N047P012nsss(0) <='0';
          end if;
        if(cVar1S2S70P017P014P062N010(0)='1' AND  D(13)='0' AND A( 6)='0' )then
          cVar2S2S70P047P007nsss(0) <='1';
          else
          cVar2S2S70P047P007nsss(0) <='0';
          end if;
        if(cVar1S3S70P017P014P062N010(0)='1' AND  D(13)='1' AND A(16)='1' )then
          cVar2S3S70P047P006nsss(0) <='1';
          else
          cVar2S3S70P047P006nsss(0) <='0';
          end if;
        if(cVar1S4S70P017P014P062N010(0)='1' AND  D(13)='1' AND A(16)='0' AND A( 5)='1' )then
          cVar2S4S70P047N006P009nsss(0) <='1';
          else
          cVar2S4S70P047N006P009nsss(0) <='0';
          end if;
        if(cVar1S5S70P017P014P062P033(0)='1' AND  A(14)='0' )then
          cVar2S5S70P010nsss(0) <='1';
          else
          cVar2S5S70P010nsss(0) <='0';
          end if;
        if(cVar1S6S70P017P014P062N033(0)='1' AND  B( 7)='0' AND E( 7)='1' AND D( 7)='0' )then
          cVar2S6S70P023P040P038nsss(0) <='1';
          else
          cVar2S6S70P023P040P038nsss(0) <='0';
          end if;
        if(cVar1S7S70P017P014P062N033(0)='1' AND  B( 7)='0' AND E( 7)='0' AND A(11)='1' )then
          cVar2S7S70P023N040P016nsss(0) <='1';
          else
          cVar2S7S70P023N040P016nsss(0) <='0';
          end if;
        if(cVar1S9S70P017P014P012N041(0)='1' AND  D(15)='0' AND E( 8)='1' AND D( 1)='1' )then
          cVar2S9S70P039P069P062nsss(0) <='1';
          else
          cVar2S9S70P039P069P062nsss(0) <='0';
          end if;
        if(cVar1S10S70P017P014P012P049(0)='1' AND  A( 9)='1' )then
          cVar2S10S70P001nsss(0) <='1';
          else
          cVar2S10S70P001nsss(0) <='0';
          end if;
        if(cVar1S11S70P017P014P012P049(0)='1' AND  A( 9)='0' AND A(10)='1' AND A(14)='0' )then
          cVar2S11S70N001P018P010nsss(0) <='1';
          else
          cVar2S11S70N001P018P010nsss(0) <='0';
          end if;
        if(cVar1S12S70P017P014P012P049(0)='1' AND  A( 9)='0' AND A(10)='0' AND A( 0)='1' )then
          cVar2S12S70N001N018P019nsss(0) <='1';
          else
          cVar2S12S70N001N018P019nsss(0) <='0';
          end if;
        if(cVar1S13S70N017P066P044P032(0)='1' AND  B(17)='0' AND E( 4)='0' AND E( 0)='0' )then
          cVar2S13S70P020P052P068nsss(0) <='1';
          else
          cVar2S13S70P020P052P068nsss(0) <='0';
          end if;
        if(cVar1S14S70N017P066P044P032(0)='1' AND  B(17)='0' AND E( 4)='1' AND D(10)='0' )then
          cVar2S14S70P020P052P059nsss(0) <='1';
          else
          cVar2S14S70P020P052P059nsss(0) <='0';
          end if;
        if(cVar1S15S70N017P066P044P032(0)='1' AND  B(17)='1' AND D(10)='0' )then
          cVar2S15S70P020P059nsss(0) <='1';
          else
          cVar2S15S70P020P059nsss(0) <='0';
          end if;
        if(cVar1S16S70N017P066P044N032(0)='1' AND  E( 8)='1' AND A(13)='0' AND D( 8)='1' )then
          cVar2S16S70P069P012P067nsss(0) <='1';
          else
          cVar2S16S70P069P012P067nsss(0) <='0';
          end if;
        if(cVar1S17S70N017P066P044N032(0)='1' AND  E( 8)='0' AND B( 4)='1' AND A(19)='0' )then
          cVar2S17S70N069P029P000nsss(0) <='1';
          else
          cVar2S17S70N069P029P000nsss(0) <='0';
          end if;
        if(cVar1S18S70N017P066P044N032(0)='1' AND  E( 8)='0' AND B( 4)='0' AND A( 2)='1' )then
          cVar2S18S70N069N029P015nsss(0) <='1';
          else
          cVar2S18S70N069N029P015nsss(0) <='0';
          end if;
        if(cVar1S19S70N017P066P044P045(0)='1' AND  E( 5)='0' AND B( 0)='1' )then
          cVar2S19S70P048P037nsss(0) <='1';
          else
          cVar2S19S70P048P037nsss(0) <='0';
          end if;
        if(cVar1S20S70N017P066P044P045(0)='1' AND  E( 5)='0' AND B( 0)='0' AND B( 7)='1' )then
          cVar2S20S70P048N037P023nsss(0) <='1';
          else
          cVar2S20S70P048N037P023nsss(0) <='0';
          end if;
        if(cVar1S21S70N017P066P044P045(0)='1' AND  E( 5)='1' AND D( 5)='0' )then
          cVar2S21S70P048P046nsss(0) <='1';
          else
          cVar2S21S70P048P046nsss(0) <='0';
          end if;
        if(cVar1S22S70N017P066P004P034(0)='1' AND  B(17)='0' AND B(11)='0' AND A(14)='0' )then
          cVar2S22S70P020P032P010nsss(0) <='1';
          else
          cVar2S22S70P020P032P010nsss(0) <='0';
          end if;
        if(cVar1S23S70N017P066P004N034(0)='1' AND  B(17)='1' AND E( 0)='1' )then
          cVar2S23S70P020P068nsss(0) <='1';
          else
          cVar2S23S70P020P068nsss(0) <='0';
          end if;
        if(cVar1S24S70N017P066P004N034(0)='1' AND  B(17)='0' AND E( 9)='0' AND B( 9)='1' )then
          cVar2S24S70N020P065P036nsss(0) <='1';
          else
          cVar2S24S70N020P065P036nsss(0) <='0';
          end if;
        if(cVar1S26S70N017P066P004N061(0)='1' AND  D( 6)='1' )then
          cVar2S26S70P042nsss(0) <='1';
          else
          cVar2S26S70P042nsss(0) <='0';
          end if;
        if(cVar1S27S70N017P066P004N061(0)='1' AND  D( 6)='0' AND B( 0)='1' AND A( 5)='1' )then
          cVar2S27S70N042P037P009nsss(0) <='1';
          else
          cVar2S27S70N042P037P009nsss(0) <='0';
          end if;
        if(cVar1S0S71P067P015P018P069(0)='1' AND  A(11)='0' AND E( 2)='0' )then
          cVar2S0S71P016P060nsss(0) <='1';
          else
          cVar2S0S71P016P060nsss(0) <='0';
          end if;
        if(cVar1S1S71P067P015P018P069(0)='1' AND  A(11)='0' AND E( 2)='1' AND A( 3)='1' )then
          cVar2S1S71P016P060P013nsss(0) <='1';
          else
          cVar2S1S71P016P060P013nsss(0) <='0';
          end if;
        if(cVar1S2S71P067P015P018P069(0)='1' AND  A(11)='1' AND D(11)='0' AND A( 6)='1' )then
          cVar2S2S71P016P055P007nsss(0) <='1';
          else
          cVar2S2S71P016P055P007nsss(0) <='0';
          end if;
        if(cVar1S3S71P067P015P018P069(0)='1' AND  A(11)='1' AND D(11)='1' AND E( 9)='1' )then
          cVar2S3S71P016P055P065nsss(0) <='1';
          else
          cVar2S3S71P016P055P065nsss(0) <='0';
          end if;
        if(cVar1S4S71P067P015P018P069(0)='1' AND  A( 0)='1' AND D( 0)='1' AND B( 0)='1' )then
          cVar2S4S71P019P066P037nsss(0) <='1';
          else
          cVar2S4S71P019P066P037nsss(0) <='0';
          end if;
        if(cVar1S5S71P067P015P018P069(0)='1' AND  A( 0)='0' AND D( 9)='1' AND A(11)='0' )then
          cVar2S5S71N019P063P016nsss(0) <='1';
          else
          cVar2S5S71N019P063P016nsss(0) <='0';
          end if;
        if(cVar1S6S71P067P015N018P002(0)='1' AND  B( 2)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar2S6S71P033P021P040nsss(0) <='1';
          else
          cVar2S6S71P033P021P040nsss(0) <='0';
          end if;
        if(cVar1S7S71P067P015N018P002(0)='1' AND  B( 2)='0' AND B( 8)='0' AND E(10)='0' )then
          cVar2S7S71P033N021P061nsss(0) <='1';
          else
          cVar2S7S71P033N021P061nsss(0) <='0';
          end if;
        if(cVar1S8S71P067P015N018N002(0)='1' AND  A(12)='1' AND A( 6)='0' AND A( 3)='0' )then
          cVar2S8S71P014P007P013nsss(0) <='1';
          else
          cVar2S8S71P014P007P013nsss(0) <='0';
          end if;
        if(cVar1S9S71P067P015N018N002(0)='1' AND  A(12)='1' AND A( 6)='1' AND B(15)='1' )then
          cVar2S9S71P014P007P024nsss(0) <='1';
          else
          cVar2S9S71P014P007P024nsss(0) <='0';
          end if;
        if(cVar1S10S71P067P015N018N002(0)='1' AND  A(12)='0' AND A(11)='1' AND A( 6)='0' )then
          cVar2S10S71N014P016P007nsss(0) <='1';
          else
          cVar2S10S71N014P016P007nsss(0) <='0';
          end if;
        if(cVar1S11S71P067P015N018N002(0)='1' AND  A(12)='0' AND A(11)='0' AND A(13)='1' )then
          cVar2S11S71N014N016P012nsss(0) <='1';
          else
          cVar2S11S71N014N016P012nsss(0) <='0';
          end if;
        if(cVar1S12S71P067P015P017P069(0)='1' AND  A( 3)='0' AND A( 0)='1' AND A(13)='0' )then
          cVar2S12S71P013P019P012nsss(0) <='1';
          else
          cVar2S12S71P013P019P012nsss(0) <='0';
          end if;
        if(cVar1S13S71P067P015P017P069(0)='1' AND  A( 3)='0' AND A( 0)='0' AND A(10)='0' )then
          cVar2S13S71P013N019P018nsss(0) <='1';
          else
          cVar2S13S71P013N019P018nsss(0) <='0';
          end if;
        if(cVar1S14S71P067P015P017P069(0)='1' AND  A( 3)='1' AND A( 0)='0' )then
          cVar2S14S71P013P019nsss(0) <='1';
          else
          cVar2S14S71P013P019nsss(0) <='0';
          end if;
        if(cVar1S15S71P067P015P017N069(0)='1' AND  B(13)='1' AND A( 0)='0' AND B( 1)='0' )then
          cVar2S15S71P028P019P035nsss(0) <='1';
          else
          cVar2S15S71P028P019P035nsss(0) <='0';
          end if;
        if(cVar1S16S71P067P015P017N069(0)='1' AND  B(13)='1' AND A( 0)='1' AND A(14)='1' )then
          cVar2S16S71P028P019P010nsss(0) <='1';
          else
          cVar2S16S71P028P019P010nsss(0) <='0';
          end if;
        if(cVar1S17S71P067P015P017N069(0)='1' AND  B(13)='0' AND A( 3)='1' )then
          cVar2S17S71N028P013nsss(0) <='1';
          else
          cVar2S17S71N028P013nsss(0) <='0';
          end if;
        if(cVar1S18S71P067P015P017N069(0)='1' AND  B(13)='0' AND A( 3)='0' AND B(16)='0' )then
          cVar2S18S71N028N013P022nsss(0) <='1';
          else
          cVar2S18S71N028N013P022nsss(0) <='0';
          end if;
        if(cVar1S19S71P067P015N017P026(0)='1' AND  B(10)='0' AND A(16)='1' AND A(15)='0' )then
          cVar2S19S71P034P006P008nsss(0) <='1';
          else
          cVar2S19S71P034P006P008nsss(0) <='0';
          end if;
        if(cVar1S20S71P067P015N017P026(0)='1' AND  B(10)='0' AND A(16)='0' AND A( 0)='0' )then
          cVar2S20S71P034N006P019nsss(0) <='1';
          else
          cVar2S20S71P034N006P019nsss(0) <='0';
          end if;
        if(cVar1S21S71P067P015N017P026(0)='1' AND  B(10)='1' AND B( 5)='1' )then
          cVar2S21S71P034P027nsss(0) <='1';
          else
          cVar2S21S71P034P027nsss(0) <='0';
          end if;
        if(cVar1S22S71P067P015N017P026(0)='1' AND  D(11)='0' AND A(17)='0' AND A( 5)='1' )then
          cVar2S22S71P055P004P009nsss(0) <='1';
          else
          cVar2S22S71P055P004P009nsss(0) <='0';
          end if;
        if(cVar1S23S71P067P001P057P037(0)='1' AND  B(10)='1' )then
          cVar2S23S71P034nsss(0) <='1';
          else
          cVar2S23S71P034nsss(0) <='0';
          end if;
        if(cVar1S24S71P067P001P057P037(0)='1' AND  B(10)='0' AND A(13)='1' AND B( 9)='0' )then
          cVar2S24S71N034P012P036nsss(0) <='1';
          else
          cVar2S24S71N034P012P036nsss(0) <='0';
          end if;
        if(cVar1S25S71P067P001P057P037(0)='1' AND  B(10)='0' AND A(13)='0' AND A( 5)='0' )then
          cVar2S25S71N034N012P009nsss(0) <='1';
          else
          cVar2S25S71N034N012P009nsss(0) <='0';
          end if;
        if(cVar1S26S71P067P001P057P037(0)='1' AND  A( 0)='1' AND A( 1)='0' )then
          cVar2S26S71P019P017nsss(0) <='1';
          else
          cVar2S26S71P019P017nsss(0) <='0';
          end if;
        if(cVar1S27S71P067N001P003P054(0)='1' AND  D( 6)='0' AND A( 3)='0' AND A( 4)='0' )then
          cVar2S27S71P042P013P011nsss(0) <='1';
          else
          cVar2S27S71P042P013P011nsss(0) <='0';
          end if;
        if(cVar1S28S71P067N001P003P054(0)='1' AND  D( 6)='0' AND A( 3)='1' AND B(10)='0' )then
          cVar2S28S71P042P013P034nsss(0) <='1';
          else
          cVar2S28S71P042P013P034nsss(0) <='0';
          end if;
        if(cVar1S29S71P067N001N003P045(0)='1' AND  A( 5)='1' AND A( 0)='1' AND A( 2)='0' )then
          cVar2S29S71P009P019P015nsss(0) <='1';
          else
          cVar2S29S71P009P019P015nsss(0) <='0';
          end if;
        if(cVar1S30S71P067N001N003P045(0)='1' AND  A( 5)='0' AND A(19)='1' AND B( 9)='1' )then
          cVar2S30S71N009P000P036nsss(0) <='1';
          else
          cVar2S30S71N009P000P036nsss(0) <='0';
          end if;
        if(cVar1S31S71P067N001N003P045(0)='1' AND  A(10)='0' AND A( 0)='1' )then
          cVar2S31S71P018P019nsss(0) <='1';
          else
          cVar2S31S71P018P019nsss(0) <='0';
          end if;
        if(cVar1S32S71P067N001N003P045(0)='1' AND  A(10)='1' AND D(13)='0' AND A( 6)='1' )then
          cVar2S32S71P018P047P007nsss(0) <='1';
          else
          cVar2S32S71P018P047P007nsss(0) <='0';
          end if;
        if(cVar1S0S72P069P045P052P056(0)='1' AND  A(16)='0' )then
          cVar2S0S72P006nsss(0) <='1';
          else
          cVar2S0S72P006nsss(0) <='0';
          end if;
        if(cVar1S1S72P069P045N052P029(0)='1' AND  A( 3)='1' AND B( 8)='0' )then
          cVar2S1S72P013P021nsss(0) <='1';
          else
          cVar2S1S72P013P021nsss(0) <='0';
          end if;
        if(cVar1S2S72P069P045N052P029(0)='1' AND  A( 3)='0' AND A(16)='1' )then
          cVar2S2S72N013P006nsss(0) <='1';
          else
          cVar2S2S72N013P006nsss(0) <='0';
          end if;
        if(cVar1S3S72P069P045N052P029(0)='1' AND  A( 3)='0' AND A(16)='0' AND E( 6)='0' )then
          cVar2S3S72N013N006P044nsss(0) <='1';
          else
          cVar2S3S72N013N006P044nsss(0) <='0';
          end if;
        if(cVar1S4S72P069P045N052P029(0)='1' AND  D( 3)='1' AND A(10)='0' )then
          cVar2S4S72P054P018nsss(0) <='1';
          else
          cVar2S4S72P054P018nsss(0) <='0';
          end if;
        if(cVar1S5S72P069P045N052P029(0)='1' AND  D( 3)='1' AND A(10)='1' AND B( 9)='0' )then
          cVar2S5S72P054P018P036nsss(0) <='1';
          else
          cVar2S5S72P054P018P036nsss(0) <='0';
          end if;
        if(cVar1S6S72P069P045N052P029(0)='1' AND  D( 3)='0' AND E( 2)='1' )then
          cVar2S6S72N054P060nsss(0) <='1';
          else
          cVar2S6S72N054P060nsss(0) <='0';
          end if;
        if(cVar1S7S72P069P045N052P029(0)='1' AND  D( 3)='0' AND E( 2)='0' AND E(12)='1' )then
          cVar2S7S72N054N060P053nsss(0) <='1';
          else
          cVar2S7S72N054N060P053nsss(0) <='0';
          end if;
        if(cVar1S9S72P069P045P018N006(0)='1' AND  D( 8)='1' )then
          cVar2S9S72P067nsss(0) <='1';
          else
          cVar2S9S72P067nsss(0) <='0';
          end if;
        if(cVar1S10S72P069P045P018P047(0)='1' AND  A( 2)='0' AND A( 0)='1' )then
          cVar2S10S72P015P019nsss(0) <='1';
          else
          cVar2S10S72P015P019nsss(0) <='0';
          end if;
        if(cVar1S11S72N069P015P027P008(0)='1' AND  A(16)='0' AND A( 1)='0' )then
          cVar2S11S72P006P017nsss(0) <='1';
          else
          cVar2S11S72P006P017nsss(0) <='0';
          end if;
        if(cVar1S12S72N069P015P027P008(0)='1' AND  A(16)='0' AND A( 1)='1' AND B( 1)='1' )then
          cVar2S12S72P006P017P035nsss(0) <='1';
          else
          cVar2S12S72P006P017P035nsss(0) <='0';
          end if;
        if(cVar1S13S72N069P015P027N008(0)='1' AND  A(13)='0' AND B( 6)='0' )then
          cVar2S13S72P012P025nsss(0) <='1';
          else
          cVar2S13S72P012P025nsss(0) <='0';
          end if;
        if(cVar1S14S72N069P015P027N008(0)='1' AND  A(13)='1' AND A(14)='0' AND A( 5)='1' )then
          cVar2S14S72P012P010P009nsss(0) <='1';
          else
          cVar2S14S72P012P010P009nsss(0) <='0';
          end if;
        if(cVar1S15S72N069P015N027P000(0)='1' AND  B(17)='1' AND D( 4)='0' )then
          cVar2S15S72P020P050nsss(0) <='1';
          else
          cVar2S15S72P020P050nsss(0) <='0';
          end if;
        if(cVar1S16S72N069P015N027P000(0)='1' AND  B(17)='0' AND A(11)='0' )then
          cVar2S16S72N020P016nsss(0) <='1';
          else
          cVar2S16S72N020P016nsss(0) <='0';
          end if;
        if(cVar1S17S72N069P015N027P000(0)='1' AND  B(17)='0' AND A(11)='1' AND E(12)='1' )then
          cVar2S17S72N020P016P053nsss(0) <='1';
          else
          cVar2S17S72N020P016P053nsss(0) <='0';
          end if;
        if(cVar1S18S72N069P015N027P000(0)='1' AND  B( 3)='1' )then
          cVar2S18S72P031nsss(0) <='1';
          else
          cVar2S18S72P031nsss(0) <='0';
          end if;
        if(cVar1S19S72N069P015N027P000(0)='1' AND  B( 3)='0' AND E(12)='0' AND B(12)='1' )then
          cVar2S19S72N031P053P030nsss(0) <='1';
          else
          cVar2S19S72N031P053P030nsss(0) <='0';
          end if;
        if(cVar1S20S72N069P015P028P026(0)='1' AND  D(10)='0' AND E(11)='1' AND A( 3)='0' )then
          cVar2S20S72P059P057P013nsss(0) <='1';
          else
          cVar2S20S72P059P057P013nsss(0) <='0';
          end if;
        if(cVar1S21S72N069P015P028P026(0)='1' AND  D(10)='0' AND E(11)='0' AND A(14)='1' )then
          cVar2S21S72P059N057P010nsss(0) <='1';
          else
          cVar2S21S72P059N057P010nsss(0) <='0';
          end if;
        if(cVar1S22S72N069P015P028P026(0)='1' AND  D(10)='1' AND B( 2)='0' )then
          cVar2S22S72P059P033nsss(0) <='1';
          else
          cVar2S22S72P059P033nsss(0) <='0';
          end if;
        if(cVar1S23S72N069P015N028P020(0)='1' AND  D(15)='0' AND E( 6)='1' )then
          cVar2S23S72P039P044nsss(0) <='1';
          else
          cVar2S23S72P039P044nsss(0) <='0';
          end if;
        if(cVar1S24S72N069P015N028P020(0)='1' AND  D(15)='1' AND A( 8)='1' )then
          cVar2S24S72P039P003nsss(0) <='1';
          else
          cVar2S24S72P039P003nsss(0) <='0';
          end if;
        if(cVar1S25S72N069P015N028P020(0)='1' AND  D(15)='1' AND A( 8)='0' AND B( 1)='1' )then
          cVar2S25S72P039N003P035nsss(0) <='1';
          else
          cVar2S25S72P039N003P035nsss(0) <='0';
          end if;
        if(cVar1S26S72N069P015N028P020(0)='1' AND  A(11)='0' AND E(10)='1' )then
          cVar2S26S72P016P061nsss(0) <='1';
          else
          cVar2S26S72P016P061nsss(0) <='0';
          end if;
        if(cVar1S27S72N069P015N028P020(0)='1' AND  A(11)='1' AND B( 2)='0' AND A(15)='1' )then
          cVar2S27S72P016P033P008nsss(0) <='1';
          else
          cVar2S27S72P016P033P008nsss(0) <='0';
          end if;
        if(cVar1S0S73P016P038P043P045(0)='1' AND  A( 8)='0' )then
          cVar2S0S73P003nsss(0) <='1';
          else
          cVar2S0S73P003nsss(0) <='0';
          end if;
        if(cVar1S1S73P016P038P043N045(0)='1' AND  E( 9)='1' )then
          cVar2S1S73P065nsss(0) <='1';
          else
          cVar2S1S73P065nsss(0) <='0';
          end if;
        if(cVar1S2S73P016P038P043N045(0)='1' AND  E( 9)='0' AND E( 0)='1' )then
          cVar2S2S73N065P068nsss(0) <='1';
          else
          cVar2S2S73N065P068nsss(0) <='0';
          end if;
        if(cVar1S3S73P016P038P043N045(0)='1' AND  E( 9)='0' AND E( 0)='0' AND A(13)='1' )then
          cVar2S3S73N065N068P012nsss(0) <='1';
          else
          cVar2S3S73N065N068P012nsss(0) <='0';
          end if;
        if(cVar1S4S73P016P038N043P045(0)='1' AND  A(10)='1' AND A( 7)='0' )then
          cVar2S4S73P018P005nsss(0) <='1';
          else
          cVar2S4S73P018P005nsss(0) <='0';
          end if;
        if(cVar1S5S73P016P038N043P045(0)='1' AND  A(10)='1' AND A( 7)='1' AND A(18)='1' )then
          cVar2S5S73P018P005P002nsss(0) <='1';
          else
          cVar2S5S73P018P005P002nsss(0) <='0';
          end if;
        if(cVar1S6S73P016P038N043P045(0)='1' AND  A(10)='0' AND D(10)='0' AND A(19)='0' )then
          cVar2S6S73N018P059P000nsss(0) <='1';
          else
          cVar2S6S73N018P059P000nsss(0) <='0';
          end if;
        if(cVar1S7S73P016P038N043P045(0)='1' AND  A(10)='0' AND D(10)='1' AND B(10)='1' )then
          cVar2S7S73N018P059P034nsss(0) <='1';
          else
          cVar2S7S73N018P059P034nsss(0) <='0';
          end if;
        if(cVar1S8S73P016P038N043P045(0)='1' AND  A( 4)='1' AND A(12)='0' )then
          cVar2S8S73P011P014nsss(0) <='1';
          else
          cVar2S8S73P011P014nsss(0) <='0';
          end if;
        if(cVar1S9S73P016P038N043P045(0)='1' AND  A( 4)='0' AND A( 5)='1' )then
          cVar2S9S73N011P009nsss(0) <='1';
          else
          cVar2S9S73N011P009nsss(0) <='0';
          end if;
        if(cVar1S10S73P016P038N043P045(0)='1' AND  A( 4)='0' AND A( 5)='0' AND B( 2)='1' )then
          cVar2S10S73N011N009P033nsss(0) <='1';
          else
          cVar2S10S73N011N009P033nsss(0) <='0';
          end if;
        if(cVar1S11S73P016P038P033P018(0)='1' AND  D( 0)='1' )then
          cVar2S11S73P066nsss(0) <='1';
          else
          cVar2S11S73P066nsss(0) <='0';
          end if;
        if(cVar1S12S73P016P038P033P018(0)='1' AND  D( 0)='0' AND A(13)='1' )then
          cVar2S12S73N066P012nsss(0) <='1';
          else
          cVar2S12S73N066P012nsss(0) <='0';
          end if;
        if(cVar1S13S73N016P036P027P014(0)='1' AND  A( 5)='1' )then
          cVar2S13S73P009nsss(0) <='1';
          else
          cVar2S13S73P009nsss(0) <='0';
          end if;
        if(cVar1S14S73N016P036P027P014(0)='1' AND  A( 5)='0' AND D( 8)='0' AND E( 5)='1' )then
          cVar2S14S73N009P067P048nsss(0) <='1';
          else
          cVar2S14S73N009P067P048nsss(0) <='0';
          end if;
        if(cVar1S15S73N016P036P027P014(0)='1' AND  A( 5)='0' AND D( 8)='1' AND A( 0)='0' )then
          cVar2S15S73N009P067P019nsss(0) <='1';
          else
          cVar2S15S73N009P067P019nsss(0) <='0';
          end if;
        if(cVar1S16S73N016P036P027P014(0)='1' AND  E( 5)='1' )then
          cVar2S16S73P048nsss(0) <='1';
          else
          cVar2S16S73P048nsss(0) <='0';
          end if;
        if(cVar1S17S73N016P036P027P014(0)='1' AND  E( 5)='0' AND D(12)='1' )then
          cVar2S17S73N048P051nsss(0) <='1';
          else
          cVar2S17S73N048P051nsss(0) <='0';
          end if;
        if(cVar1S18S73N016P036P027P014(0)='1' AND  E( 5)='0' AND D(12)='0' AND A( 4)='1' )then
          cVar2S18S73N048N051P011nsss(0) <='1';
          else
          cVar2S18S73N048N051P011nsss(0) <='0';
          end if;
        if(cVar1S19S73N016P036N027P038(0)='1' AND  A(18)='1' )then
          cVar2S19S73P002nsss(0) <='1';
          else
          cVar2S19S73P002nsss(0) <='0';
          end if;
        if(cVar1S20S73N016P036N027P038(0)='1' AND  A(18)='0' AND A(19)='1' )then
          cVar2S20S73N002P000nsss(0) <='1';
          else
          cVar2S20S73N002P000nsss(0) <='0';
          end if;
        if(cVar1S21S73N016P036N027P038(0)='1' AND  A(18)='0' AND A(19)='0' AND B( 8)='1' )then
          cVar2S21S73N002N000P021nsss(0) <='1';
          else
          cVar2S21S73N002N000P021nsss(0) <='0';
          end if;
        if(cVar1S22S73N016P036N027N038(0)='1' AND  B(13)='1' AND D(14)='1' )then
          cVar2S22S73P028P043nsss(0) <='1';
          else
          cVar2S22S73P028P043nsss(0) <='0';
          end if;
        if(cVar1S23S73N016P036N027N038(0)='1' AND  B(13)='1' AND D(14)='0' AND B(12)='0' )then
          cVar2S23S73P028N043P030nsss(0) <='1';
          else
          cVar2S23S73P028N043P030nsss(0) <='0';
          end if;
        if(cVar1S24S73N016P036N027N038(0)='1' AND  B(13)='0' AND D( 8)='1' AND B(10)='0' )then
          cVar2S24S73N028P067P034nsss(0) <='1';
          else
          cVar2S24S73N028P067P034nsss(0) <='0';
          end if;
        if(cVar1S25S73N016P036N027N038(0)='1' AND  B(13)='0' AND D( 8)='0' AND B( 1)='1' )then
          cVar2S25S73N028N067P035nsss(0) <='1';
          else
          cVar2S25S73N028N067P035nsss(0) <='0';
          end if;
        if(cVar1S26S73N016P036P045P068(0)='1' AND  A( 3)='1' AND A( 5)='0' )then
          cVar2S26S73P013P009nsss(0) <='1';
          else
          cVar2S26S73P013P009nsss(0) <='0';
          end if;
        if(cVar1S27S73N016P036P045P068(0)='1' AND  A( 3)='0' AND D(13)='1' AND E(13)='1' )then
          cVar2S27S73N013P047P049nsss(0) <='1';
          else
          cVar2S27S73N013P047P049nsss(0) <='0';
          end if;
        if(cVar1S28S73N016P036P045P068(0)='1' AND  D( 0)='1' AND E( 1)='1' AND D(10)='1' )then
          cVar2S28S73P066P064P059nsss(0) <='1';
          else
          cVar2S28S73P066P064P059nsss(0) <='0';
          end if;
        if(cVar1S29S73N016P036P045P068(0)='1' AND  D( 0)='0' AND A( 0)='1' AND E( 8)='1' )then
          cVar2S29S73N066P019P069nsss(0) <='1';
          else
          cVar2S29S73N066P019P069nsss(0) <='0';
          end if;
        if(cVar1S30S73N016P036P045P043(0)='1' AND  D( 8)='1' )then
          cVar2S30S73P067nsss(0) <='1';
          else
          cVar2S30S73P067nsss(0) <='0';
          end if;
        if(cVar1S0S74P016P053P035P026(0)='1' AND  E(13)='1' AND D( 2)='1' )then
          cVar2S0S74P049P058nsss(0) <='1';
          else
          cVar2S0S74P049P058nsss(0) <='0';
          end if;
        if(cVar1S1S74P016P053P035P026(0)='1' AND  E(13)='1' AND D( 2)='0' AND B(15)='0' )then
          cVar2S1S74P049N058P024nsss(0) <='1';
          else
          cVar2S1S74P049N058P024nsss(0) <='0';
          end if;
        if(cVar1S2S74P016P053P035P026(0)='1' AND  E(13)='0' AND D( 4)='1' )then
          cVar2S2S74N049P050nsss(0) <='1';
          else
          cVar2S2S74N049P050nsss(0) <='0';
          end if;
        if(cVar1S3S74P016P053P035P026(0)='1' AND  E(13)='0' AND D( 4)='0' AND E( 5)='1' )then
          cVar2S3S74N049N050P048nsss(0) <='1';
          else
          cVar2S3S74N049N050P048nsss(0) <='0';
          end if;
        if(cVar1S4S74P016P053P035N026(0)='1' AND  D(11)='1' AND A( 2)='1' )then
          cVar2S4S74P055P015nsss(0) <='1';
          else
          cVar2S4S74P055P015nsss(0) <='0';
          end if;
        if(cVar1S5S74P016P053P035N026(0)='1' AND  D(11)='1' AND A( 2)='0' AND D(12)='0' )then
          cVar2S5S74P055N015P051nsss(0) <='1';
          else
          cVar2S5S74P055N015P051nsss(0) <='0';
          end if;
        if(cVar1S6S74P016P053P035N026(0)='1' AND  D(11)='0' AND E(11)='0' AND B(16)='1' )then
          cVar2S6S74N055P057P022nsss(0) <='1';
          else
          cVar2S6S74N055P057P022nsss(0) <='0';
          end if;
        if(cVar1S7S74P016P053P035P052(0)='1' AND  A(14)='1' )then
          cVar2S7S74P010nsss(0) <='1';
          else
          cVar2S7S74P010nsss(0) <='0';
          end if;
        if(cVar1S8S74P016P053P035P052(0)='1' AND  A(14)='0' AND A(15)='1' )then
          cVar2S8S74N010P008nsss(0) <='1';
          else
          cVar2S8S74N010P008nsss(0) <='0';
          end if;
        if(cVar1S9S74P016P053P035P052(0)='1' AND  A(14)='0' AND A(15)='0' AND A(12)='1' )then
          cVar2S9S74N010N008P014nsss(0) <='1';
          else
          cVar2S9S74N010N008P014nsss(0) <='0';
          end if;
        if(cVar1S10S74P016P053P035N052(0)='1' AND  B(14)='0' AND B( 0)='1' AND A( 3)='0' )then
          cVar2S10S74P026P037P013nsss(0) <='1';
          else
          cVar2S10S74P026P037P013nsss(0) <='0';
          end if;
        if(cVar1S11S74P016P053P030P019(0)='1' AND  B(13)='1' )then
          cVar2S11S74P028nsss(0) <='1';
          else
          cVar2S11S74P028nsss(0) <='0';
          end if;
        if(cVar1S12S74P016P053P030P019(0)='1' AND  B(13)='0' AND D(12)='1' )then
          cVar2S12S74N028P051nsss(0) <='1';
          else
          cVar2S12S74N028P051nsss(0) <='0';
          end if;
        if(cVar1S13S74P016P053P030P019(0)='1' AND  B(13)='0' AND D(12)='0' AND D(11)='1' )then
          cVar2S13S74N028N051P055nsss(0) <='1';
          else
          cVar2S13S74N028N051P055nsss(0) <='0';
          end if;
        if(cVar1S14S74P016P053N030P059(0)='1' AND  E(11)='0' AND A( 4)='1' AND A(14)='0' )then
          cVar2S14S74P057P011P010nsss(0) <='1';
          else
          cVar2S14S74P057P011P010nsss(0) <='0';
          end if;
        if(cVar1S15S74P016P053N030P059(0)='1' AND  E(11)='1' AND D( 0)='0' AND D(12)='1' )then
          cVar2S15S74P057P066P051nsss(0) <='1';
          else
          cVar2S15S74P057P066P051nsss(0) <='0';
          end if;
        if(cVar1S16S74P016P053N030P059(0)='1' AND  B( 1)='1' )then
          cVar2S16S74P035nsss(0) <='1';
          else
          cVar2S16S74P035nsss(0) <='0';
          end if;
        if(cVar1S19S74P016P043N062N022(0)='1' AND  A(16)='1' )then
          cVar2S19S74P006nsss(0) <='1';
          else
          cVar2S19S74P006nsss(0) <='0';
          end if;
        if(cVar1S20S74P016P043N062N022(0)='1' AND  A(16)='0' AND E( 0)='1' AND A( 0)='0' )then
          cVar2S20S74N006P068P019nsss(0) <='1';
          else
          cVar2S20S74N006P068P019nsss(0) <='0';
          end if;
        if(cVar1S21S74P016N043P038P056(0)='1' AND  A(14)='1' AND E( 4)='1' )then
          cVar2S21S74P010P052nsss(0) <='1';
          else
          cVar2S21S74P010P052nsss(0) <='0';
          end if;
        if(cVar1S22S74P016N043P038P056(0)='1' AND  A(14)='1' AND E( 4)='0' AND B( 4)='0' )then
          cVar2S22S74P010N052P029nsss(0) <='1';
          else
          cVar2S22S74P010N052P029nsss(0) <='0';
          end if;
        if(cVar1S23S74P016N043P038P056(0)='1' AND  A(14)='0' AND D( 3)='1' AND A(12)='1' )then
          cVar2S23S74N010P054P014nsss(0) <='1';
          else
          cVar2S23S74N010P054P014nsss(0) <='0';
          end if;
        if(cVar1S24S74P016N043P038P056(0)='1' AND  A( 4)='0' AND B(14)='0' AND D( 8)='1' )then
          cVar2S24S74P011P026P067nsss(0) <='1';
          else
          cVar2S24S74P011P026P067nsss(0) <='0';
          end if;
        if(cVar1S25S74P016N043P038P056(0)='1' AND  A( 4)='1' AND A(14)='0' AND D(11)='1' )then
          cVar2S25S74P011P010P055nsss(0) <='1';
          else
          cVar2S25S74P011P010P055nsss(0) <='0';
          end if;
        if(cVar1S26S74P016N043P038P033(0)='1' AND  A(10)='0' AND D( 0)='1' )then
          cVar2S26S74P018P066nsss(0) <='1';
          else
          cVar2S26S74P018P066nsss(0) <='0';
          end if;
        if(cVar1S27S74P016N043P038P033(0)='1' AND  A(10)='0' AND D( 0)='0' AND A( 1)='1' )then
          cVar2S27S74P018N066P017nsss(0) <='1';
          else
          cVar2S27S74P018N066P017nsss(0) <='0';
          end if;
        if(cVar1S0S75P064P027P026P006(0)='1' AND  B( 0)='0' AND E( 5)='1' )then
          cVar2S0S75P037P048nsss(0) <='1';
          else
          cVar2S0S75P037P048nsss(0) <='0';
          end if;
        if(cVar1S1S75P064P027P026P006(0)='1' AND  B( 0)='0' AND E( 5)='0' AND E( 4)='1' )then
          cVar2S1S75P037N048P052nsss(0) <='1';
          else
          cVar2S1S75P037N048P052nsss(0) <='0';
          end if;
        if(cVar1S2S75P064P027P026N006(0)='1' AND  E(14)='0' AND A(12)='0' )then
          cVar2S2S75P045P014nsss(0) <='1';
          else
          cVar2S2S75P045P014nsss(0) <='0';
          end if;
        if(cVar1S3S75P064P027P026N006(0)='1' AND  E(14)='0' AND A(12)='1' AND D( 5)='1' )then
          cVar2S3S75P045P014P046nsss(0) <='1';
          else
          cVar2S3S75P045P014P046nsss(0) <='0';
          end if;
        if(cVar1S4S75P064P027P026P010(0)='1' AND  A( 5)='1' )then
          cVar2S4S75P009nsss(0) <='1';
          else
          cVar2S4S75P009nsss(0) <='0';
          end if;
        if(cVar1S5S75P064N027P060P054(0)='1' AND  E( 3)='0' AND B( 3)='1' AND B( 2)='0' )then
          cVar2S5S75P056P031P033nsss(0) <='1';
          else
          cVar2S5S75P056P031P033nsss(0) <='0';
          end if;
        if(cVar1S6S75P064N027P060P054(0)='1' AND  E( 3)='0' AND B( 3)='0' AND A(17)='0' )then
          cVar2S6S75P056N031P004nsss(0) <='1';
          else
          cVar2S6S75P056N031P004nsss(0) <='0';
          end if;
        if(cVar1S7S75P064N027P060P054(0)='1' AND  E( 3)='1' AND B(11)='1' )then
          cVar2S7S75P056P032nsss(0) <='1';
          else
          cVar2S7S75P056P032nsss(0) <='0';
          end if;
        if(cVar1S8S75P064N027P060P054(0)='1' AND  E( 3)='1' AND B(11)='0' AND A( 3)='1' )then
          cVar2S8S75P056N032P013nsss(0) <='1';
          else
          cVar2S8S75P056N032P013nsss(0) <='0';
          end if;
        if(cVar1S9S75P064N027P060P054(0)='1' AND  A( 4)='1' AND D( 0)='0' )then
          cVar2S9S75P011P066nsss(0) <='1';
          else
          cVar2S9S75P011P066nsss(0) <='0';
          end if;
        if(cVar1S10S75P064N027P060P054(0)='1' AND  A( 4)='0' AND D( 8)='0' AND A(13)='0' )then
          cVar2S10S75N011P067P012nsss(0) <='1';
          else
          cVar2S10S75N011P067P012nsss(0) <='0';
          end if;
        if(cVar1S11S75P064N027N060P062(0)='1' AND  A( 6)='1' AND A(15)='0' )then
          cVar2S11S75P007P008nsss(0) <='1';
          else
          cVar2S11S75P007P008nsss(0) <='0';
          end if;
        if(cVar1S12S75P064N027N060P062(0)='1' AND  A( 6)='0' AND A(11)='0' AND E(14)='0' )then
          cVar2S12S75N007P016P045nsss(0) <='1';
          else
          cVar2S12S75N007P016P045nsss(0) <='0';
          end if;
        if(cVar1S13S75P064N027N060P062(0)='1' AND  E( 9)='1' AND B( 0)='1' AND E( 8)='0' )then
          cVar2S13S75P065P037P069nsss(0) <='1';
          else
          cVar2S13S75P065P037P069nsss(0) <='0';
          end if;
        if(cVar1S14S75P064N027N060P062(0)='1' AND  E( 9)='1' AND B( 0)='0' AND D( 0)='0' )then
          cVar2S14S75P065N037P066nsss(0) <='1';
          else
          cVar2S14S75P065N037P066nsss(0) <='0';
          end if;
        if(cVar1S15S75P064N027N060P062(0)='1' AND  E( 9)='0' AND B(12)='1' AND A( 0)='1' )then
          cVar2S15S75N065P030P019nsss(0) <='1';
          else
          cVar2S15S75N065P030P019nsss(0) <='0';
          end if;
        if(cVar1S16S75P064N027N060P062(0)='1' AND  E( 9)='0' AND B(12)='0' AND D(12)='1' )then
          cVar2S16S75N065N030P051nsss(0) <='1';
          else
          cVar2S16S75N065N030P051nsss(0) <='0';
          end if;
        if(cVar1S17S75P064P003P046P058(0)='1' AND  A(13)='0' )then
          cVar2S17S75P012nsss(0) <='1';
          else
          cVar2S17S75P012nsss(0) <='0';
          end if;
        if(cVar1S18S75P064P003P046N058(0)='1' AND  A( 5)='1' AND B( 2)='0' )then
          cVar2S18S75P009P033nsss(0) <='1';
          else
          cVar2S18S75P009P033nsss(0) <='0';
          end if;
        if(cVar1S19S75P064P003P046N058(0)='1' AND  A( 5)='0' AND A(12)='1' AND D( 1)='1' )then
          cVar2S19S75N009P014P062nsss(0) <='1';
          else
          cVar2S19S75N009P014P062nsss(0) <='0';
          end if;
        if(cVar1S20S75P064P003P046N058(0)='1' AND  A( 5)='0' AND A(12)='0' AND B(11)='0' )then
          cVar2S20S75N009N014P032nsss(0) <='1';
          else
          cVar2S20S75N009N014P032nsss(0) <='0';
          end if;
        if(cVar1S21S75P064N003P018P065(0)='1' AND  A( 1)='0' AND E( 0)='0' AND D( 9)='1' )then
          cVar2S21S75P017P068P063nsss(0) <='1';
          else
          cVar2S21S75P017P068P063nsss(0) <='0';
          end if;
        if(cVar1S22S75P064N003P018P065(0)='1' AND  A( 1)='0' AND E( 0)='1' AND D( 1)='1' )then
          cVar2S22S75P017P068P062nsss(0) <='1';
          else
          cVar2S22S75P017P068P062nsss(0) <='0';
          end if;
        if(cVar1S23S75P064N003P018P065(0)='1' AND  A( 1)='1' AND D( 9)='0' )then
          cVar2S23S75P017P063nsss(0) <='1';
          else
          cVar2S23S75P017P063nsss(0) <='0';
          end if;
        if(cVar1S24S75P064N003P018P065(0)='1' AND  A( 1)='1' AND D( 9)='1' AND D( 8)='1' )then
          cVar2S24S75P017P063P067nsss(0) <='1';
          else
          cVar2S24S75P017P063P067nsss(0) <='0';
          end if;
        if(cVar1S25S75P064N003P018N065(0)='1' AND  A( 0)='0' AND A(13)='1' )then
          cVar2S25S75P019P012nsss(0) <='1';
          else
          cVar2S25S75P019P012nsss(0) <='0';
          end if;
        if(cVar1S26S75P064N003P018N065(0)='1' AND  A( 0)='0' AND A(13)='0' AND A(11)='0' )then
          cVar2S26S75P019N012P016nsss(0) <='1';
          else
          cVar2S26S75P019N012P016nsss(0) <='0';
          end if;
        if(cVar1S27S75P064N003P018N065(0)='1' AND  A( 0)='1' AND A( 2)='0' AND A( 4)='1' )then
          cVar2S27S75P019P015P011nsss(0) <='1';
          else
          cVar2S27S75P019P015P011nsss(0) <='0';
          end if;
        if(cVar1S28S75P064N003N018P013(0)='1' AND  B( 1)='1' )then
          cVar2S28S75P035nsss(0) <='1';
          else
          cVar2S28S75P035nsss(0) <='0';
          end if;
        if(cVar1S29S75P064N003N018P013(0)='1' AND  B( 1)='0' AND D( 8)='0' AND D( 9)='1' )then
          cVar2S29S75N035P067P063nsss(0) <='1';
          else
          cVar2S29S75N035P067P063nsss(0) <='0';
          end if;
        if(cVar1S30S75P064N003N018P013(0)='1' AND  B( 1)='0' AND D( 8)='1' AND A(12)='1' )then
          cVar2S30S75N035P067P014nsss(0) <='1';
          else
          cVar2S30S75N035P067P014nsss(0) <='0';
          end if;
        if(cVar1S31S75P064N003N018N013(0)='1' AND  D(11)='0' AND B(15)='1' )then
          cVar2S31S75P055P024nsss(0) <='1';
          else
          cVar2S31S75P055P024nsss(0) <='0';
          end if;
        if(cVar1S32S75P064N003N018N013(0)='1' AND  D(11)='1' AND E( 0)='1' )then
          cVar2S32S75P055P068nsss(0) <='1';
          else
          cVar2S32S75P055P068nsss(0) <='0';
          end if;
        if(cVar1S33S75P064N003N018N013(0)='1' AND  D(11)='1' AND E( 0)='0' AND E( 3)='1' )then
          cVar2S33S75P055N068P056nsss(0) <='1';
          else
          cVar2S33S75P055N068P056nsss(0) <='0';
          end if;
        if(cVar1S0S76P016P060P056P067(0)='1' AND  B( 2)='1' AND E( 9)='1' AND E( 0)='0' )then
          cVar2S0S76P033P065P068nsss(0) <='1';
          else
          cVar2S0S76P033P065P068nsss(0) <='0';
          end if;
        if(cVar1S1S76P016P060P056P067(0)='1' AND  B( 2)='1' AND E( 9)='0' AND D(10)='1' )then
          cVar2S1S76P033N065P059nsss(0) <='1';
          else
          cVar2S1S76P033N065P059nsss(0) <='0';
          end if;
        if(cVar1S2S76P016P060P056P067(0)='1' AND  B( 2)='0' AND B( 6)='0' )then
          cVar2S2S76N033P025nsss(0) <='1';
          else
          cVar2S2S76N033P025nsss(0) <='0';
          end if;
        if(cVar1S3S76P016P060P056P067(0)='1' AND  E( 4)='1' AND B( 4)='1' )then
          cVar2S3S76P052P029nsss(0) <='1';
          else
          cVar2S3S76P052P029nsss(0) <='0';
          end if;
        if(cVar1S4S76P016P060P056P067(0)='1' AND  E( 4)='1' AND B( 4)='0' AND A( 2)='0' )then
          cVar2S4S76P052N029P015nsss(0) <='1';
          else
          cVar2S4S76P052N029P015nsss(0) <='0';
          end if;
        if(cVar1S5S76P016P060P056P067(0)='1' AND  E( 4)='0' AND B( 4)='0' )then
          cVar2S5S76N052P029nsss(0) <='1';
          else
          cVar2S5S76N052P029nsss(0) <='0';
          end if;
        if(cVar1S6S76P016P060P056P011(0)='1' AND  B(14)='0' AND A(10)='1' )then
          cVar2S6S76P026P018nsss(0) <='1';
          else
          cVar2S6S76P026P018nsss(0) <='0';
          end if;
        if(cVar1S7S76P016P060P056P011(0)='1' AND  B(14)='0' AND A(10)='0' AND B(12)='1' )then
          cVar2S7S76P026N018P030nsss(0) <='1';
          else
          cVar2S7S76P026N018P030nsss(0) <='0';
          end if;
        if(cVar1S8S76P016P060P056P011(0)='1' AND  A(14)='0' AND E(11)='1' )then
          cVar2S8S76P010P057nsss(0) <='1';
          else
          cVar2S8S76P010P057nsss(0) <='0';
          end if;
        if(cVar1S9S76P016P060P015P064(0)='1' AND  B( 0)='0' )then
          cVar2S9S76P037nsss(0) <='1';
          else
          cVar2S9S76P037nsss(0) <='0';
          end if;
        if(cVar1S10S76P016P060P015P064(0)='1' AND  B( 0)='1' AND B( 1)='1' AND A( 0)='1' )then
          cVar2S10S76P037P035P019nsss(0) <='1';
          else
          cVar2S10S76P037P035P019nsss(0) <='0';
          end if;
        if(cVar1S11S76P016P060P015P064(0)='1' AND  B( 0)='1' AND B( 1)='0' AND B(10)='1' )then
          cVar2S11S76P037N035P034nsss(0) <='1';
          else
          cVar2S11S76P037N035P034nsss(0) <='0';
          end if;
        if(cVar1S12S76P016P060P015P064(0)='1' AND  D( 0)='1' AND D( 2)='1' )then
          cVar2S12S76P066P058nsss(0) <='1';
          else
          cVar2S12S76P066P058nsss(0) <='0';
          end if;
        if(cVar1S13S76P016P060P015P064(0)='1' AND  D( 0)='0' AND B( 2)='1' )then
          cVar2S13S76N066P033nsss(0) <='1';
          else
          cVar2S13S76N066P033nsss(0) <='0';
          end if;
        if(cVar1S14S76P016P060P015P020(0)='1' AND  B( 9)='0' AND A(15)='0' AND B( 1)='1' )then
          cVar2S14S76P036P008P035nsss(0) <='1';
          else
          cVar2S14S76P036P008P035nsss(0) <='0';
          end if;
        if(cVar1S15S76P016P060P015P020(0)='1' AND  B( 9)='1' AND D( 0)='1' AND A( 0)='0' )then
          cVar2S15S76P036P066P019nsss(0) <='1';
          else
          cVar2S15S76P036P066P019nsss(0) <='0';
          end if;
        if(cVar1S16S76N016P064P048P062(0)='1' AND  A( 9)='1' AND E( 0)='1' )then
          cVar2S16S76P001P068nsss(0) <='1';
          else
          cVar2S16S76P001P068nsss(0) <='0';
          end if;
        if(cVar1S17S76N016P064P048P062(0)='1' AND  A( 9)='1' AND E( 0)='0' AND B( 0)='0' )then
          cVar2S17S76P001N068P037nsss(0) <='1';
          else
          cVar2S17S76P001N068P037nsss(0) <='0';
          end if;
        if(cVar1S18S76N016P064P048P062(0)='1' AND  A( 9)='0' AND A( 4)='0' )then
          cVar2S18S76N001P011nsss(0) <='1';
          else
          cVar2S18S76N001P011nsss(0) <='0';
          end if;
        if(cVar1S19S76N016P064P048N062(0)='1' AND  B(11)='1' AND B( 0)='0' )then
          cVar2S19S76P032P037nsss(0) <='1';
          else
          cVar2S19S76P032P037nsss(0) <='0';
          end if;
        if(cVar1S20S76N016P064P048N062(0)='1' AND  B(11)='1' AND B( 0)='1' AND A( 1)='0' )then
          cVar2S20S76P032P037P017nsss(0) <='1';
          else
          cVar2S20S76P032P037P017nsss(0) <='0';
          end if;
        if(cVar1S21S76N016P064P048N062(0)='1' AND  B(11)='0' AND E( 4)='1' )then
          cVar2S21S76N032P052nsss(0) <='1';
          else
          cVar2S21S76N032P052nsss(0) <='0';
          end if;
        if(cVar1S22S76N016P064P048P058(0)='1' AND  B( 6)='1' )then
          cVar2S22S76P025nsss(0) <='1';
          else
          cVar2S22S76P025nsss(0) <='0';
          end if;
        if(cVar1S23S76N016P064P048P058(0)='1' AND  B( 6)='0' AND D( 0)='1' AND A( 0)='0' )then
          cVar2S23S76N025P066P019nsss(0) <='1';
          else
          cVar2S23S76N025P066P019nsss(0) <='0';
          end if;
        if(cVar1S24S76N016N064P027P006(0)='1' AND  B( 0)='0' )then
          cVar2S24S76P037nsss(0) <='1';
          else
          cVar2S24S76P037nsss(0) <='0';
          end if;
        if(cVar1S25S76N016N064P027N006(0)='1' AND  B( 3)='0' AND B(12)='1' )then
          cVar2S25S76P031P030nsss(0) <='1';
          else
          cVar2S25S76P031P030nsss(0) <='0';
          end if;
        if(cVar1S26S76N016N064P027N006(0)='1' AND  B( 3)='0' AND B(12)='0' AND A(15)='1' )then
          cVar2S26S76P031N030P008nsss(0) <='1';
          else
          cVar2S26S76P031N030P008nsss(0) <='0';
          end if;
        if(cVar1S27S76N016N064N027P057(0)='1' AND  B( 1)='0' AND E(12)='0' AND A( 6)='1' )then
          cVar2S27S76P035P053P007nsss(0) <='1';
          else
          cVar2S27S76P035P053P007nsss(0) <='0';
          end if;
        if(cVar1S28S76N016N064N027P057(0)='1' AND  B( 1)='0' AND E(12)='1' AND A(10)='1' )then
          cVar2S28S76P035P053P018nsss(0) <='1';
          else
          cVar2S28S76P035P053P018nsss(0) <='0';
          end if;
        if(cVar1S29S76N016N064N027P057(0)='1' AND  B( 1)='1' AND B( 2)='1' AND A(17)='0' )then
          cVar2S29S76P035P033P004nsss(0) <='1';
          else
          cVar2S29S76P035P033P004nsss(0) <='0';
          end if;
        if(cVar1S30S76N016N064N027P057(0)='1' AND  A( 2)='1' AND A( 4)='1' AND B( 2)='0' )then
          cVar2S30S76P015P011P033nsss(0) <='1';
          else
          cVar2S30S76P015P011P033nsss(0) <='0';
          end if;
        if(cVar1S31S76N016N064N027P057(0)='1' AND  A( 2)='1' AND A( 4)='0' AND D( 3)='1' )then
          cVar2S31S76P015N011P054nsss(0) <='1';
          else
          cVar2S31S76P015N011P054nsss(0) <='0';
          end if;
        if(cVar1S32S76N016N064N027P057(0)='1' AND  A( 2)='0' AND A(14)='1' AND E( 3)='0' )then
          cVar2S32S76N015P010P056nsss(0) <='1';
          else
          cVar2S32S76N015P010P056nsss(0) <='0';
          end if;
        if(cVar1S33S76N016N064N027P057(0)='1' AND  A( 2)='0' AND A(14)='0' AND A(12)='1' )then
          cVar2S33S76N015N010P014nsss(0) <='1';
          else
          cVar2S33S76N015N010P014nsss(0) <='0';
          end if;
        if(cVar1S0S77P035P053P016P057(0)='1' AND  E( 1)='0' AND A(10)='0' )then
          cVar2S0S77P064P018nsss(0) <='1';
          else
          cVar2S0S77P064P018nsss(0) <='0';
          end if;
        if(cVar1S1S77P035P053P016P057(0)='1' AND  E( 1)='0' AND A(10)='1' AND D( 1)='0' )then
          cVar2S1S77P064P018P062nsss(0) <='1';
          else
          cVar2S1S77P064P018P062nsss(0) <='0';
          end if;
        if(cVar1S2S77P035P053P016P057(0)='1' AND  E( 1)='1' AND A(19)='0' AND E( 6)='0' )then
          cVar2S2S77P064P000P044nsss(0) <='1';
          else
          cVar2S2S77P064P000P044nsss(0) <='0';
          end if;
        if(cVar1S3S77P035P053P016P057(0)='1' AND  E( 1)='1' AND A(19)='1' AND B( 2)='1' )then
          cVar2S3S77P064P000P033nsss(0) <='1';
          else
          cVar2S3S77P064P000P033nsss(0) <='0';
          end if;
        if(cVar1S4S77P035P053P016P057(0)='1' AND  D(12)='0' AND A(10)='1' )then
          cVar2S4S77P051P018nsss(0) <='1';
          else
          cVar2S4S77P051P018nsss(0) <='0';
          end if;
        if(cVar1S5S77P035P053P016P057(0)='1' AND  D(12)='0' AND A(10)='0' AND A( 4)='1' )then
          cVar2S5S77P051N018P011nsss(0) <='1';
          else
          cVar2S5S77P051N018P011nsss(0) <='0';
          end if;
        if(cVar1S6S77P035P053P016P028(0)='1' AND  A(12)='1' AND B(12)='0' )then
          cVar2S6S77P014P030nsss(0) <='1';
          else
          cVar2S6S77P014P030nsss(0) <='0';
          end if;
        if(cVar1S7S77P035P053P016P028(0)='1' AND  A(12)='1' AND B(12)='1' AND D( 1)='1' )then
          cVar2S7S77P014P030P062nsss(0) <='1';
          else
          cVar2S7S77P014P030P062nsss(0) <='0';
          end if;
        if(cVar1S8S77P035P053P016P028(0)='1' AND  A(12)='0' AND A( 4)='0' AND B(17)='0' )then
          cVar2S8S77N014P011P020nsss(0) <='1';
          else
          cVar2S8S77N014P011P020nsss(0) <='0';
          end if;
        if(cVar1S9S77P035P053P016P028(0)='1' AND  A(12)='0' AND A( 4)='1' AND B( 2)='1' )then
          cVar2S9S77N014P011P033nsss(0) <='1';
          else
          cVar2S9S77N014P011P033nsss(0) <='0';
          end if;
        if(cVar1S10S77P035P053P016P028(0)='1' AND  A( 3)='0' AND B( 0)='1' AND A( 0)='1' )then
          cVar2S10S77P013P037P019nsss(0) <='1';
          else
          cVar2S10S77P013P037P019nsss(0) <='0';
          end if;
        if(cVar1S11S77P035P053P016P028(0)='1' AND  A( 4)='1' )then
          cVar2S11S77P011nsss(0) <='1';
          else
          cVar2S11S77P011nsss(0) <='0';
          end if;
        if(cVar1S12S77P035P053P016P028(0)='1' AND  A( 4)='0' AND A( 2)='1' )then
          cVar2S12S77N011P015nsss(0) <='1';
          else
          cVar2S12S77N011P015nsss(0) <='0';
          end if;
        if(cVar1S13S77P035P053P016P028(0)='1' AND  A( 4)='0' AND A( 2)='0' AND A(14)='1' )then
          cVar2S13S77N011N015P010nsss(0) <='1';
          else
          cVar2S13S77N011N015P010nsss(0) <='0';
          end if;
        if(cVar1S14S77P035P053P016N028(0)='1' AND  A(19)='0' AND D(13)='0' AND A( 5)='1' )then
          cVar2S14S77P000P047P009nsss(0) <='1';
          else
          cVar2S14S77P000P047P009nsss(0) <='0';
          end if;
        if(cVar1S15S77P035P053N016P059(0)='1' AND  A( 2)='1' AND A(14)='1' AND B(13)='1' )then
          cVar2S15S77P015P010P028nsss(0) <='1';
          else
          cVar2S15S77P015P010P028nsss(0) <='0';
          end if;
        if(cVar1S16S77P035P053N016P059(0)='1' AND  A( 2)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar2S16S77P015N010P011nsss(0) <='1';
          else
          cVar2S16S77P015N010P011nsss(0) <='0';
          end if;
        if(cVar1S17S77P035P053N016P059(0)='1' AND  A( 2)='0' AND A( 9)='1' )then
          cVar2S17S77N015P001nsss(0) <='1';
          else
          cVar2S17S77N015P001nsss(0) <='0';
          end if;
        if(cVar1S18S77P035P053N016P059(0)='1' AND  A( 2)='0' AND A( 9)='0' AND B( 3)='1' )then
          cVar2S18S77N015N001P031nsss(0) <='1';
          else
          cVar2S18S77N015N001P031nsss(0) <='0';
          end if;
        if(cVar1S19S77P035P053N016P059(0)='1' AND  E( 8)='0' AND E( 2)='0' AND B(11)='1' )then
          cVar2S19S77P069P060P032nsss(0) <='1';
          else
          cVar2S19S77P069P060P032nsss(0) <='0';
          end if;
        if(cVar1S21S77P035P052P012N029(0)='1' AND  E( 2)='0' AND D( 8)='1' )then
          cVar2S21S77P060P067nsss(0) <='1';
          else
          cVar2S21S77P060P067nsss(0) <='0';
          end if;
        if(cVar1S22S77P035P052P012N029(0)='1' AND  E( 2)='0' AND D( 8)='0' AND B( 5)='1' )then
          cVar2S22S77P060N067P027nsss(0) <='1';
          else
          cVar2S22S77P060N067P027nsss(0) <='0';
          end if;
        if(cVar1S24S77P035N052P046P033(0)='1' AND  A( 0)='0' )then
          cVar2S24S77P019nsss(0) <='1';
          else
          cVar2S24S77P019nsss(0) <='0';
          end if;
        if(cVar1S25S77P035N052P046P033(0)='1' AND  A( 0)='1' AND A(11)='1' )then
          cVar2S25S77P019P016nsss(0) <='1';
          else
          cVar2S25S77P019P016nsss(0) <='0';
          end if;
        if(cVar1S26S77P035N052N046P051(0)='1' AND  B( 0)='1' )then
          cVar2S26S77P037nsss(0) <='1';
          else
          cVar2S26S77P037nsss(0) <='0';
          end if;
        if(cVar1S27S77P035N052N046P051(0)='1' AND  B( 0)='0' AND E(12)='1' )then
          cVar2S27S77N037P053nsss(0) <='1';
          else
          cVar2S27S77N037P053nsss(0) <='0';
          end if;
        if(cVar1S28S77P035N052N046N051(0)='1' AND  A( 6)='0' AND A(16)='0' AND E( 1)='0' )then
          cVar2S28S77P007P006P064nsss(0) <='1';
          else
          cVar2S28S77P007P006P064nsss(0) <='0';
          end if;
        if(cVar1S29S77P035N052N046N051(0)='1' AND  A( 6)='0' AND A(16)='1' AND E(14)='1' )then
          cVar2S29S77P007P006P045nsss(0) <='1';
          else
          cVar2S29S77P007P006P045nsss(0) <='0';
          end if;
        if(cVar1S30S77P035N052N046N051(0)='1' AND  A( 6)='1' AND E(11)='0' AND D(13)='1' )then
          cVar2S30S77P007P057P047nsss(0) <='1';
          else
          cVar2S30S77P007P057P047nsss(0) <='0';
          end if;
        if(cVar1S1S78P035P064P052N036(0)='1' AND  A( 2)='1' )then
          cVar2S1S78P015nsss(0) <='1';
          else
          cVar2S1S78P015nsss(0) <='0';
          end if;
        if(cVar1S2S78P035P064P052N036(0)='1' AND  A( 2)='0' AND B( 4)='1' )then
          cVar2S2S78N015P029nsss(0) <='1';
          else
          cVar2S2S78N015P029nsss(0) <='0';
          end if;
        if(cVar1S3S78P035P064P052N036(0)='1' AND  A( 2)='0' AND B( 4)='0' AND A( 1)='1' )then
          cVar2S3S78N015N029P017nsss(0) <='1';
          else
          cVar2S3S78N015N029P017nsss(0) <='0';
          end if;
        if(cVar1S4S78P035P064N052P037(0)='1' AND  B(10)='0' AND D( 8)='0' )then
          cVar2S4S78P034P067nsss(0) <='1';
          else
          cVar2S4S78P034P067nsss(0) <='0';
          end if;
        if(cVar1S5S78P035P064N052P037(0)='1' AND  B(10)='0' AND D( 8)='1' AND A( 0)='0' )then
          cVar2S5S78P034P067P019nsss(0) <='1';
          else
          cVar2S5S78P034P067P019nsss(0) <='0';
          end if;
        if(cVar1S6S78P035P064N052P037(0)='1' AND  B(10)='1' AND A(13)='1' )then
          cVar2S6S78P034P012nsss(0) <='1';
          else
          cVar2S6S78P034P012nsss(0) <='0';
          end if;
        if(cVar1S7S78P035P064N052P037(0)='1' AND  B(10)='1' AND A(13)='0' AND A( 3)='1' )then
          cVar2S7S78P034N012P013nsss(0) <='1';
          else
          cVar2S7S78P034N012P013nsss(0) <='0';
          end if;
        if(cVar1S8S78P035P064N052N037(0)='1' AND  D( 1)='1' AND B(17)='1' )then
          cVar2S8S78P062P020nsss(0) <='1';
          else
          cVar2S8S78P062P020nsss(0) <='0';
          end if;
        if(cVar1S9S78P035P064N052N037(0)='1' AND  D( 1)='1' AND B(17)='0' AND A( 9)='1' )then
          cVar2S9S78P062N020P001nsss(0) <='1';
          else
          cVar2S9S78P062N020P001nsss(0) <='0';
          end if;
        if(cVar1S10S78P035P064N052N037(0)='1' AND  D( 1)='0' AND E( 0)='1' )then
          cVar2S10S78N062P068nsss(0) <='1';
          else
          cVar2S10S78N062P068nsss(0) <='0';
          end if;
        if(cVar1S11S78P035N064P012P001(0)='1' AND  A( 3)='0' AND B( 3)='0' )then
          cVar2S11S78P013P031nsss(0) <='1';
          else
          cVar2S11S78P013P031nsss(0) <='0';
          end if;
        if(cVar1S12S78P035N064P012P001(0)='1' AND  A( 3)='1' AND A( 2)='0' AND A( 0)='0' )then
          cVar2S12S78P013P015P019nsss(0) <='1';
          else
          cVar2S12S78P013P015P019nsss(0) <='0';
          end if;
        if(cVar1S13S78P035N064P012P001(0)='1' AND  A( 3)='1' AND A( 2)='1' AND D( 9)='1' )then
          cVar2S13S78P013P015P063nsss(0) <='1';
          else
          cVar2S13S78P013P015P063nsss(0) <='0';
          end if;
        if(cVar1S14S78P035N064P012P036(0)='1' AND  B(14)='0' AND A( 5)='0' AND E( 8)='1' )then
          cVar2S14S78P026P009P069nsss(0) <='1';
          else
          cVar2S14S78P026P009P069nsss(0) <='0';
          end if;
        if(cVar1S15S78P035N064P012P036(0)='1' AND  B(14)='0' AND A( 5)='1' AND D( 8)='0' )then
          cVar2S15S78P026P009P067nsss(0) <='1';
          else
          cVar2S15S78P026P009P067nsss(0) <='0';
          end if;
        if(cVar1S16S78P035N064P012N036(0)='1' AND  E( 3)='1' AND D( 3)='1' )then
          cVar2S16S78P056P054nsss(0) <='1';
          else
          cVar2S16S78P056P054nsss(0) <='0';
          end if;
        if(cVar1S17S78N035P016P064P015(0)='1' AND  A(10)='0' AND A( 6)='0' AND E(13)='0' )then
          cVar2S17S78P018P007P049nsss(0) <='1';
          else
          cVar2S17S78P018P007P049nsss(0) <='0';
          end if;
        if(cVar1S18S78N035P016P064P015(0)='1' AND  A(10)='1' AND D( 9)='0' AND A( 4)='1' )then
          cVar2S18S78P018P063P011nsss(0) <='1';
          else
          cVar2S18S78P018P063P011nsss(0) <='0';
          end if;
        if(cVar1S19S78N035P016P064N015(0)='1' AND  A( 1)='1' AND E( 3)='1' AND E( 2)='0' )then
          cVar2S19S78P017P056P060nsss(0) <='1';
          else
          cVar2S19S78P017P056P060nsss(0) <='0';
          end if;
        if(cVar1S20S78N035P016P064N015(0)='1' AND  A( 1)='1' AND E( 3)='0' AND A(16)='1' )then
          cVar2S20S78P017N056P006nsss(0) <='1';
          else
          cVar2S20S78P017N056P006nsss(0) <='0';
          end if;
        if(cVar1S21S78N035P016P064N015(0)='1' AND  A( 1)='0' AND E( 9)='0' AND B(17)='1' )then
          cVar2S21S78N017P065P020nsss(0) <='1';
          else
          cVar2S21S78N017P065P020nsss(0) <='0';
          end if;
        if(cVar1S22S78N035P016P064P048(0)='1' AND  D(12)='0' AND E(11)='1' AND E( 2)='0' )then
          cVar2S22S78P051P057P060nsss(0) <='1';
          else
          cVar2S22S78P051P057P060nsss(0) <='0';
          end if;
        if(cVar1S23S78N035P016P064P048(0)='1' AND  D(12)='0' AND E(11)='0' AND E( 7)='1' )then
          cVar2S23S78P051N057P040nsss(0) <='1';
          else
          cVar2S23S78P051N057P040nsss(0) <='0';
          end if;
        if(cVar1S24S78N035P016P064P048(0)='1' AND  D(12)='1' AND B(14)='1' )then
          cVar2S24S78P051P026nsss(0) <='1';
          else
          cVar2S24S78P051P026nsss(0) <='0';
          end if;
        if(cVar1S25S78N035P016P064P048(0)='1' AND  D( 2)='0' AND A(15)='1' )then
          cVar2S25S78P058P008nsss(0) <='1';
          else
          cVar2S25S78P058P008nsss(0) <='0';
          end if;
        if(cVar1S26S78N035P016P053P004(0)='1' AND  B(13)='1' AND A( 4)='1' )then
          cVar2S26S78P028P011nsss(0) <='1';
          else
          cVar2S26S78P028P011nsss(0) <='0';
          end if;
        if(cVar1S27S78N035P016P053P004(0)='1' AND  B(13)='1' AND A( 4)='0' AND B( 0)='0' )then
          cVar2S27S78P028N011P037nsss(0) <='1';
          else
          cVar2S27S78P028N011P037nsss(0) <='0';
          end if;
        if(cVar1S28S78N035P016P053P004(0)='1' AND  B(13)='0' AND D(13)='0' AND A(19)='0' )then
          cVar2S28S78N028P047P000nsss(0) <='1';
          else
          cVar2S28S78N028P047P000nsss(0) <='0';
          end if;
        if(cVar1S29S78N035P016N053P028(0)='1' AND  A(12)='1' AND A( 0)='1' AND D(10)='0' )then
          cVar2S29S78P014P019P059nsss(0) <='1';
          else
          cVar2S29S78P014P019P059nsss(0) <='0';
          end if;
        if(cVar1S30S78N035P016N053P028(0)='1' AND  A(12)='1' AND A( 0)='0' AND E(10)='1' )then
          cVar2S30S78P014N019P061nsss(0) <='1';
          else
          cVar2S30S78P014N019P061nsss(0) <='0';
          end if;
        if(cVar1S31S78N035P016N053P028(0)='1' AND  A(12)='0' AND E(14)='1' AND E( 1)='1' )then
          cVar2S31S78N014P045P064nsss(0) <='1';
          else
          cVar2S31S78N014P045P064nsss(0) <='0';
          end if;
        if(cVar1S32S78N035P016N053P028(0)='1' AND  A(12)='0' AND E(14)='0' AND E(11)='1' )then
          cVar2S32S78N014N045P057nsss(0) <='1';
          else
          cVar2S32S78N014N045P057nsss(0) <='0';
          end if;
        if(cVar1S33S78N035P016N053P028(0)='1' AND  A( 3)='0' AND E( 9)='0' AND E( 8)='1' )then
          cVar2S33S78P013P065P069nsss(0) <='1';
          else
          cVar2S33S78P013P065P069nsss(0) <='0';
          end if;
        if(cVar1S1S79P064P035N052P055(0)='1' AND  D( 5)='1' AND A( 0)='0' )then
          cVar2S1S79P046P019nsss(0) <='1';
          else
          cVar2S1S79P046P019nsss(0) <='0';
          end if;
        if(cVar1S2S79P064P035N052P055(0)='1' AND  D( 5)='0' AND E(11)='1' AND D(10)='1' )then
          cVar2S2S79N046P057P059nsss(0) <='1';
          else
          cVar2S2S79N046P057P059nsss(0) <='0';
          end if;
        if(cVar1S3S79P064P035N052P055(0)='1' AND  D( 5)='0' AND E(11)='0' )then
          cVar2S3S79N046N057psss(0) <='1';
          else
          cVar2S3S79N046N057psss(0) <='0';
          end if;
        if(cVar1S4S79P064P035N052P055(0)='1' AND  E( 3)='1' )then
          cVar2S4S79P056nsss(0) <='1';
          else
          cVar2S4S79P056nsss(0) <='0';
          end if;
        if(cVar1S5S79P064P035N052P055(0)='1' AND  E( 3)='0' AND A( 3)='1' AND A(11)='0' )then
          cVar2S5S79N056P013P016nsss(0) <='1';
          else
          cVar2S5S79N056P013P016nsss(0) <='0';
          end if;
        if(cVar1S6S79P064N035P051P048(0)='1' AND  A( 5)='1' )then
          cVar2S6S79P009nsss(0) <='1';
          else
          cVar2S6S79P009nsss(0) <='0';
          end if;
        if(cVar1S7S79P064N035P051P048(0)='1' AND  A( 5)='0' AND D( 4)='0' )then
          cVar2S7S79N009P050nsss(0) <='1';
          else
          cVar2S7S79N009P050nsss(0) <='0';
          end if;
        if(cVar1S8S79P064N035P051P048(0)='1' AND  A( 5)='0' AND D( 4)='1' AND A(15)='1' )then
          cVar2S8S79N009P050P008nsss(0) <='1';
          else
          cVar2S8S79N009P050P008nsss(0) <='0';
          end if;
        if(cVar1S9S79P064N035P051P048(0)='1' AND  D( 2)='0' AND B(10)='0' AND A( 1)='0' )then
          cVar2S9S79P058P034P017nsss(0) <='1';
          else
          cVar2S9S79P058P034P017nsss(0) <='0';
          end if;
        if(cVar1S10S79P064N035P051P069(0)='1' AND  A( 0)='0' AND B(14)='1' )then
          cVar2S10S79P019P026nsss(0) <='1';
          else
          cVar2S10S79P019P026nsss(0) <='0';
          end if;
        if(cVar1S11S79N064P035P016P026(0)='1' AND  D( 4)='1' )then
          cVar2S11S79P050nsss(0) <='1';
          else
          cVar2S11S79P050nsss(0) <='0';
          end if;
        if(cVar1S12S79N064P035P016P026(0)='1' AND  D( 4)='0' AND B( 4)='0' AND E( 6)='0' )then
          cVar2S12S79N050P029P044nsss(0) <='1';
          else
          cVar2S12S79N050P029P044nsss(0) <='0';
          end if;
        if(cVar1S13S79N064P035P016N026(0)='1' AND  A( 2)='0' AND A( 8)='0' )then
          cVar2S13S79P015P003nsss(0) <='1';
          else
          cVar2S13S79P015P003nsss(0) <='0';
          end if;
        if(cVar1S14S79N064P035P016N026(0)='1' AND  A( 2)='0' AND A( 8)='1' AND E(14)='1' )then
          cVar2S14S79P015P003P045nsss(0) <='1';
          else
          cVar2S14S79P015P003P045nsss(0) <='0';
          end if;
        if(cVar1S15S79N064P035P016N026(0)='1' AND  A( 2)='1' AND D(11)='1' AND B( 2)='0' )then
          cVar2S15S79P015P055P033nsss(0) <='1';
          else
          cVar2S15S79P015P055P033nsss(0) <='0';
          end if;
        if(cVar1S16S79N064P035P016N026(0)='1' AND  A( 2)='1' AND D(11)='0' AND D( 2)='1' )then
          cVar2S16S79P015N055P058nsss(0) <='1';
          else
          cVar2S16S79P015N055P058nsss(0) <='0';
          end if;
        if(cVar1S17S79N064P035P016P052(0)='1' AND  B( 4)='1' )then
          cVar2S17S79P029nsss(0) <='1';
          else
          cVar2S17S79P029nsss(0) <='0';
          end if;
        if(cVar1S18S79N064P035P016P052(0)='1' AND  B( 4)='0' AND B( 5)='1' )then
          cVar2S18S79N029P027nsss(0) <='1';
          else
          cVar2S18S79N029P027nsss(0) <='0';
          end if;
        if(cVar1S19S79N064P035P016P052(0)='1' AND  B( 4)='0' AND B( 5)='0' AND B(13)='1' )then
          cVar2S19S79N029N027P028nsss(0) <='1';
          else
          cVar2S19S79N029N027P028nsss(0) <='0';
          end if;
        if(cVar1S20S79N064P035P016N052(0)='1' AND  E( 9)='1' AND E( 8)='0' AND E( 2)='0' )then
          cVar2S20S79P065P069P060nsss(0) <='1';
          else
          cVar2S20S79P065P069P060nsss(0) <='0';
          end if;
        if(cVar1S21S79N064P035P016N052(0)='1' AND  E( 9)='0' AND B( 0)='1' AND D( 9)='0' )then
          cVar2S21S79N065P037P063nsss(0) <='1';
          else
          cVar2S21S79N065P037P063nsss(0) <='0';
          end if;
        if(cVar1S22S79N064P035P013P016(0)='1' AND  B( 4)='0' AND A( 1)='0' AND A(14)='0' )then
          cVar2S22S79P029P017P010nsss(0) <='1';
          else
          cVar2S22S79P029P017P010nsss(0) <='0';
          end if;
        if(cVar1S23S79N064P035P013N016(0)='1' AND  B(11)='0' AND D(10)='1' AND A(12)='1' )then
          cVar2S23S79P032P059P014nsss(0) <='1';
          else
          cVar2S23S79P032P059P014nsss(0) <='0';
          end if;
        if(cVar1S24S79N064P035P013N016(0)='1' AND  B(11)='1' AND D(10)='0' AND E( 2)='1' )then
          cVar2S24S79P032P059P060nsss(0) <='1';
          else
          cVar2S24S79P032P059P060nsss(0) <='0';
          end if;
        if(cVar1S25S79N064P035P013N016(0)='1' AND  B(11)='1' AND D(10)='1' AND D( 9)='1' )then
          cVar2S25S79P032P059P063nsss(0) <='1';
          else
          cVar2S25S79P032P059P063nsss(0) <='0';
          end if;
        if(cVar1S26S79N064P035P013P030(0)='1' AND  E(11)='1' )then
          cVar2S26S79P057nsss(0) <='1';
          else
          cVar2S26S79P057nsss(0) <='0';
          end if;
        if(cVar1S27S79N064P035P013P030(0)='1' AND  E(11)='0' AND A(13)='1' )then
          cVar2S27S79N057P012nsss(0) <='1';
          else
          cVar2S27S79N057P012nsss(0) <='0';
          end if;
        if(cVar1S28S79N064P035P013N030(0)='1' AND  A( 2)='0' AND D(10)='0' AND E( 0)='0' )then
          cVar2S28S79P015P059P068nsss(0) <='1';
          else
          cVar2S28S79P015P059P068nsss(0) <='0';
          end if;
        if(cVar1S29S79N064P035P013N030(0)='1' AND  A( 2)='1' AND D( 9)='1' AND A(11)='0' )then
          cVar2S29S79P015P063P016nsss(0) <='1';
          else
          cVar2S29S79P015P063P016nsss(0) <='0';
          end if;
        if(cVar1S0S80P037P034P057P058(0)='1' AND  B(11)='0' AND A(14)='0' )then
          cVar2S0S80P032P010nsss(0) <='1';
          else
          cVar2S0S80P032P010nsss(0) <='0';
          end if;
        if(cVar1S1S80P037P034P057P058(0)='1' AND  B(11)='0' AND A(14)='1' AND B( 5)='1' )then
          cVar2S1S80P032P010P027nsss(0) <='1';
          else
          cVar2S1S80P032P010P027nsss(0) <='0';
          end if;
        if(cVar1S2S80P037P034P057P058(0)='1' AND  B(11)='1' AND E(10)='1' AND A(12)='1' )then
          cVar2S2S80P032P061P014nsss(0) <='1';
          else
          cVar2S2S80P032P061P014nsss(0) <='0';
          end if;
        if(cVar1S3S80P037P034P057P058(0)='1' AND  A(12)='0' AND B( 3)='1' )then
          cVar2S3S80P014P031nsss(0) <='1';
          else
          cVar2S3S80P014P031nsss(0) <='0';
          end if;
        if(cVar1S4S80P037P034P057P058(0)='1' AND  A(12)='0' AND B( 3)='0' AND A( 5)='1' )then
          cVar2S4S80P014N031P009nsss(0) <='1';
          else
          cVar2S4S80P014N031P009nsss(0) <='0';
          end if;
        if(cVar1S5S80P037P034P057P058(0)='1' AND  A(12)='1' AND B( 3)='0' AND A( 2)='0' )then
          cVar2S5S80P014P031P015nsss(0) <='1';
          else
          cVar2S5S80P014P031P015nsss(0) <='0';
          end if;
        if(cVar1S6S80P037P034P057P014(0)='1' AND  A(11)='1' )then
          cVar2S6S80P016nsss(0) <='1';
          else
          cVar2S6S80P016nsss(0) <='0';
          end if;
        if(cVar1S7S80P037P034P057P014(0)='1' AND  A(11)='0' AND B(12)='1' )then
          cVar2S7S80N016P030nsss(0) <='1';
          else
          cVar2S7S80N016P030nsss(0) <='0';
          end if;
        if(cVar1S8S80P037P034P057N014(0)='1' AND  A(13)='0' AND B( 1)='1' )then
          cVar2S8S80P012P035nsss(0) <='1';
          else
          cVar2S8S80P012P035nsss(0) <='0';
          end if;
        if(cVar1S9S80P037N034P017P012(0)='1' AND  E( 6)='1' )then
          cVar2S9S80P044nsss(0) <='1';
          else
          cVar2S9S80P044nsss(0) <='0';
          end if;
        if(cVar1S10S80P037N034P017P012(0)='1' AND  E( 6)='0' AND A( 4)='0' )then
          cVar2S10S80N044P011nsss(0) <='1';
          else
          cVar2S10S80N044P011nsss(0) <='0';
          end if;
        if(cVar1S11S80P037N034P017P012(0)='1' AND  E( 6)='0' AND A( 4)='1' AND D( 2)='1' )then
          cVar2S11S80N044P011P058nsss(0) <='1';
          else
          cVar2S11S80N044P011P058nsss(0) <='0';
          end if;
        if(cVar1S12S80P037N034P017P012(0)='1' AND  B( 3)='1' AND D( 1)='0' )then
          cVar2S12S80P031P062nsss(0) <='1';
          else
          cVar2S12S80P031P062nsss(0) <='0';
          end if;
        if(cVar1S13S80P037N034P017P012(0)='1' AND  B( 3)='0' AND B(11)='1' AND A( 5)='0' )then
          cVar2S13S80N031P032P009nsss(0) <='1';
          else
          cVar2S13S80N031P032P009nsss(0) <='0';
          end if;
        if(cVar1S14S80P037N034N017P012(0)='1' AND  E(10)='0' AND A( 3)='0' )then
          cVar2S14S80P061P013nsss(0) <='1';
          else
          cVar2S14S80P061P013nsss(0) <='0';
          end if;
        if(cVar1S15S80P037N034N017P012(0)='1' AND  E(10)='1' AND B( 3)='0' AND D( 2)='0' )then
          cVar2S15S80P061P031P058nsss(0) <='1';
          else
          cVar2S15S80P061P031P058nsss(0) <='0';
          end if;
        if(cVar1S16S80P037N034N017P012(0)='1' AND  E(10)='1' AND B( 3)='1' AND A( 3)='1' )then
          cVar2S16S80P061P031P013nsss(0) <='1';
          else
          cVar2S16S80P061P031P013nsss(0) <='0';
          end if;
        if(cVar1S17S80P037N034N017N012(0)='1' AND  B(11)='1' AND A( 7)='0' )then
          cVar2S17S80P032P005nsss(0) <='1';
          else
          cVar2S17S80P032P005nsss(0) <='0';
          end if;
        if(cVar1S18S80P037N034N017N012(0)='1' AND  B(11)='0' AND D( 2)='0' AND B( 3)='1' )then
          cVar2S18S80N032P058P031nsss(0) <='1';
          else
          cVar2S18S80N032P058P031nsss(0) <='0';
          end if;
        if(cVar1S19S80P037N034N017N012(0)='1' AND  B(11)='0' AND D( 2)='1' AND A(11)='1' )then
          cVar2S19S80N032P058P016nsss(0) <='1';
          else
          cVar2S19S80N032P058P016nsss(0) <='0';
          end if;
        if(cVar1S21S80P037P015P052N029(0)='1' AND  A(10)='0' AND A(11)='0' )then
          cVar2S21S80P018P016nsss(0) <='1';
          else
          cVar2S21S80P018P016nsss(0) <='0';
          end if;
        if(cVar1S22S80P037P015N052P025(0)='1' AND  A(11)='0' AND E( 0)='1' )then
          cVar2S22S80P016P068nsss(0) <='1';
          else
          cVar2S22S80P016P068nsss(0) <='0';
          end if;
        if(cVar1S23S80P037P015N052P025(0)='1' AND  A(11)='0' AND E( 0)='0' AND A(10)='1' )then
          cVar2S23S80P016N068P018nsss(0) <='1';
          else
          cVar2S23S80P016N068P018nsss(0) <='0';
          end if;
        if(cVar1S24S80P037P015N052N025(0)='1' AND  B(14)='0' AND D(13)='0' AND B(15)='0' )then
          cVar2S24S80P026P047P024nsss(0) <='1';
          else
          cVar2S24S80P026P047P024nsss(0) <='0';
          end if;
        if(cVar1S25S80P037P015N052N025(0)='1' AND  B(14)='1' AND E(12)='0' AND E( 0)='1' )then
          cVar2S25S80P026P053P068nsss(0) <='1';
          else
          cVar2S25S80P026P053P068nsss(0) <='0';
          end if;
        if(cVar1S26S80P037N015P018P055(0)='1' AND  B(10)='1' AND B( 1)='0' )then
          cVar2S26S80P034P035nsss(0) <='1';
          else
          cVar2S26S80P034P035nsss(0) <='0';
          end if;
        if(cVar1S27S80P037N015P018P055(0)='1' AND  B(10)='1' AND B( 1)='1' AND A( 1)='0' )then
          cVar2S27S80P034P035P017nsss(0) <='1';
          else
          cVar2S27S80P034P035P017nsss(0) <='0';
          end if;
        if(cVar1S28S80P037N015P018P055(0)='1' AND  B(10)='0' AND D( 1)='0' AND E(10)='0' )then
          cVar2S28S80N034P062P061nsss(0) <='1';
          else
          cVar2S28S80N034P062P061nsss(0) <='0';
          end if;
        if(cVar1S29S80P037N015P018P055(0)='1' AND  B(10)='0' AND D( 1)='1' AND D(10)='1' )then
          cVar2S29S80N034P062P059nsss(0) <='1';
          else
          cVar2S29S80N034P062P059nsss(0) <='0';
          end if;
        if(cVar1S30S80P037N015P018P055(0)='1' AND  E(12)='0' AND D( 1)='1' )then
          cVar2S30S80P053P062nsss(0) <='1';
          else
          cVar2S30S80P053P062nsss(0) <='0';
          end if;
        if(cVar1S31S80P037N015N018P034(0)='1' AND  E( 7)='1' AND D( 1)='1' )then
          cVar2S31S80P040P062nsss(0) <='1';
          else
          cVar2S31S80P040P062nsss(0) <='0';
          end if;
        if(cVar1S32S80P037N015N018P034(0)='1' AND  E( 7)='1' AND D( 1)='0' AND D( 7)='1' )then
          cVar2S32S80P040N062P038nsss(0) <='1';
          else
          cVar2S32S80P040N062P038nsss(0) <='0';
          end if;
        if(cVar1S33S80P037N015N018P034(0)='1' AND  E( 7)='0' AND D(11)='1' AND A(15)='0' )then
          cVar2S33S80N040P055P008nsss(0) <='1';
          else
          cVar2S33S80N040P055P008nsss(0) <='0';
          end if;
        if(cVar1S34S80P037N015N018P034(0)='1' AND  E( 7)='0' AND D(11)='0' AND B( 1)='1' )then
          cVar2S34S80N040N055P035nsss(0) <='1';
          else
          cVar2S34S80N040N055P035nsss(0) <='0';
          end if;
        if(cVar1S35S80P037N015N018P034(0)='1' AND  E( 2)='1' AND E( 8)='1' )then
          cVar2S35S80P060P069nsss(0) <='1';
          else
          cVar2S35S80P060P069nsss(0) <='0';
          end if;
        if(cVar1S36S80P037N015N018P034(0)='1' AND  E( 2)='1' AND E( 8)='0' AND A( 0)='1' )then
          cVar2S36S80P060N069P019nsss(0) <='1';
          else
          cVar2S36S80P060N069P019nsss(0) <='0';
          end if;
        if(cVar1S37S80P037N015N018P034(0)='1' AND  E( 2)='0' AND B(12)='1' )then
          cVar2S37S80N060P030nsss(0) <='1';
          else
          cVar2S37S80N060P030nsss(0) <='0';
          end if;
        if(cVar1S0S81P037P032P017P056(0)='1' AND  B( 4)='1' AND B(12)='0' AND E( 4)='1' )then
          cVar2S0S81P029P030P052nsss(0) <='1';
          else
          cVar2S0S81P029P030P052nsss(0) <='0';
          end if;
        if(cVar1S1S81P037P032P017P056(0)='1' AND  B( 4)='0' AND D( 3)='0' )then
          cVar2S1S81N029P054nsss(0) <='1';
          else
          cVar2S1S81N029P054nsss(0) <='0';
          end if;
        if(cVar1S2S81P037P032P017P056(0)='1' AND  B( 4)='0' AND D( 3)='1' AND B(13)='1' )then
          cVar2S2S81N029P054P028nsss(0) <='1';
          else
          cVar2S2S81N029P054P028nsss(0) <='0';
          end if;
        if(cVar1S3S81P037P032P017P056(0)='1' AND  A( 3)='1' AND E( 9)='0' AND B(13)='0' )then
          cVar2S3S81P013P065P028nsss(0) <='1';
          else
          cVar2S3S81P013P065P028nsss(0) <='0';
          end if;
        if(cVar1S4S81P037P032P017P056(0)='1' AND  A( 3)='0' AND E( 4)='0' AND A(12)='1' )then
          cVar2S4S81N013P052P014nsss(0) <='1';
          else
          cVar2S4S81N013P052P014nsss(0) <='0';
          end if;
        if(cVar1S5S81P037P032P017P056(0)='1' AND  A( 3)='0' AND E( 4)='1' AND A( 5)='1' )then
          cVar2S5S81N013P052P009nsss(0) <='1';
          else
          cVar2S5S81N013P052P009nsss(0) <='0';
          end if;
        if(cVar1S6S81P037P032P017P036(0)='1' AND  E( 8)='1' AND E(10)='0' AND A(10)='1' )then
          cVar2S6S81P069P061P018nsss(0) <='1';
          else
          cVar2S6S81P069P061P018nsss(0) <='0';
          end if;
        if(cVar1S7S81P037P032P017P036(0)='1' AND  E( 8)='0' AND D( 1)='1' AND A(12)='0' )then
          cVar2S7S81N069P062P014nsss(0) <='1';
          else
          cVar2S7S81N069P062P014nsss(0) <='0';
          end if;
        if(cVar1S8S81P037P032P017N036(0)='1' AND  E( 8)='0' AND B(14)='1' AND B( 3)='0' )then
          cVar2S8S81P069P026P031nsss(0) <='1';
          else
          cVar2S8S81P069P026P031nsss(0) <='0';
          end if;
        if(cVar1S9S81P037P032P017N036(0)='1' AND  E( 8)='1' AND B( 4)='1' )then
          cVar2S9S81P069P029nsss(0) <='1';
          else
          cVar2S9S81P069P029nsss(0) <='0';
          end if;
        if(cVar1S10S81P037P032P013P031(0)='1' AND  B( 5)='0' AND E(14)='0' AND A(12)='0' )then
          cVar2S10S81P027P045P014nsss(0) <='1';
          else
          cVar2S10S81P027P045P014nsss(0) <='0';
          end if;
        if(cVar1S11S81P037P032P013P031(0)='1' AND  B( 5)='0' AND E(14)='1' AND D(14)='1' )then
          cVar2S11S81P027P045P043nsss(0) <='1';
          else
          cVar2S11S81P027P045P043nsss(0) <='0';
          end if;
        if(cVar1S12S81P037P032P013P031(0)='1' AND  A(14)='1' )then
          cVar2S12S81P010nsss(0) <='1';
          else
          cVar2S12S81P010nsss(0) <='0';
          end if;
        if(cVar1S13S81P037P032P013P031(0)='1' AND  A(14)='0' AND A( 0)='1' )then
          cVar2S13S81N010P019nsss(0) <='1';
          else
          cVar2S13S81N010P019nsss(0) <='0';
          end if;
        if(cVar1S14S81P037P032P013P059(0)='1' AND  B(12)='1' )then
          cVar2S14S81P030nsss(0) <='1';
          else
          cVar2S14S81P030nsss(0) <='0';
          end if;
        if(cVar1S15S81P037P032P013P059(0)='1' AND  B(12)='0' AND A( 2)='0' AND B( 9)='0' )then
          cVar2S15S81N030P015P036nsss(0) <='1';
          else
          cVar2S15S81N030P015P036nsss(0) <='0';
          end if;
        if(cVar1S16S81P037P032P013P059(0)='1' AND  B(12)='0' AND A( 2)='1' AND A( 0)='1' )then
          cVar2S16S81N030P015P019nsss(0) <='1';
          else
          cVar2S16S81N030P015P019nsss(0) <='0';
          end if;
        if(cVar1S17S81P037P032P013N059(0)='1' AND  A(13)='0' AND D( 2)='1' )then
          cVar2S17S81P012P058nsss(0) <='1';
          else
          cVar2S17S81P012P058nsss(0) <='0';
          end if;
        if(cVar1S18S81P037P032P013N059(0)='1' AND  A(13)='0' AND D( 2)='0' AND E( 9)='1' )then
          cVar2S18S81P012N058P065nsss(0) <='1';
          else
          cVar2S18S81P012N058P065nsss(0) <='0';
          end if;
        if(cVar1S20S81P037P052P008N013(0)='1' AND  B( 5)='1' )then
          cVar2S20S81P027nsss(0) <='1';
          else
          cVar2S20S81P027nsss(0) <='0';
          end if;
        if(cVar1S21S81P037P052P008N013(0)='1' AND  B( 5)='0' AND A( 1)='1' )then
          cVar2S21S81N027P017nsss(0) <='1';
          else
          cVar2S21S81N027P017nsss(0) <='0';
          end if;
        if(cVar1S22S81P037P052P008N013(0)='1' AND  B( 5)='0' AND A( 1)='0' AND E( 0)='0' )then
          cVar2S22S81N027N017P068nsss(0) <='1';
          else
          cVar2S22S81N027N017P068nsss(0) <='0';
          end if;
        if(cVar1S23S81P037P052N008P068(0)='1' AND  A( 1)='1' )then
          cVar2S23S81P017nsss(0) <='1';
          else
          cVar2S23S81P017nsss(0) <='0';
          end if;
        if(cVar1S24S81P037P052N008P068(0)='1' AND  A( 1)='0' AND D( 8)='1' )then
          cVar2S24S81N017P067nsss(0) <='1';
          else
          cVar2S24S81N017P067nsss(0) <='0';
          end if;
        if(cVar1S25S81P037P052N008P068(0)='1' AND  A( 1)='0' AND D( 8)='0' AND A(14)='1' )then
          cVar2S25S81N017N067P010nsss(0) <='1';
          else
          cVar2S25S81N017N067P010nsss(0) <='0';
          end if;
        if(cVar1S26S81P037P052N008N068(0)='1' AND  B( 2)='1' )then
          cVar2S26S81P033nsss(0) <='1';
          else
          cVar2S26S81P033nsss(0) <='0';
          end if;
        if(cVar1S27S81P037P052N008N068(0)='1' AND  B( 2)='0' AND E( 9)='1' )then
          cVar2S27S81N033P065nsss(0) <='1';
          else
          cVar2S27S81N033P065nsss(0) <='0';
          end if;
        if(cVar1S28S81P037P052N008N068(0)='1' AND  B( 2)='0' AND E( 9)='0' AND A( 4)='1' )then
          cVar2S28S81N033N065P011nsss(0) <='1';
          else
          cVar2S28S81N033N065P011nsss(0) <='0';
          end if;
        if(cVar1S30S81P037N052P025N044(0)='1' AND  B( 9)='1' AND A(11)='0' )then
          cVar2S30S81P036P016nsss(0) <='1';
          else
          cVar2S30S81P036P016nsss(0) <='0';
          end if;
        if(cVar1S31S81P037N052P025N044(0)='1' AND  B( 9)='0' AND D( 1)='1' AND D( 0)='1' )then
          cVar2S31S81N036P062P066nsss(0) <='1';
          else
          cVar2S31S81N036P062P066nsss(0) <='0';
          end if;
        if(cVar1S32S81P037N052N025P024(0)='1' AND  B( 8)='1' )then
          cVar2S32S81P021nsss(0) <='1';
          else
          cVar2S32S81P021nsss(0) <='0';
          end if;
        if(cVar1S33S81P037N052N025P024(0)='1' AND  B( 8)='0' AND D( 0)='0' )then
          cVar2S33S81N021P066nsss(0) <='1';
          else
          cVar2S33S81N021P066nsss(0) <='0';
          end if;
        if(cVar1S34S81P037N052N025P024(0)='1' AND  B( 8)='0' AND D( 0)='1' AND A( 7)='1' )then
          cVar2S34S81N021P066P005nsss(0) <='1';
          else
          cVar2S34S81N021P066P005nsss(0) <='0';
          end if;
        if(cVar1S35S81P037N052N025N024(0)='1' AND  D(13)='0' AND A( 6)='0' AND D( 3)='1' )then
          cVar2S35S81P047P007P054nsss(0) <='1';
          else
          cVar2S35S81P047P007P054nsss(0) <='0';
          end if;
        if(cVar1S36S81P037N052N025N024(0)='1' AND  D(13)='0' AND A( 6)='1' AND B(16)='1' )then
          cVar2S36S81P047P007P022nsss(0) <='1';
          else
          cVar2S36S81P047P007P022nsss(0) <='0';
          end if;
        if(cVar1S37S81P037N052N025N024(0)='1' AND  D(13)='1' AND B(14)='1' AND A(15)='0' )then
          cVar2S37S81P047P026P008nsss(0) <='1';
          else
          cVar2S37S81P047P026P008nsss(0) <='0';
          end if;
        if(cVar1S38S81P037N052N025N024(0)='1' AND  D(13)='1' AND B(14)='0' AND A(14)='1' )then
          cVar2S38S81P047N026P010nsss(0) <='1';
          else
          cVar2S38S81P047N026P010nsss(0) <='0';
          end if;
        if(cVar1S0S82P037P031P054P034(0)='1' AND  E( 6)='1' AND A( 6)='0' )then
          cVar2S0S82P044P007nsss(0) <='1';
          else
          cVar2S0S82P044P007nsss(0) <='0';
          end if;
        if(cVar1S1S82P037P031P054P034(0)='1' AND  E( 6)='0' AND D( 8)='0' )then
          cVar2S1S82N044P067nsss(0) <='1';
          else
          cVar2S1S82N044P067nsss(0) <='0';
          end if;
        if(cVar1S2S82P037P031P054P034(0)='1' AND  E( 6)='0' AND D( 8)='1' AND D( 9)='0' )then
          cVar2S2S82N044P067P063nsss(0) <='1';
          else
          cVar2S2S82N044P067P063nsss(0) <='0';
          end if;
        if(cVar1S3S82P037P031P054P034(0)='1' AND  B( 1)='0' AND B( 9)='1' )then
          cVar2S3S82P035P036nsss(0) <='1';
          else
          cVar2S3S82P035P036nsss(0) <='0';
          end if;
        if(cVar1S4S82P037P031P054P034(0)='1' AND  B( 1)='1' AND A( 6)='1' )then
          cVar2S4S82P035P007nsss(0) <='1';
          else
          cVar2S4S82P035P007nsss(0) <='0';
          end if;
        if(cVar1S5S82P037P031P054P034(0)='1' AND  B( 1)='1' AND A( 6)='0' AND A(13)='1' )then
          cVar2S5S82P035N007P012nsss(0) <='1';
          else
          cVar2S5S82P035N007P012nsss(0) <='0';
          end if;
        if(cVar1S6S82P037P031P054P065(0)='1' AND  A(13)='0' )then
          cVar2S6S82P012nsss(0) <='1';
          else
          cVar2S6S82P012nsss(0) <='0';
          end if;
        if(cVar1S7S82P037P031P054N065(0)='1' AND  D( 8)='1' AND B( 4)='1' )then
          cVar2S7S82P067P029nsss(0) <='1';
          else
          cVar2S7S82P067P029nsss(0) <='0';
          end if;
        if(cVar1S8S82P037P031P054N065(0)='1' AND  D( 8)='1' AND B( 4)='0' AND A(13)='1' )then
          cVar2S8S82P067N029P012nsss(0) <='1';
          else
          cVar2S8S82P067N029P012nsss(0) <='0';
          end if;
        if(cVar1S9S82P037P031P054N065(0)='1' AND  D( 8)='0' AND A( 0)='1' AND A(14)='1' )then
          cVar2S9S82N067P019P010nsss(0) <='1';
          else
          cVar2S9S82N067P019P010nsss(0) <='0';
          end if;
        if(cVar1S10S82P037P031P058P007(0)='1' AND  D( 3)='0' )then
          cVar2S10S82P054nsss(0) <='1';
          else
          cVar2S10S82P054nsss(0) <='0';
          end if;
        if(cVar1S11S82P037P031N058P054(0)='1' AND  A(10)='0' AND E( 0)='0' )then
          cVar2S11S82P018P068nsss(0) <='1';
          else
          cVar2S11S82P018P068nsss(0) <='0';
          end if;
        if(cVar1S12S82P037P031N058P054(0)='1' AND  A(10)='0' AND E( 0)='1' AND A(14)='0' )then
          cVar2S12S82P018P068P010nsss(0) <='1';
          else
          cVar2S12S82P018P068P010nsss(0) <='0';
          end if;
        if(cVar1S13S82P037P031N058N054(0)='1' AND  A( 3)='1' AND A( 4)='0' AND E(11)='1' )then
          cVar2S13S82P013P011P057nsss(0) <='1';
          else
          cVar2S13S82P013P011P057nsss(0) <='0';
          end if;
        if(cVar1S14S82N037P017P044P060(0)='1' AND  A(14)='0' )then
          cVar2S14S82P010nsss(0) <='1';
          else
          cVar2S14S82P010nsss(0) <='0';
          end if;
        if(cVar1S15S82N037P017N044P023(0)='1' AND  A( 0)='1' AND D( 6)='0' )then
          cVar2S15S82P019P042nsss(0) <='1';
          else
          cVar2S15S82P019P042nsss(0) <='0';
          end if;
        if(cVar1S16S82N037P017N044P023(0)='1' AND  A( 0)='0' AND E( 8)='0' AND B( 9)='0' )then
          cVar2S16S82N019P069P036nsss(0) <='1';
          else
          cVar2S16S82N019P069P036nsss(0) <='0';
          end if;
        if(cVar1S17S82N037P017N044P023(0)='1' AND  A( 0)='0' AND E( 8)='1' AND A(10)='1' )then
          cVar2S17S82N019P069P018nsss(0) <='1';
          else
          cVar2S17S82N019P069P018nsss(0) <='0';
          end if;
        if(cVar1S18S82N037P017N044P023(0)='1' AND  A( 7)='1' )then
          cVar2S18S82P005nsss(0) <='1';
          else
          cVar2S18S82P005nsss(0) <='0';
          end if;
        if(cVar1S19S82N037P017N044P023(0)='1' AND  A( 7)='0' AND A(12)='1' AND A(10)='1' )then
          cVar2S19S82N005P014P018nsss(0) <='1';
          else
          cVar2S19S82N005P014P018nsss(0) <='0';
          end if;
        if(cVar1S20S82N037N017P029P009(0)='1' AND  D( 8)='0' AND B( 9)='0' )then
          cVar2S20S82P067P036nsss(0) <='1';
          else
          cVar2S20S82P067P036nsss(0) <='0';
          end if;
        if(cVar1S21S82N037N017P029P009(0)='1' AND  D( 8)='1' AND B( 9)='1' )then
          cVar2S21S82P067P036nsss(0) <='1';
          else
          cVar2S21S82P067P036nsss(0) <='0';
          end if;
        if(cVar1S22S82N037N017P029N009(0)='1' AND  E( 3)='0' AND B(12)='0' )then
          cVar2S22S82P056P030nsss(0) <='1';
          else
          cVar2S22S82P056P030nsss(0) <='0';
          end if;
        if(cVar1S23S82N037N017P029N009(0)='1' AND  E( 3)='1' AND E( 4)='0' AND B( 3)='0' )then
          cVar2S23S82P056P052P031nsss(0) <='1';
          else
          cVar2S23S82P056P052P031nsss(0) <='0';
          end if;
        if(cVar1S24S82N037N017N029P067(0)='1' AND  B(14)='1' )then
          cVar2S24S82P026nsss(0) <='1';
          else
          cVar2S24S82P026nsss(0) <='0';
          end if;
        if(cVar1S25S82N037N017N029N067(0)='1' AND  A(19)='0' AND E( 6)='1' AND A(14)='1' )then
          cVar2S25S82P000P044P010nsss(0) <='1';
          else
          cVar2S25S82P000P044P010nsss(0) <='0';
          end if;
        if(cVar1S0S83P017P037P000P047(0)='1' AND  A(16)='1' AND D( 5)='0' )then
          cVar2S0S83P006P046nsss(0) <='1';
          else
          cVar2S0S83P006P046nsss(0) <='0';
          end if;
        if(cVar1S1S83P017P037P000P047(0)='1' AND  A(16)='0' AND E( 2)='1' AND E(13)='1' )then
          cVar2S1S83N006P060P049nsss(0) <='1';
          else
          cVar2S1S83N006P060P049nsss(0) <='0';
          end if;
        if(cVar1S2S83P017P037P000P047(0)='1' AND  A(16)='0' AND E( 2)='0' AND A(10)='1' )then
          cVar2S2S83N006N060P018nsss(0) <='1';
          else
          cVar2S2S83N006N060P018nsss(0) <='0';
          end if;
        if(cVar1S3S83P017P037P000N047(0)='1' AND  B(15)='0' AND E(13)='0' )then
          cVar2S3S83P024P049nsss(0) <='1';
          else
          cVar2S3S83P024P049nsss(0) <='0';
          end if;
        if(cVar1S4S83P017P037P000N047(0)='1' AND  B(15)='0' AND E(13)='1' AND D(12)='1' )then
          cVar2S4S83P024P049P051nsss(0) <='1';
          else
          cVar2S4S83P024P049P051nsss(0) <='0';
          end if;
        if(cVar1S5S83P017P037P000N047(0)='1' AND  B(15)='1' AND A(18)='0' AND B(17)='1' )then
          cVar2S5S83P024P002P020nsss(0) <='1';
          else
          cVar2S5S83P024P002P020nsss(0) <='0';
          end if;
        if(cVar1S7S83P017P037P000N021(0)='1' AND  A( 8)='1' AND E( 8)='1' )then
          cVar2S7S83P003P069nsss(0) <='1';
          else
          cVar2S7S83P003P069nsss(0) <='0';
          end if;
        if(cVar1S8S83P017P037P019P003(0)='1' AND  A( 7)='0' )then
          cVar2S8S83P005nsss(0) <='1';
          else
          cVar2S8S83P005nsss(0) <='0';
          end if;
        if(cVar1S9S83P017P037P019N003(0)='1' AND  B( 4)='1' )then
          cVar2S9S83P029nsss(0) <='1';
          else
          cVar2S9S83P029nsss(0) <='0';
          end if;
        if(cVar1S10S83P017P037P019N003(0)='1' AND  B( 4)='0' AND D( 8)='0' AND E(10)='0' )then
          cVar2S10S83N029P067P061nsss(0) <='1';
          else
          cVar2S10S83N029P067P061nsss(0) <='0';
          end if;
        if(cVar1S11S83P017P037P019N003(0)='1' AND  B( 4)='0' AND D( 8)='1' AND E( 3)='1' )then
          cVar2S11S83N029P067P056nsss(0) <='1';
          else
          cVar2S11S83N029P067P056nsss(0) <='0';
          end if;
        if(cVar1S12S83P017P037N019P001(0)='1' AND  D( 1)='0' AND D( 8)='1' AND A(19)='0' )then
          cVar2S12S83P062P067P000nsss(0) <='1';
          else
          cVar2S12S83P062P067P000nsss(0) <='0';
          end if;
        if(cVar1S13S83P017P037N019P001(0)='1' AND  D( 1)='0' AND D( 8)='0' AND B(10)='1' )then
          cVar2S13S83P062N067P034nsss(0) <='1';
          else
          cVar2S13S83P062N067P034nsss(0) <='0';
          end if;
        if(cVar1S14S83P017P037N019P001(0)='1' AND  D( 1)='1' AND D( 0)='0' AND B(12)='1' )then
          cVar2S14S83P062P066P030nsss(0) <='1';
          else
          cVar2S14S83P062P066P030nsss(0) <='0';
          end if;
        if(cVar1S15S83P017P044P060P010(0)='1' AND  D( 4)='0' )then
          cVar2S15S83P050nsss(0) <='1';
          else
          cVar2S15S83P050nsss(0) <='0';
          end if;
        if(cVar1S16S83P017P044P060P010(0)='1' AND  A( 2)='1' )then
          cVar2S16S83P015nsss(0) <='1';
          else
          cVar2S16S83P015nsss(0) <='0';
          end if;
        if(cVar1S17S83P017N044P023P052(0)='1' AND  E( 8)='1' )then
          cVar2S17S83P069nsss(0) <='1';
          else
          cVar2S17S83P069nsss(0) <='0';
          end if;
        if(cVar1S18S83P017N044P023P052(0)='1' AND  E( 8)='0' AND A(14)='1' AND A(13)='0' )then
          cVar2S18S83N069P010P012nsss(0) <='1';
          else
          cVar2S18S83N069P010P012nsss(0) <='0';
          end if;
        if(cVar1S19S83P017N044P023N052(0)='1' AND  D( 9)='1' AND A( 7)='1' )then
          cVar2S19S83P063P005nsss(0) <='1';
          else
          cVar2S19S83P063P005nsss(0) <='0';
          end if;
        if(cVar1S20S83P017N044P023N052(0)='1' AND  D( 9)='1' AND A( 7)='0' AND B( 1)='0' )then
          cVar2S20S83P063N005P035nsss(0) <='1';
          else
          cVar2S20S83P063N005P035nsss(0) <='0';
          end if;
        if(cVar1S21S83P017N044P023N052(0)='1' AND  D( 9)='0' AND E( 1)='1' AND A(15)='0' )then
          cVar2S21S83N063P064P008nsss(0) <='1';
          else
          cVar2S21S83N063P064P008nsss(0) <='0';
          end if;
        if(cVar1S23S83P017N044P023N065(0)='1' AND  A( 7)='1' )then
          cVar2S23S83P005nsss(0) <='1';
          else
          cVar2S23S83P005nsss(0) <='0';
          end if;
        if(cVar1S0S84P019P018P057P064(0)='1' AND  B( 1)='0' )then
          cVar2S0S84P035nsss(0) <='1';
          else
          cVar2S0S84P035nsss(0) <='0';
          end if;
        if(cVar1S1S84P019P018P057P064(0)='1' AND  B( 1)='1' AND D( 8)='1' AND E( 0)='0' )then
          cVar2S1S84P035P067P068nsss(0) <='1';
          else
          cVar2S1S84P035P067P068nsss(0) <='0';
          end if;
        if(cVar1S2S84P019P018P057P064(0)='1' AND  A( 9)='1' )then
          cVar2S2S84P001nsss(0) <='1';
          else
          cVar2S2S84P001nsss(0) <='0';
          end if;
        if(cVar1S3S84P019P018P057P064(0)='1' AND  A( 9)='0' AND B( 9)='0' AND D( 1)='1' )then
          cVar2S3S84N001P036P062nsss(0) <='1';
          else
          cVar2S3S84N001P036P062nsss(0) <='0';
          end if;
        if(cVar1S4S84P019P018P057P064(0)='1' AND  A( 9)='0' AND B( 9)='1' AND A( 8)='1' )then
          cVar2S4S84N001P036P003nsss(0) <='1';
          else
          cVar2S4S84N001P036P003nsss(0) <='0';
          end if;
        if(cVar1S5S84P019P018P057P003(0)='1' AND  A(12)='0' )then
          cVar2S5S84P014nsss(0) <='1';
          else
          cVar2S5S84P014nsss(0) <='0';
          end if;
        if(cVar1S6S84P019P018P057N003(0)='1' AND  E( 0)='0' AND B( 9)='0' AND B( 0)='0' )then
          cVar2S6S84P068P036P037nsss(0) <='1';
          else
          cVar2S6S84P068P036P037nsss(0) <='0';
          end if;
        if(cVar1S7S84P019P018P057N003(0)='1' AND  E( 0)='0' AND B( 9)='1' AND B(12)='1' )then
          cVar2S7S84P068P036P030nsss(0) <='1';
          else
          cVar2S7S84P068P036P030nsss(0) <='0';
          end if;
        if(cVar1S8S84P019P018P057N003(0)='1' AND  E( 0)='1' AND B( 0)='1' AND A( 4)='1' )then
          cVar2S8S84P068P037P011nsss(0) <='1';
          else
          cVar2S8S84P068P037P011nsss(0) <='0';
          end if;
        if(cVar1S9S84P019P018P033P014(0)='1' AND  B(12)='1' AND E(11)='1' )then
          cVar2S9S84P030P057nsss(0) <='1';
          else
          cVar2S9S84P030P057nsss(0) <='0';
          end if;
        if(cVar1S10S84P019P018P033P014(0)='1' AND  B(12)='1' AND E(11)='0' AND E( 0)='1' )then
          cVar2S10S84P030N057P068nsss(0) <='1';
          else
          cVar2S10S84P030N057P068nsss(0) <='0';
          end if;
        if(cVar1S11S84P019P018P033P014(0)='1' AND  B(12)='0' AND B( 3)='1' )then
          cVar2S11S84N030P031nsss(0) <='1';
          else
          cVar2S11S84N030P031nsss(0) <='0';
          end if;
        if(cVar1S12S84P019P018P033P014(0)='1' AND  E( 9)='1' AND D( 2)='1' )then
          cVar2S12S84P065P058nsss(0) <='1';
          else
          cVar2S12S84P065P058nsss(0) <='0';
          end if;
        if(cVar1S13S84P019P018P033P014(0)='1' AND  E( 9)='1' AND D( 2)='0' AND A(13)='0' )then
          cVar2S13S84P065N058P012nsss(0) <='1';
          else
          cVar2S13S84P065N058P012nsss(0) <='0';
          end if;
        if(cVar1S14S84P019P018P033P014(0)='1' AND  E( 9)='0' AND B( 9)='1' AND A( 1)='0' )then
          cVar2S14S84N065P036P017nsss(0) <='1';
          else
          cVar2S14S84N065P036P017nsss(0) <='0';
          end if;
        if(cVar1S15S84P019P018P033P014(0)='1' AND  E( 9)='0' AND B( 9)='0' AND B( 6)='1' )then
          cVar2S15S84N065N036P025nsss(0) <='1';
          else
          cVar2S15S84N065N036P025nsss(0) <='0';
          end if;
        if(cVar1S16S84P019P018P033P013(0)='1' AND  D( 8)='0' )then
          cVar2S16S84P067nsss(0) <='1';
          else
          cVar2S16S84P067nsss(0) <='0';
          end if;
        if(cVar1S17S84P019P018P033P013(0)='1' AND  D( 8)='1' AND B( 0)='1' )then
          cVar2S17S84P067P037nsss(0) <='1';
          else
          cVar2S17S84P067P037nsss(0) <='0';
          end if;
        if(cVar1S18S84P019P018P033P013(0)='1' AND  D( 8)='1' AND B( 0)='0' AND E( 2)='1' )then
          cVar2S18S84P067N037P060nsss(0) <='1';
          else
          cVar2S18S84P067N037P060nsss(0) <='0';
          end if;
        if(cVar1S19S84P019P018P033N013(0)='1' AND  D(10)='1' AND A(13)='0' )then
          cVar2S19S84P059P012nsss(0) <='1';
          else
          cVar2S19S84P059P012nsss(0) <='0';
          end if;
        if(cVar1S20S84P019P018P033N013(0)='1' AND  D(10)='0' AND B(10)='1' AND E( 2)='1' )then
          cVar2S20S84N059P034P060nsss(0) <='1';
          else
          cVar2S20S84N059P034P060nsss(0) <='0';
          end if;
        if(cVar1S21S84N019P047P006P064(0)='1' AND  D( 5)='0' AND A(15)='0' )then
          cVar2S21S84P046P008nsss(0) <='1';
          else
          cVar2S21S84P046P008nsss(0) <='0';
          end if;
        if(cVar1S22S84N019P047P006P064(0)='1' AND  D( 5)='1' AND E(13)='1' )then
          cVar2S22S84P046P049nsss(0) <='1';
          else
          cVar2S22S84P046P049nsss(0) <='0';
          end if;
        if(cVar1S23S84N019P047N006P066(0)='1' AND  E(13)='1' AND D( 5)='0' AND D(12)='0' )then
          cVar2S23S84P049P046P051nsss(0) <='1';
          else
          cVar2S23S84P049P046P051nsss(0) <='0';
          end if;
        if(cVar1S24S84N019P047N006P066(0)='1' AND  E(13)='0' AND D( 5)='1' )then
          cVar2S24S84N049P046nsss(0) <='1';
          else
          cVar2S24S84N049P046nsss(0) <='0';
          end if;
        if(cVar1S25S84N019P047N006P066(0)='1' AND  E(13)='0' AND D( 5)='0' AND B(15)='1' )then
          cVar2S25S84N049N046P024nsss(0) <='1';
          else
          cVar2S25S84N049N046P024nsss(0) <='0';
          end if;
        if(cVar1S26S84N019P047N006P066(0)='1' AND  E( 8)='1' AND B( 9)='0' )then
          cVar2S26S84P069P036nsss(0) <='1';
          else
          cVar2S26S84P069P036nsss(0) <='0';
          end if;
        if(cVar1S27S84N019P047N006P066(0)='1' AND  E( 8)='0' AND A(10)='1' AND B(14)='1' )then
          cVar2S27S84N069P018P026nsss(0) <='1';
          else
          cVar2S27S84N069P018P026nsss(0) <='0';
          end if;
        if(cVar1S28S84N019N047P043P044(0)='1' AND  A(13)='0' AND E( 8)='0' )then
          cVar2S28S84P012P069nsss(0) <='1';
          else
          cVar2S28S84P012P069nsss(0) <='0';
          end if;
        if(cVar1S29S84N019N047P043P044(0)='1' AND  A(13)='0' AND E( 8)='1' AND E( 0)='0' )then
          cVar2S29S84P012P069P068nsss(0) <='1';
          else
          cVar2S29S84P012P069P068nsss(0) <='0';
          end if;
        if(cVar1S30S84N019N047P043P044(0)='1' AND  A(13)='1' AND A(10)='1' )then
          cVar2S30S84P012P018nsss(0) <='1';
          else
          cVar2S30S84P012P018nsss(0) <='0';
          end if;
        if(cVar1S31S84N019N047P043P044(0)='1' AND  A( 1)='1' )then
          cVar2S31S84P017nsss(0) <='1';
          else
          cVar2S31S84P017nsss(0) <='0';
          end if;
        if(cVar1S32S84N019N047N043P024(0)='1' AND  A( 7)='0' AND D(12)='1' AND D( 4)='0' )then
          cVar2S32S84P005P051P050nsss(0) <='1';
          else
          cVar2S32S84P005P051P050nsss(0) <='0';
          end if;
        if(cVar1S33S84N019N047N043P024(0)='1' AND  A( 7)='1' AND D(15)='1' )then
          cVar2S33S84P005P039nsss(0) <='1';
          else
          cVar2S33S84P005P039nsss(0) <='0';
          end if;
        if(cVar1S34S84N019N047N043P024(0)='1' AND  A( 7)='1' AND D(15)='0' AND D( 6)='1' )then
          cVar2S34S84P005N039P042nsss(0) <='1';
          else
          cVar2S34S84P005N039P042nsss(0) <='0';
          end if;
        if(cVar1S35S84N019N047N043P024(0)='1' AND  D(10)='1' AND A(14)='0' )then
          cVar2S35S84P059P010nsss(0) <='1';
          else
          cVar2S35S84P059P010nsss(0) <='0';
          end if;
        if(cVar1S36S84N019N047N043P024(0)='1' AND  D(10)='0' AND D( 5)='1' AND A( 3)='0' )then
          cVar2S36S84N059P046P013nsss(0) <='1';
          else
          cVar2S36S84N059P046P013nsss(0) <='0';
          end if;
        if(cVar1S37S84N019N047N043P024(0)='1' AND  D(10)='0' AND D( 5)='0' AND E(15)='1' )then
          cVar2S37S84N059N046P041nsss(0) <='1';
          else
          cVar2S37S84N059N046P041nsss(0) <='0';
          end if;
        if(cVar1S0S85P019P051P067P007(0)='1' AND  B( 8)='0' AND D( 2)='1' )then
          cVar2S0S85P021P058nsss(0) <='1';
          else
          cVar2S0S85P021P058nsss(0) <='0';
          end if;
        if(cVar1S1S85P019P051P067P007(0)='1' AND  B( 8)='0' AND D( 2)='0' AND E( 2)='0' )then
          cVar2S1S85P021N058P060nsss(0) <='1';
          else
          cVar2S1S85P021N058P060nsss(0) <='0';
          end if;
        if(cVar1S2S85P019P051P067P007(0)='1' AND  B( 8)='1' AND A(14)='0' AND A( 1)='1' )then
          cVar2S2S85P021P010P017nsss(0) <='1';
          else
          cVar2S2S85P021P010P017nsss(0) <='0';
          end if;
        if(cVar1S3S85P019P051P067P007(0)='1' AND  E( 9)='1' AND A( 4)='1' )then
          cVar2S3S85P065P011nsss(0) <='1';
          else
          cVar2S3S85P065P011nsss(0) <='0';
          end if;
        if(cVar1S4S85P019P051P067P007(0)='1' AND  E( 9)='1' AND A( 4)='0' AND A(11)='1' )then
          cVar2S4S85P065N011P016nsss(0) <='1';
          else
          cVar2S4S85P065N011P016nsss(0) <='0';
          end if;
        if(cVar1S5S85P019P051P067P007(0)='1' AND  E( 9)='0' AND A(13)='1' AND B( 9)='1' )then
          cVar2S5S85N065P012P036nsss(0) <='1';
          else
          cVar2S5S85N065P012P036nsss(0) <='0';
          end if;
        if(cVar1S6S85P019P051P067P007(0)='1' AND  E( 9)='0' AND A(13)='0' AND A( 5)='1' )then
          cVar2S6S85N065N012P009nsss(0) <='1';
          else
          cVar2S6S85N065N012P009nsss(0) <='0';
          end if;
        if(cVar1S7S85P019P051N067P001(0)='1' AND  A( 1)='1' AND A(17)='0' )then
          cVar2S7S85P017P004nsss(0) <='1';
          else
          cVar2S7S85P017P004nsss(0) <='0';
          end if;
        if(cVar1S8S85P019P051N067P001(0)='1' AND  A( 1)='1' AND A(17)='1' AND E( 9)='1' )then
          cVar2S8S85P017P004P065nsss(0) <='1';
          else
          cVar2S8S85P017P004P065nsss(0) <='0';
          end if;
        if(cVar1S9S85P019P051N067P001(0)='1' AND  A( 1)='0' AND E( 8)='0' AND E( 6)='0' )then
          cVar2S9S85N017P069P044nsss(0) <='1';
          else
          cVar2S9S85N017P069P044nsss(0) <='0';
          end if;
        if(cVar1S10S85P019P051N067P001(0)='1' AND  A( 1)='0' AND E( 8)='1' AND A(11)='1' )then
          cVar2S10S85N017P069P016nsss(0) <='1';
          else
          cVar2S10S85N017P069P016nsss(0) <='0';
          end if;
        if(cVar1S11S85P019P051N067P001(0)='1' AND  A(12)='1' AND A(14)='1' )then
          cVar2S11S85P014P010nsss(0) <='1';
          else
          cVar2S11S85P014P010nsss(0) <='0';
          end if;
        if(cVar1S12S85P019P051N067P001(0)='1' AND  A(12)='1' AND A(14)='0' AND E( 2)='1' )then
          cVar2S12S85P014N010P060nsss(0) <='1';
          else
          cVar2S12S85P014N010P060nsss(0) <='0';
          end if;
        if(cVar1S13S85P019P051N067P001(0)='1' AND  A(12)='0' AND E(10)='1' )then
          cVar2S13S85N014P061nsss(0) <='1';
          else
          cVar2S13S85N014P061nsss(0) <='0';
          end if;
        if(cVar1S15S85P019P051P008N027(0)='1' AND  A( 6)='0' AND D( 4)='0' )then
          cVar2S15S85P007P050nsss(0) <='1';
          else
          cVar2S15S85P007P050nsss(0) <='0';
          end if;
        if(cVar1S16S85P019P051P008N027(0)='1' AND  A( 6)='0' AND D( 4)='1' AND B(14)='0' )then
          cVar2S16S85P007P050P026nsss(0) <='1';
          else
          cVar2S16S85P007P050P026nsss(0) <='0';
          end if;
        if(cVar1S17S85P019P051N008P057(0)='1' AND  B(14)='1' AND E( 8)='0' )then
          cVar2S17S85P026P069nsss(0) <='1';
          else
          cVar2S17S85P026P069nsss(0) <='0';
          end if;
        if(cVar1S18S85P019P051N008P057(0)='1' AND  B(14)='0' AND A(16)='1' )then
          cVar2S18S85N026P006nsss(0) <='1';
          else
          cVar2S18S85N026P006nsss(0) <='0';
          end if;
        if(cVar1S19S85P019P051N008P057(0)='1' AND  B(14)='0' AND A(16)='0' AND B(12)='1' )then
          cVar2S19S85N026N006P030nsss(0) <='1';
          else
          cVar2S19S85N026N006P030nsss(0) <='0';
          end if;
        if(cVar1S20S85P019P051N008P057(0)='1' AND  B(12)='1' )then
          cVar2S20S85P030nsss(0) <='1';
          else
          cVar2S20S85P030nsss(0) <='0';
          end if;
        if(cVar1S21S85P019P018P014P033(0)='1' AND  B(10)='0' AND B( 9)='0' AND E(12)='0' )then
          cVar2S21S85P034P036P053nsss(0) <='1';
          else
          cVar2S21S85P034P036P053nsss(0) <='0';
          end if;
        if(cVar1S22S85P019P018P014P033(0)='1' AND  B(10)='0' AND B( 9)='1' AND D(13)='0' )then
          cVar2S22S85P034P036P047nsss(0) <='1';
          else
          cVar2S22S85P034P036P047nsss(0) <='0';
          end if;
        if(cVar1S23S85P019P018P014P033(0)='1' AND  B(10)='1' AND A( 2)='0' AND E( 0)='1' )then
          cVar2S23S85P034P015P068nsss(0) <='1';
          else
          cVar2S23S85P034P015P068nsss(0) <='0';
          end if;
        if(cVar1S24S85P019P018P014P033(0)='1' AND  A( 3)='1' AND D( 9)='1' )then
          cVar2S24S85P013P063nsss(0) <='1';
          else
          cVar2S24S85P013P063nsss(0) <='0';
          end if;
        if(cVar1S25S85P019P018P014P033(0)='1' AND  A( 3)='1' AND D( 9)='0' AND A( 4)='1' )then
          cVar2S25S85P013N063P011nsss(0) <='1';
          else
          cVar2S25S85P013N063P011nsss(0) <='0';
          end if;
        if(cVar1S26S85P019P018P014P033(0)='1' AND  A( 3)='0' AND D(10)='1' )then
          cVar2S26S85N013P059nsss(0) <='1';
          else
          cVar2S26S85N013P059nsss(0) <='0';
          end if;
        if(cVar1S27S85P019P018P014P023(0)='1' AND  A( 3)='0' )then
          cVar2S27S85P013nsss(0) <='1';
          else
          cVar2S27S85P013nsss(0) <='0';
          end if;
        if(cVar1S28S85P019P018P014N023(0)='1' AND  B(10)='1' AND E( 8)='1' )then
          cVar2S28S85P034P069nsss(0) <='1';
          else
          cVar2S28S85P034P069nsss(0) <='0';
          end if;
        if(cVar1S29S85P019P018P014N023(0)='1' AND  B(10)='1' AND E( 8)='0' AND A( 1)='1' )then
          cVar2S29S85P034N069P017nsss(0) <='1';
          else
          cVar2S29S85P034N069P017nsss(0) <='0';
          end if;
        if(cVar1S30S85P019P018P014N023(0)='1' AND  B(10)='0' AND E( 0)='1' AND E( 9)='1' )then
          cVar2S30S85N034P068P065nsss(0) <='1';
          else
          cVar2S30S85N034P068P065nsss(0) <='0';
          end if;
        if(cVar1S31S85P019P018P014N023(0)='1' AND  B(10)='0' AND E( 0)='0' AND B( 1)='1' )then
          cVar2S31S85N034N068P035nsss(0) <='1';
          else
          cVar2S31S85N034N068P035nsss(0) <='0';
          end if;
        if(cVar1S32S85P019N018P033P012(0)='1' AND  A(12)='0' AND E( 9)='0' )then
          cVar2S32S85P014P065nsss(0) <='1';
          else
          cVar2S32S85P014P065nsss(0) <='0';
          end if;
        if(cVar1S33S85P019N018P033P012(0)='1' AND  A(12)='1' AND E( 0)='0' AND B( 0)='0' )then
          cVar2S33S85P014P068P037nsss(0) <='1';
          else
          cVar2S33S85P014P068P037nsss(0) <='0';
          end if;
        if(cVar1S34S85P019N018P033N012(0)='1' AND  A(18)='0' AND D(13)='1' )then
          cVar2S34S85P002P047nsss(0) <='1';
          else
          cVar2S34S85P002P047nsss(0) <='0';
          end if;
        if(cVar1S35S85P019N018P033N012(0)='1' AND  A(18)='0' AND D(13)='0' AND D( 9)='1' )then
          cVar2S35S85P002N047P063nsss(0) <='1';
          else
          cVar2S35S85P002N047P063nsss(0) <='0';
          end if;
        if(cVar1S36S85P019N018N033P010(0)='1' AND  D( 4)='1' )then
          cVar2S36S85P050nsss(0) <='1';
          else
          cVar2S36S85P050nsss(0) <='0';
          end if;
        if(cVar1S37S85P019N018N033P010(0)='1' AND  D( 4)='0' AND A( 1)='1' AND A( 5)='0' )then
          cVar2S37S85N050P017P009nsss(0) <='1';
          else
          cVar2S37S85N050P017P009nsss(0) <='0';
          end if;
        if(cVar1S38S85P019N018N033P010(0)='1' AND  D( 4)='0' AND A( 1)='0' AND D(13)='1' )then
          cVar2S38S85N050N017P047nsss(0) <='1';
          else
          cVar2S38S85N050N017P047nsss(0) <='0';
          end if;
        if(cVar1S39S85P019N018N033N010(0)='1' AND  E( 4)='0' AND D( 2)='1' AND B( 0)='1' )then
          cVar2S39S85P052P058P037nsss(0) <='1';
          else
          cVar2S39S85P052P058P037nsss(0) <='0';
          end if;
        if(cVar1S40S85P019N018N033N010(0)='1' AND  E( 4)='1' AND A( 3)='1' AND A( 2)='0' )then
          cVar2S40S85P052P013P015nsss(0) <='1';
          else
          cVar2S40S85P052P013P015nsss(0) <='0';
          end if;
        if(cVar1S41S85P019N018N033N010(0)='1' AND  E( 4)='1' AND A( 3)='0' AND B(14)='1' )then
          cVar2S41S85P052N013P026nsss(0) <='1';
          else
          cVar2S41S85P052N013P026nsss(0) <='0';
          end if;
        if(cVar1S0S86P019P018P036P014(0)='1' AND  E( 3)='1' )then
          cVar2S0S86P056nsss(0) <='1';
          else
          cVar2S0S86P056nsss(0) <='0';
          end if;
        if(cVar1S1S86P019P018P036P014(0)='1' AND  E( 3)='0' AND A( 8)='1' )then
          cVar2S1S86N056P003nsss(0) <='1';
          else
          cVar2S1S86N056P003nsss(0) <='0';
          end if;
        if(cVar1S2S86P019P018P036P014(0)='1' AND  E( 3)='0' AND A( 8)='0' AND A(15)='0' )then
          cVar2S2S86N056N003P008nsss(0) <='1';
          else
          cVar2S2S86N056N003P008nsss(0) <='0';
          end if;
        if(cVar1S3S86P019P018P036N014(0)='1' AND  E( 0)='1' AND A( 3)='0' AND D(10)='0' )then
          cVar2S3S86P068P013P059nsss(0) <='1';
          else
          cVar2S3S86P068P013P059nsss(0) <='0';
          end if;
        if(cVar1S4S86P019P018P036N014(0)='1' AND  E( 0)='1' AND A( 3)='1' AND A( 2)='1' )then
          cVar2S4S86P068P013P015nsss(0) <='1';
          else
          cVar2S4S86P068P013P015nsss(0) <='0';
          end if;
        if(cVar1S5S86P019P018P036N014(0)='1' AND  E( 0)='0' AND D( 0)='0' AND A( 2)='1' )then
          cVar2S5S86N068P066P015nsss(0) <='1';
          else
          cVar2S5S86N068P066P015nsss(0) <='0';
          end if;
        if(cVar1S6S86P019P018N036P069(0)='1' AND  A(16)='0' AND A( 7)='1' )then
          cVar2S6S86P006P005nsss(0) <='1';
          else
          cVar2S6S86P006P005nsss(0) <='0';
          end if;
        if(cVar1S7S86P019P018N036P069(0)='1' AND  A(16)='0' AND A( 7)='0' AND A(11)='0' )then
          cVar2S7S86P006N005P016nsss(0) <='1';
          else
          cVar2S7S86P006N005P016nsss(0) <='0';
          end if;
        if(cVar1S8S86P019P018N036P069(0)='1' AND  A(16)='1' AND A( 9)='1' )then
          cVar2S8S86P006P001nsss(0) <='1';
          else
          cVar2S8S86P006P001nsss(0) <='0';
          end if;
        if(cVar1S9S86P019P018N036P069(0)='1' AND  A(16)='1' AND A( 9)='0' AND B( 8)='1' )then
          cVar2S9S86P006N001P021nsss(0) <='1';
          else
          cVar2S9S86P006N001P021nsss(0) <='0';
          end if;
        if(cVar1S10S86P019P018N036P069(0)='1' AND  B(17)='1' )then
          cVar2S10S86P020nsss(0) <='1';
          else
          cVar2S10S86P020nsss(0) <='0';
          end if;
        if(cVar1S11S86P019P018N036P069(0)='1' AND  B(17)='0' AND A(18)='1' )then
          cVar2S11S86N020P002nsss(0) <='1';
          else
          cVar2S11S86N020P002nsss(0) <='0';
          end if;
        if(cVar1S12S86P019P018P055P030(0)='1' AND  B( 0)='0' )then
          cVar2S12S86P037nsss(0) <='1';
          else
          cVar2S12S86P037nsss(0) <='0';
          end if;
        if(cVar1S13S86P019P018P055P030(0)='1' AND  B( 0)='1' AND A( 3)='1' )then
          cVar2S13S86P037P013nsss(0) <='1';
          else
          cVar2S13S86P037P013nsss(0) <='0';
          end if;
        if(cVar1S14S86P019P018P055N030(0)='1' AND  A( 4)='1' AND D( 0)='0' )then
          cVar2S14S86P011P066nsss(0) <='1';
          else
          cVar2S14S86P011P066nsss(0) <='0';
          end if;
        if(cVar1S15S86P019P018P055N030(0)='1' AND  A( 4)='0' AND E(10)='1' )then
          cVar2S15S86N011P061nsss(0) <='1';
          else
          cVar2S15S86N011P061nsss(0) <='0';
          end if;
        if(cVar1S16S86P019P018P055N030(0)='1' AND  A( 4)='0' AND E(10)='0' AND E( 8)='1' )then
          cVar2S16S86N011N061P069nsss(0) <='1';
          else
          cVar2S16S86N011N061P069nsss(0) <='0';
          end if;
        if(cVar1S17S86P019P018N055P046(0)='1' AND  B( 2)='0' AND E(11)='0' AND D( 1)='1' )then
          cVar2S17S86P033P057P062nsss(0) <='1';
          else
          cVar2S17S86P033P057P062nsss(0) <='0';
          end if;
        if(cVar1S18S86P019P018N055P046(0)='1' AND  B( 2)='0' AND E(11)='1' AND D(10)='1' )then
          cVar2S18S86P033P057P059nsss(0) <='1';
          else
          cVar2S18S86P033P057P059nsss(0) <='0';
          end if;
        if(cVar1S19S86P019P018N055P046(0)='1' AND  B( 2)='1' AND A( 3)='1' AND D( 8)='0' )then
          cVar2S19S86P033P013P067nsss(0) <='1';
          else
          cVar2S19S86P033P013P067nsss(0) <='0';
          end if;
        if(cVar1S20S86P019P018N055P046(0)='1' AND  B( 6)='1' )then
          cVar2S20S86P025nsss(0) <='1';
          else
          cVar2S20S86P025nsss(0) <='0';
          end if;
        if(cVar1S21S86N019P067P002P031(0)='1' AND  B(17)='0' AND A( 7)='0' AND A( 1)='0' )then
          cVar2S21S86P020P005P017nsss(0) <='1';
          else
          cVar2S21S86P020P005P017nsss(0) <='0';
          end if;
        if(cVar1S22S86N019P067P002P031(0)='1' AND  B(17)='0' AND A( 7)='1' AND D( 1)='1' )then
          cVar2S22S86P020P005P062nsss(0) <='1';
          else
          cVar2S22S86P020P005P062nsss(0) <='0';
          end if;
        if(cVar1S23S86N019P067P002P031(0)='1' AND  B(17)='1' AND D( 0)='1' )then
          cVar2S23S86P020P066nsss(0) <='1';
          else
          cVar2S23S86P020P066nsss(0) <='0';
          end if;
        if(cVar1S24S86N019P067P002P031(0)='1' AND  D(10)='1' AND A( 3)='1' )then
          cVar2S24S86P059P013nsss(0) <='1';
          else
          cVar2S24S86P059P013nsss(0) <='0';
          end if;
        if(cVar1S25S86N019P067P002P031(0)='1' AND  D(10)='0' AND A(13)='1' AND E( 3)='0' )then
          cVar2S25S86N059P012P056nsss(0) <='1';
          else
          cVar2S25S86N059P012P056nsss(0) <='0';
          end if;
        if(cVar1S27S86N019P067P002N064(0)='1' AND  D( 9)='0' AND A( 1)='1' AND A(10)='1' )then
          cVar2S27S86P063P017P018nsss(0) <='1';
          else
          cVar2S27S86P063P017P018nsss(0) <='0';
          end if;
        if(cVar1S28S86N019N067P017P011(0)='1' AND  D(15)='0' AND D(10)='1' )then
          cVar2S28S86P039P059nsss(0) <='1';
          else
          cVar2S28S86P039P059nsss(0) <='0';
          end if;
        if(cVar1S29S86N019N067P017P011(0)='1' AND  D(15)='0' AND D(10)='0' AND B(11)='0' )then
          cVar2S29S86P039N059P032nsss(0) <='1';
          else
          cVar2S29S86P039N059P032nsss(0) <='0';
          end if;
        if(cVar1S30S86N019N067P017N011(0)='1' AND  B( 4)='0' AND D( 4)='1' )then
          cVar2S30S86P029P050nsss(0) <='1';
          else
          cVar2S30S86P029P050nsss(0) <='0';
          end if;
        if(cVar1S31S86N019N067P017N011(0)='1' AND  B( 4)='0' AND D( 4)='0' AND A(18)='1' )then
          cVar2S31S86P029N050P002nsss(0) <='1';
          else
          cVar2S31S86P029N050P002nsss(0) <='0';
          end if;
        if(cVar1S32S86N019N067P017N011(0)='1' AND  B( 4)='1' AND B(14)='0' AND B( 1)='1' )then
          cVar2S32S86P029P026P035nsss(0) <='1';
          else
          cVar2S32S86P029P026P035nsss(0) <='0';
          end if;
        if(cVar1S33S86N019N067N017P069(0)='1' AND  B( 5)='1' AND D( 4)='1' )then
          cVar2S33S86P027P050nsss(0) <='1';
          else
          cVar2S33S86P027P050nsss(0) <='0';
          end if;
        if(cVar1S34S86N019N067N017P069(0)='1' AND  B( 5)='1' AND D( 4)='0' AND A(15)='1' )then
          cVar2S34S86P027N050P008nsss(0) <='1';
          else
          cVar2S34S86P027N050P008nsss(0) <='0';
          end if;
        if(cVar1S35S86N019N067N017P069(0)='1' AND  B( 5)='0' AND E( 5)='0' AND A(14)='1' )then
          cVar2S35S86N027P048P010nsss(0) <='1';
          else
          cVar2S35S86N027P048P010nsss(0) <='0';
          end if;
        if(cVar1S36S86N019N067N017P069(0)='1' AND  B( 5)='0' AND E( 5)='1' AND B( 6)='1' )then
          cVar2S36S86N027P048P025nsss(0) <='1';
          else
          cVar2S36S86N027P048P025nsss(0) <='0';
          end if;
        if(cVar1S37S86N019N067N017P069(0)='1' AND  E( 9)='1' AND B( 9)='1' )then
          cVar2S37S86P065P036nsss(0) <='1';
          else
          cVar2S37S86P065P036nsss(0) <='0';
          end if;
        if(cVar1S38S86N019N067N017P069(0)='1' AND  E( 9)='1' AND B( 9)='0' AND A(11)='1' )then
          cVar2S38S86P065N036P016nsss(0) <='1';
          else
          cVar2S38S86P065N036P016nsss(0) <='0';
          end if;
        if(cVar1S39S86N019N067N017P069(0)='1' AND  E( 9)='0' AND D(13)='1' )then
          cVar2S39S86N065P047nsss(0) <='1';
          else
          cVar2S39S86N065P047nsss(0) <='0';
          end if;
        if(cVar1S40S86N019N067N017P069(0)='1' AND  E( 9)='0' AND D(13)='0' AND E(11)='1' )then
          cVar2S40S86N065N047P057nsss(0) <='1';
          else
          cVar2S40S86N065N047P057nsss(0) <='0';
          end if;
        if(cVar1S0S87P017P002P038P066(0)='1' AND  A( 5)='1' AND A(15)='0' )then
          cVar2S0S87P009P008nsss(0) <='1';
          else
          cVar2S0S87P009P008nsss(0) <='0';
          end if;
        if(cVar1S1S87P017P002P038P066(0)='1' AND  A( 5)='1' AND A(15)='1' AND A(11)='0' )then
          cVar2S1S87P009P008P016nsss(0) <='1';
          else
          cVar2S1S87P009P008P016nsss(0) <='0';
          end if;
        if(cVar1S2S87P017P002P038P066(0)='1' AND  A( 5)='0' AND E( 8)='1' )then
          cVar2S2S87N009P069nsss(0) <='1';
          else
          cVar2S2S87N009P069nsss(0) <='0';
          end if;
        if(cVar1S3S87P017P002P038P066(0)='1' AND  A( 5)='0' AND E( 8)='0' AND A(10)='1' )then
          cVar2S3S87N009N069P018nsss(0) <='1';
          else
          cVar2S3S87N009N069P018nsss(0) <='0';
          end if;
        if(cVar1S4S87P017P002P038N066(0)='1' AND  A( 5)='0' AND E( 0)='0' AND A(10)='0' )then
          cVar2S4S87P009P068P018nsss(0) <='1';
          else
          cVar2S4S87P009P068P018nsss(0) <='0';
          end if;
        if(cVar1S5S87P017P002P038N066(0)='1' AND  A( 5)='1' AND D( 4)='1' AND A(13)='0' )then
          cVar2S5S87P009P050P012nsss(0) <='1';
          else
          cVar2S5S87P009P050P012nsss(0) <='0';
          end if;
        if(cVar1S6S87P017P002P038N066(0)='1' AND  A( 5)='1' AND D( 4)='0' AND D(13)='1' )then
          cVar2S6S87P009N050P047nsss(0) <='1';
          else
          cVar2S6S87P009N050P047nsss(0) <='0';
          end if;
        if(cVar1S8S87P017P002P038N004(0)='1' AND  E( 1)='0' AND A( 5)='1' )then
          cVar2S8S87N064P009nsss(0) <='1';
          else
          cVar2S8S87N064P009nsss(0) <='0';
          end if;
        if(cVar1S10S87P017P002N040P013(0)='1' AND  B( 9)='1' )then
          cVar2S10S87P036nsss(0) <='1';
          else
          cVar2S10S87P036nsss(0) <='0';
          end if;
        if(cVar1S11S87P017P002N040P013(0)='1' AND  B( 9)='0' AND A( 0)='1' AND A(12)='0' )then
          cVar2S11S87N036P019P014nsss(0) <='1';
          else
          cVar2S11S87N036P019P014nsss(0) <='0';
          end if;
        if(cVar1S12S87P017P002N040N013(0)='1' AND  B( 1)='1' AND D( 8)='1' )then
          cVar2S12S87P035P067nsss(0) <='1';
          else
          cVar2S12S87P035P067nsss(0) <='0';
          end if;
        if(cVar1S13S87P017P002N040N013(0)='1' AND  B( 1)='1' AND D( 8)='0' AND A(10)='0' )then
          cVar2S13S87P035N067P018nsss(0) <='1';
          else
          cVar2S13S87P035N067P018nsss(0) <='0';
          end if;
        if(cVar1S14S87P017P002N040N013(0)='1' AND  B( 1)='0' AND B( 0)='1' AND A( 0)='0' )then
          cVar2S14S87N035P037P019nsss(0) <='1';
          else
          cVar2S14S87N035P037P019nsss(0) <='0';
          end if;
        if(cVar1S15S87N017P019P052P003(0)='1' AND  E(11)='1' )then
          cVar2S15S87P057nsss(0) <='1';
          else
          cVar2S15S87P057nsss(0) <='0';
          end if;
        if(cVar1S16S87N017P019P052P003(0)='1' AND  E(11)='0' AND B( 0)='1' AND E(12)='0' )then
          cVar2S16S87N057P037P053nsss(0) <='1';
          else
          cVar2S16S87N057P037P053nsss(0) <='0';
          end if;
        if(cVar1S17S87N017P019P052P003(0)='1' AND  E(11)='0' AND B( 0)='0' AND D(12)='1' )then
          cVar2S17S87N057N037P051nsss(0) <='1';
          else
          cVar2S17S87N057N037P051nsss(0) <='0';
          end if;
        if(cVar1S18S87N017P019P052N003(0)='1' AND  D( 6)='1' AND D( 9)='0' )then
          cVar2S18S87P042P063nsss(0) <='1';
          else
          cVar2S18S87P042P063nsss(0) <='0';
          end if;
        if(cVar1S19S87N017P019P052N003(0)='1' AND  D( 6)='0' AND E( 3)='1' AND E(12)='0' )then
          cVar2S19S87N042P056P053nsss(0) <='1';
          else
          cVar2S19S87N042P056P053nsss(0) <='0';
          end if;
        if(cVar1S20S87N017P019P052N003(0)='1' AND  D( 6)='0' AND E( 3)='0' AND A(14)='0' )then
          cVar2S20S87N042N056P010nsss(0) <='1';
          else
          cVar2S20S87N042N056P010nsss(0) <='0';
          end if;
        if(cVar1S21S87N017P019P052P009(0)='1' AND  B( 4)='1' )then
          cVar2S21S87P029nsss(0) <='1';
          else
          cVar2S21S87P029nsss(0) <='0';
          end if;
        if(cVar1S22S87N017P019P052P009(0)='1' AND  B( 4)='0' AND A(10)='0' )then
          cVar2S22S87N029P018nsss(0) <='1';
          else
          cVar2S22S87N029P018nsss(0) <='0';
          end if;
        if(cVar1S23S87N017P019P052N009(0)='1' AND  A(14)='1' AND D( 4)='1' )then
          cVar2S23S87P010P050nsss(0) <='1';
          else
          cVar2S23S87P010P050nsss(0) <='0';
          end if;
        if(cVar1S24S87N017P019P052N009(0)='1' AND  A(14)='0' AND B(14)='1' AND A(15)='1' )then
          cVar2S24S87N010P026P008nsss(0) <='1';
          else
          cVar2S24S87N010P026P008nsss(0) <='0';
          end if;
        if(cVar1S25S87N017P019P052N009(0)='1' AND  A(14)='0' AND B(14)='0' AND A( 3)='1' )then
          cVar2S25S87N010N026P013nsss(0) <='1';
          else
          cVar2S25S87N010N026P013nsss(0) <='0';
          end if;
        if(cVar1S26S87N017N019P069P067(0)='1' AND  A(10)='1' AND E( 3)='1' )then
          cVar2S26S87P018P056nsss(0) <='1';
          else
          cVar2S26S87P018P056nsss(0) <='0';
          end if;
        if(cVar1S27S87N017N019P069P067(0)='1' AND  A(10)='1' AND E( 3)='0' AND A(14)='0' )then
          cVar2S27S87P018N056P010nsss(0) <='1';
          else
          cVar2S27S87P018N056P010nsss(0) <='0';
          end if;
        if(cVar1S28S87N017N019P069P067(0)='1' AND  A(10)='0' AND B( 8)='1' )then
          cVar2S28S87N018P021nsss(0) <='1';
          else
          cVar2S28S87N018P021nsss(0) <='0';
          end if;
        if(cVar1S29S87N017N019P069P067(0)='1' AND  A(10)='0' AND B( 8)='0' AND A(12)='1' )then
          cVar2S29S87N018N021P014nsss(0) <='1';
          else
          cVar2S29S87N018N021P014nsss(0) <='0';
          end if;
        if(cVar1S30S87N017N019P069P067(0)='1' AND  B(11)='1' AND D(10)='1' )then
          cVar2S30S87P032P059nsss(0) <='1';
          else
          cVar2S30S87P032P059nsss(0) <='0';
          end if;
        if(cVar1S31S87N017N019P069P067(0)='1' AND  B(11)='0' AND D(13)='1' )then
          cVar2S31S87N032P047nsss(0) <='1';
          else
          cVar2S31S87N032P047nsss(0) <='0';
          end if;
        if(cVar1S32S87N017N019P069P067(0)='1' AND  B(11)='0' AND D(13)='0' AND E(14)='1' )then
          cVar2S32S87N032N047P045nsss(0) <='1';
          else
          cVar2S32S87N032N047P045nsss(0) <='0';
          end if;
        if(cVar1S33S87N017N019P069P064(0)='1' AND  A(10)='0' AND B( 0)='0' AND A(11)='1' )then
          cVar2S33S87P018P037P016nsss(0) <='1';
          else
          cVar2S33S87P018P037P016nsss(0) <='0';
          end if;
        if(cVar1S34S87N017N019P069P064(0)='1' AND  A(10)='0' AND B( 0)='1' AND A( 2)='1' )then
          cVar2S34S87P018P037P015nsss(0) <='1';
          else
          cVar2S34S87P018P037P015nsss(0) <='0';
          end if;
        if(cVar1S35S87N017N019P069P064(0)='1' AND  A(10)='1' AND B( 9)='1' AND A( 2)='0' )then
          cVar2S35S87P018P036P015nsss(0) <='1';
          else
          cVar2S35S87P018P036P015nsss(0) <='0';
          end if;
        if(cVar1S36S87N017N019P069P064(0)='1' AND  A(10)='1' AND B( 9)='0' AND A(12)='1' )then
          cVar2S36S87P018N036P014nsss(0) <='1';
          else
          cVar2S36S87P018N036P014nsss(0) <='0';
          end if;
        if(cVar1S37S87N017N019P069N064(0)='1' AND  D( 1)='0' AND B( 0)='1' AND B(15)='0' )then
          cVar2S37S87P062P037P024nsss(0) <='1';
          else
          cVar2S37S87P062P037P024nsss(0) <='0';
          end if;
        if(cVar1S38S87N017N019P069N064(0)='1' AND  D( 1)='0' AND B( 0)='0' AND D( 2)='1' )then
          cVar2S38S87P062N037P058nsss(0) <='1';
          else
          cVar2S38S87P062N037P058nsss(0) <='0';
          end if;
        if(cVar1S39S87N017N019P069N064(0)='1' AND  D( 1)='1' AND A( 4)='1' )then
          cVar2S39S87P062P011nsss(0) <='1';
          else
          cVar2S39S87P062P011nsss(0) <='0';
          end if;
        if(cVar1S0S88P014P016P018P012(0)='1' AND  A( 0)='0' AND A( 1)='0' )then
          cVar2S0S88P019P017nsss(0) <='1';
          else
          cVar2S0S88P019P017nsss(0) <='0';
          end if;
        if(cVar1S1S88P014P016P018P012(0)='1' AND  A( 0)='1' AND A( 2)='1' )then
          cVar2S1S88P019P015nsss(0) <='1';
          else
          cVar2S1S88P019P015nsss(0) <='0';
          end if;
        if(cVar1S2S88P014P016P018P012(0)='1' AND  A( 0)='1' AND A( 2)='0' AND D( 5)='1' )then
          cVar2S2S88P019N015P046nsss(0) <='1';
          else
          cVar2S2S88P019N015P046nsss(0) <='0';
          end if;
        if(cVar1S3S88P014P016P018P012(0)='1' AND  D( 2)='1' AND D( 9)='1' )then
          cVar2S3S88P058P063nsss(0) <='1';
          else
          cVar2S3S88P058P063nsss(0) <='0';
          end if;
        if(cVar1S4S88P014P016P018P012(0)='1' AND  D( 2)='1' AND D( 9)='0' AND E( 1)='0' )then
          cVar2S4S88P058N063P064nsss(0) <='1';
          else
          cVar2S4S88P058N063P064nsss(0) <='0';
          end if;
        if(cVar1S5S88P014P016P018P012(0)='1' AND  D( 2)='0' AND D( 3)='1' AND A( 0)='0' )then
          cVar2S5S88N058P054P019nsss(0) <='1';
          else
          cVar2S5S88N058P054P019nsss(0) <='0';
          end if;
        if(cVar1S6S88P014P016P018P033(0)='1' AND  A( 8)='0' AND A( 2)='0' )then
          cVar2S6S88P003P015nsss(0) <='1';
          else
          cVar2S6S88P003P015nsss(0) <='0';
          end if;
        if(cVar1S7S88P014P016P018P033(0)='1' AND  A( 8)='0' AND A( 2)='1' AND D(10)='1' )then
          cVar2S7S88P003P015P059nsss(0) <='1';
          else
          cVar2S7S88P003P015P059nsss(0) <='0';
          end if;
        if(cVar1S8S88P014P016P018P033(0)='1' AND  A( 8)='1' AND D( 2)='0' AND A( 0)='1' )then
          cVar2S8S88P003P058P019nsss(0) <='1';
          else
          cVar2S8S88P003P058P019nsss(0) <='0';
          end if;
        if(cVar1S9S88P014P016P018N033(0)='1' AND  B( 1)='1' AND E( 8)='0' )then
          cVar2S9S88P035P069nsss(0) <='1';
          else
          cVar2S9S88P035P069nsss(0) <='0';
          end if;
        if(cVar1S10S88P014P016P018N033(0)='1' AND  B( 1)='1' AND E( 8)='1' AND B( 0)='0' )then
          cVar2S10S88P035P069P037nsss(0) <='1';
          else
          cVar2S10S88P035P069P037nsss(0) <='0';
          end if;
        if(cVar1S11S88P014P016P018N033(0)='1' AND  B( 1)='0' AND A( 0)='1' AND E( 2)='0' )then
          cVar2S11S88N035P019P060nsss(0) <='1';
          else
          cVar2S11S88N035P019P060nsss(0) <='0';
          end if;
        if(cVar1S12S88P014P016P018N033(0)='1' AND  B( 1)='0' AND A( 0)='0' AND D( 2)='1' )then
          cVar2S12S88N035N019P058nsss(0) <='1';
          else
          cVar2S12S88N035N019P058nsss(0) <='0';
          end if;
        if(cVar1S13S88P014N016P021P040(0)='1' AND  A(18)='1' )then
          cVar2S13S88P002nsss(0) <='1';
          else
          cVar2S13S88P002nsss(0) <='0';
          end if;
        if(cVar1S14S88P014N016P021P040(0)='1' AND  A(18)='0' AND D( 6)='1' )then
          cVar2S14S88N002P042nsss(0) <='1';
          else
          cVar2S14S88N002P042nsss(0) <='0';
          end if;
        if(cVar1S15S88P014N016P021P040(0)='1' AND  A(18)='0' AND D( 6)='0' AND A( 1)='0' )then
          cVar2S15S88N002N042P017nsss(0) <='1';
          else
          cVar2S15S88N002N042P017nsss(0) <='0';
          end if;
        if(cVar1S16S88P014N016P021N040(0)='1' AND  E( 6)='1' )then
          cVar2S16S88P044nsss(0) <='1';
          else
          cVar2S16S88P044nsss(0) <='0';
          end if;
        if(cVar1S17S88P014N016P021N040(0)='1' AND  E( 6)='0' AND A(17)='0' AND E( 1)='1' )then
          cVar2S17S88N044P004P064nsss(0) <='1';
          else
          cVar2S17S88N044P004P064nsss(0) <='0';
          end if;
        if(cVar1S18S88P014N016N021P054(0)='1' AND  E( 5)='0' AND B( 2)='1' )then
          cVar2S18S88P048P033nsss(0) <='1';
          else
          cVar2S18S88P048P033nsss(0) <='0';
          end if;
        if(cVar1S19S88P014N016N021P054(0)='1' AND  E( 5)='0' AND B( 2)='0' AND A(10)='0' )then
          cVar2S19S88P048N033P018nsss(0) <='1';
          else
          cVar2S19S88P048N033P018nsss(0) <='0';
          end if;
        if(cVar1S20S88P014N016N021P054(0)='1' AND  E( 5)='1' AND B( 3)='0' AND A( 5)='1' )then
          cVar2S20S88P048N031P009nsss(0) <='1';
          else
          cVar2S20S88P048N031P009nsss(0) <='0';
          end if;
        if(cVar1S21S88P014N016N021N054(0)='1' AND  A( 1)='1' AND A( 5)='1' )then
          cVar2S21S88P017P009nsss(0) <='1';
          else
          cVar2S21S88P017P009nsss(0) <='0';
          end if;
        if(cVar1S22S88P014P021P003P019(0)='1' AND  B( 5)='0' )then
          cVar2S22S88P027nsss(0) <='1';
          else
          cVar2S22S88P027nsss(0) <='0';
          end if;
        if(cVar1S23S88P014P021P003N019(0)='1' AND  A( 4)='0' AND B(13)='0' AND A(19)='0' )then
          cVar2S23S88P011P028P000nsss(0) <='1';
          else
          cVar2S23S88P011P028P000nsss(0) <='0';
          end if;
        if(cVar1S24S88P014P021N003P023(0)='1' AND  D( 6)='1' )then
          cVar2S24S88P042nsss(0) <='1';
          else
          cVar2S24S88P042nsss(0) <='0';
          end if;
        if(cVar1S25S88P014P021N003P023(0)='1' AND  D( 6)='0' AND A( 2)='1' AND A( 5)='1' )then
          cVar2S25S88N042P015P009nsss(0) <='1';
          else
          cVar2S25S88N042P015P009nsss(0) <='0';
          end if;
        if(cVar1S26S88P014P021N003P023(0)='1' AND  D( 6)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar2S26S88N042N015P017nsss(0) <='1';
          else
          cVar2S26S88N042N015P017nsss(0) <='0';
          end if;
        if(cVar1S27S88P014P021N003N023(0)='1' AND  A(13)='0' AND A( 1)='1' AND E( 1)='0' )then
          cVar2S27S88P012P017P064nsss(0) <='1';
          else
          cVar2S27S88P012P017P064nsss(0) <='0';
          end if;
        if(cVar1S28S88P014P021N003N023(0)='1' AND  A(13)='0' AND A( 1)='0' AND A(17)='1' )then
          cVar2S28S88P012N017P004nsss(0) <='1';
          else
          cVar2S28S88P012N017P004nsss(0) <='0';
          end if;
        if(cVar1S29S88P014P021N003N023(0)='1' AND  A(13)='1' AND E(15)='0' AND D(10)='1' )then
          cVar2S29S88P012P041P059nsss(0) <='1';
          else
          cVar2S29S88P012P041P059nsss(0) <='0';
          end if;
        if(cVar1S30S88P014P021P026P037(0)='1' AND  B( 9)='1' )then
          cVar2S30S88P036nsss(0) <='1';
          else
          cVar2S30S88P036nsss(0) <='0';
          end if;
        if(cVar1S31S88P014P021P026P037(0)='1' AND  B( 9)='0' AND A(10)='0' AND A( 4)='1' )then
          cVar2S31S88N036P018P011nsss(0) <='1';
          else
          cVar2S31S88N036P018P011nsss(0) <='0';
          end if;
        if(cVar1S32S88P014P021P026N037(0)='1' AND  B(11)='1' AND E(10)='1' )then
          cVar2S32S88P032P061nsss(0) <='1';
          else
          cVar2S32S88P032P061nsss(0) <='0';
          end if;
        if(cVar1S0S89P014P017P015P037(0)='1' AND  B(10)='1' )then
          cVar2S0S89P034nsss(0) <='1';
          else
          cVar2S0S89P034nsss(0) <='0';
          end if;
        if(cVar1S1S89P014P017P015P037(0)='1' AND  B(10)='0' AND B(14)='0' )then
          cVar2S1S89N034P026nsss(0) <='1';
          else
          cVar2S1S89N034P026nsss(0) <='0';
          end if;
        if(cVar1S2S89P014P017P015P037(0)='1' AND  B(10)='0' AND B(14)='1' AND A(10)='0' )then
          cVar2S2S89N034P026P018nsss(0) <='1';
          else
          cVar2S2S89N034P026P018nsss(0) <='0';
          end if;
        if(cVar1S3S89P014P017P015N037(0)='1' AND  B( 9)='1' )then
          cVar2S3S89P036nsss(0) <='1';
          else
          cVar2S3S89P036nsss(0) <='0';
          end if;
        if(cVar1S4S89P014P017P015N037(0)='1' AND  B( 9)='0' AND B(17)='1' AND A( 5)='0' )then
          cVar2S4S89N036P020P009nsss(0) <='1';
          else
          cVar2S4S89N036P020P009nsss(0) <='0';
          end if;
        if(cVar1S5S89P014P017P015N037(0)='1' AND  B( 9)='0' AND B(17)='0' AND D( 7)='1' )then
          cVar2S5S89N036N020P038nsss(0) <='1';
          else
          cVar2S5S89N036N020P038nsss(0) <='0';
          end if;
        if(cVar1S6S89P014P017P015P030(0)='1' AND  E( 1)='1' )then
          cVar2S6S89P064nsss(0) <='1';
          else
          cVar2S6S89P064nsss(0) <='0';
          end if;
        if(cVar1S7S89P014P017P015P030(0)='1' AND  E( 1)='0' AND D( 0)='1' )then
          cVar2S7S89N064P066nsss(0) <='1';
          else
          cVar2S7S89N064P066nsss(0) <='0';
          end if;
        if(cVar1S8S89P014P017P015P030(0)='1' AND  E( 1)='0' AND D( 0)='0' AND E( 3)='1' )then
          cVar2S8S89N064N066P056nsss(0) <='1';
          else
          cVar2S8S89N064N066P056nsss(0) <='0';
          end if;
        if(cVar1S9S89P014P017P015N030(0)='1' AND  E( 1)='0' AND E(15)='0' )then
          cVar2S9S89P064P041nsss(0) <='1';
          else
          cVar2S9S89P064P041nsss(0) <='0';
          end if;
        if(cVar1S10S89P014P017P015N030(0)='1' AND  E( 1)='1' AND E( 4)='1' )then
          cVar2S10S89P064P052nsss(0) <='1';
          else
          cVar2S10S89P064P052nsss(0) <='0';
          end if;
        if(cVar1S11S89P014N017P044P015(0)='1' AND  D( 5)='1' )then
          cVar2S11S89P046nsss(0) <='1';
          else
          cVar2S11S89P046nsss(0) <='0';
          end if;
        if(cVar1S12S89P014N017P044P015(0)='1' AND  D( 5)='0' AND B( 2)='1' )then
          cVar2S12S89N046P033nsss(0) <='1';
          else
          cVar2S12S89N046P033nsss(0) <='0';
          end if;
        if(cVar1S13S89P014N017P044P015(0)='1' AND  D( 5)='0' AND B( 2)='0' AND A(10)='1' )then
          cVar2S13S89N046N033P018nsss(0) <='1';
          else
          cVar2S13S89N046N033P018nsss(0) <='0';
          end if;
        if(cVar1S14S89P014N017P044N015(0)='1' AND  B( 4)='1' )then
          cVar2S14S89P029nsss(0) <='1';
          else
          cVar2S14S89P029nsss(0) <='0';
          end if;
        if(cVar1S15S89P014N017P044N015(0)='1' AND  B( 4)='0' AND D( 5)='0' )then
          cVar2S15S89N029P046nsss(0) <='1';
          else
          cVar2S15S89N029P046nsss(0) <='0';
          end if;
        if(cVar1S16S89P014N017P044N015(0)='1' AND  B( 4)='0' AND D( 5)='1' AND B( 0)='1' )then
          cVar2S16S89N029P046P037nsss(0) <='1';
          else
          cVar2S16S89N029P046P037nsss(0) <='0';
          end if;
        if(cVar1S17S89P014N017N044P027(0)='1' AND  B( 7)='0' AND A(16)='1' )then
          cVar2S17S89P023P006nsss(0) <='1';
          else
          cVar2S17S89P023P006nsss(0) <='0';
          end if;
        if(cVar1S18S89P014N017N044P027(0)='1' AND  B( 7)='0' AND A(16)='0' AND B( 9)='0' )then
          cVar2S18S89P023N006P036nsss(0) <='1';
          else
          cVar2S18S89P023N006P036nsss(0) <='0';
          end if;
        if(cVar1S19S89P014N017N044N027(0)='1' AND  E( 5)='0' AND D( 5)='0' AND A(17)='0' )then
          cVar2S19S89P048P046P004nsss(0) <='1';
          else
          cVar2S19S89P048P046P004nsss(0) <='0';
          end if;
        if(cVar1S20S89P014N017N044N027(0)='1' AND  E( 5)='1' AND D( 1)='0' AND E( 7)='0' )then
          cVar2S20S89P048P062P040nsss(0) <='1';
          else
          cVar2S20S89P048P062P040nsss(0) <='0';
          end if;
        if(cVar1S21S89P014P021P012P040(0)='1' AND  B( 5)='0' AND B(11)='1' )then
          cVar2S21S89P027P032nsss(0) <='1';
          else
          cVar2S21S89P027P032nsss(0) <='0';
          end if;
        if(cVar1S22S89P014P021P012P040(0)='1' AND  B( 5)='0' AND B(11)='0' AND D( 1)='1' )then
          cVar2S22S89P027N032P062nsss(0) <='1';
          else
          cVar2S22S89P027N032P062nsss(0) <='0';
          end if;
        if(cVar1S23S89P014P021P012P040(0)='1' AND  B( 5)='1' AND D(12)='1' )then
          cVar2S23S89P027P051nsss(0) <='1';
          else
          cVar2S23S89P027P051nsss(0) <='0';
          end if;
        if(cVar1S24S89P014P021P012P040(0)='1' AND  B( 5)='1' AND D(12)='0' AND E( 5)='1' )then
          cVar2S24S89P027N051P048nsss(0) <='1';
          else
          cVar2S24S89P027N051P048nsss(0) <='0';
          end if;
        if(cVar1S25S89P014P021P012P040(0)='1' AND  A(14)='0' AND A( 0)='0' AND A(10)='1' )then
          cVar2S25S89P010P019P018nsss(0) <='1';
          else
          cVar2S25S89P010P019P018nsss(0) <='0';
          end if;
        if(cVar1S26S89P014P021P012P039(0)='1' AND  B( 9)='1' AND E( 3)='1' )then
          cVar2S26S89P036P056nsss(0) <='1';
          else
          cVar2S26S89P036P056nsss(0) <='0';
          end if;
        if(cVar1S27S89P014P021P012P039(0)='1' AND  B( 9)='1' AND E( 3)='0' AND B( 3)='0' )then
          cVar2S27S89P036N056P031nsss(0) <='1';
          else
          cVar2S27S89P036N056P031nsss(0) <='0';
          end if;
        if(cVar1S28S89P014P021P012P039(0)='1' AND  B( 9)='0' AND A(11)='1' AND A( 0)='1' )then
          cVar2S28S89N036P016P019nsss(0) <='1';
          else
          cVar2S28S89N036P016P019nsss(0) <='0';
          end if;
        if(cVar1S29S89P014P021P012P039(0)='1' AND  B( 9)='0' AND A(11)='0' AND B(12)='1' )then
          cVar2S29S89N036N016P030nsss(0) <='1';
          else
          cVar2S29S89N036N016P030nsss(0) <='0';
          end if;
        if(cVar1S30S89P014P021P026P037(0)='1' AND  B( 9)='1' )then
          cVar2S30S89P036nsss(0) <='1';
          else
          cVar2S30S89P036nsss(0) <='0';
          end if;
        if(cVar1S31S89P014P021P026P037(0)='1' AND  B( 9)='0' AND A(10)='0' AND A( 0)='1' )then
          cVar2S31S89N036P018P019nsss(0) <='1';
          else
          cVar2S31S89N036P018P019nsss(0) <='0';
          end if;
        if(cVar1S32S89P014P021P026N037(0)='1' AND  E( 2)='1' )then
          cVar2S32S89P060nsss(0) <='1';
          else
          cVar2S32S89P060nsss(0) <='0';
          end if;
        if(cVar1S0S90P017P014P019P042(0)='1' AND  B( 9)='1' )then
          cVar2S0S90P036nsss(0) <='1';
          else
          cVar2S0S90P036nsss(0) <='0';
          end if;
        if(cVar1S1S90P017P014P019P042(0)='1' AND  B( 9)='0' AND B( 1)='1' )then
          cVar2S1S90N036P035nsss(0) <='1';
          else
          cVar2S1S90N036P035nsss(0) <='0';
          end if;
        if(cVar1S2S90P017P014P019P042(0)='1' AND  B( 9)='0' AND B( 1)='0' AND A( 2)='1' )then
          cVar2S2S90N036N035P015nsss(0) <='1';
          else
          cVar2S2S90N036N035P015nsss(0) <='0';
          end if;
        if(cVar1S3S90P017P014P019N042(0)='1' AND  A(19)='1' AND B(10)='1' )then
          cVar2S3S90P000P034nsss(0) <='1';
          else
          cVar2S3S90P000P034nsss(0) <='0';
          end if;
        if(cVar1S4S90P017P014P019N042(0)='1' AND  A(19)='1' AND B(10)='0' AND E( 0)='1' )then
          cVar2S4S90P000N034P068nsss(0) <='1';
          else
          cVar2S4S90P000N034P068nsss(0) <='0';
          end if;
        if(cVar1S5S90P017P014P019N042(0)='1' AND  A(19)='0' AND A(17)='0' )then
          cVar2S5S90N000P004nsss(0) <='1';
          else
          cVar2S5S90N000P004nsss(0) <='0';
          end if;
        if(cVar1S6S90P017P014P019P042(0)='1' AND  B( 7)='0' AND B( 5)='1' )then
          cVar2S6S90P023P027nsss(0) <='1';
          else
          cVar2S6S90P023P027nsss(0) <='0';
          end if;
        if(cVar1S7S90P017P014P019P042(0)='1' AND  B( 7)='0' AND B( 5)='0' AND E( 0)='1' )then
          cVar2S7S90P023N027P068nsss(0) <='1';
          else
          cVar2S7S90P023N027P068nsss(0) <='0';
          end if;
        if(cVar1S8S90P017P014P019P042(0)='1' AND  B( 7)='1' )then
          cVar2S8S90P023nsss(0) <='1';
          else
          cVar2S8S90P023nsss(0) <='0';
          end if;
        if(cVar1S9S90P017P014P047P024(0)='1' AND  E( 8)='1' AND E( 2)='1' AND B(11)='0' )then
          cVar2S9S90P069P060P032nsss(0) <='1';
          else
          cVar2S9S90P069P060P032nsss(0) <='0';
          end if;
        if(cVar1S10S90P017P014P047P024(0)='1' AND  E( 8)='1' AND E( 2)='0' AND B( 0)='1' )then
          cVar2S10S90P069N060P037nsss(0) <='1';
          else
          cVar2S10S90P069N060P037nsss(0) <='0';
          end if;
        if(cVar1S11S90P017P014P047P024(0)='1' AND  D( 0)='1' AND A( 0)='0' )then
          cVar2S11S90P066P019nsss(0) <='1';
          else
          cVar2S11S90P066P019nsss(0) <='0';
          end if;
        if(cVar1S12S90P017P014P047P024(0)='1' AND  D( 0)='1' AND A( 0)='1' AND A(11)='1' )then
          cVar2S12S90P066P019P016nsss(0) <='1';
          else
          cVar2S12S90P066P019P016nsss(0) <='0';
          end if;
        if(cVar1S13S90P017P014P047P024(0)='1' AND  D( 0)='0' AND A(11)='0' AND A(13)='1' )then
          cVar2S13S90N066P016P012nsss(0) <='1';
          else
          cVar2S13S90N066P016P012nsss(0) <='0';
          end if;
        if(cVar1S15S90N017P068P004P025(0)='1' AND  D( 5)='1' )then
          cVar2S15S90P046nsss(0) <='1';
          else
          cVar2S15S90P046nsss(0) <='0';
          end if;
        if(cVar1S16S90N017P068P004N025(0)='1' AND  E( 7)='1' )then
          cVar2S16S90P040nsss(0) <='1';
          else
          cVar2S16S90P040nsss(0) <='0';
          end if;
        if(cVar1S17S90N017P068P004N025(0)='1' AND  E( 7)='0' AND A(18)='0' AND E( 6)='1' )then
          cVar2S17S90N040P002P044nsss(0) <='1';
          else
          cVar2S17S90N040P002P044nsss(0) <='0';
          end if;
        if(cVar1S18S90N017P068P004N025(0)='1' AND  E( 7)='0' AND A(18)='1' AND A(12)='1' )then
          cVar2S18S90N040P002P014nsss(0) <='1';
          else
          cVar2S18S90N040P002P014nsss(0) <='0';
          end if;
        if(cVar1S19S90N017P068N004P028(0)='1' AND  D( 0)='0' )then
          cVar2S19S90P066nsss(0) <='1';
          else
          cVar2S19S90P066nsss(0) <='0';
          end if;
        if(cVar1S20S90N017P068N004N028(0)='1' AND  D(15)='1' AND D( 0)='0' AND E( 7)='0' )then
          cVar2S20S90P039P066P040nsss(0) <='1';
          else
          cVar2S20S90P039P066P040nsss(0) <='0';
          end if;
        if(cVar1S21S90N017P068N004N028(0)='1' AND  D(15)='0' AND B(17)='1' AND D(14)='1' )then
          cVar2S21S90N039P020P043nsss(0) <='1';
          else
          cVar2S21S90N039P020P043nsss(0) <='0';
          end if;
        if(cVar1S22S90N017P068P064P062(0)='1' AND  D(12)='1' AND D(11)='0' AND A(10)='1' )then
          cVar2S22S90P051P055P018nsss(0) <='1';
          else
          cVar2S22S90P051P055P018nsss(0) <='0';
          end if;
        if(cVar1S23S90N017P068P064P062(0)='1' AND  D(12)='0' AND D( 6)='1' )then
          cVar2S23S90N051P042nsss(0) <='1';
          else
          cVar2S23S90N051P042nsss(0) <='0';
          end if;
        if(cVar1S24S90N017P068P064P062(0)='1' AND  B(11)='1' )then
          cVar2S24S90P032nsss(0) <='1';
          else
          cVar2S24S90P032nsss(0) <='0';
          end if;
        if(cVar1S25S90N017P068P064P062(0)='1' AND  B(11)='0' AND A(15)='1' AND A( 2)='0' )then
          cVar2S25S90N032P008P015nsss(0) <='1';
          else
          cVar2S25S90N032P008P015nsss(0) <='0';
          end if;
        if(cVar1S26S90N017P068P064P019(0)='1' AND  D( 1)='1' AND D( 0)='1' AND A(10)='0' )then
          cVar2S26S90P062P066P018nsss(0) <='1';
          else
          cVar2S26S90P062P066P018nsss(0) <='0';
          end if;
        if(cVar1S27S90N017P068P064P019(0)='1' AND  D( 1)='0' AND E( 9)='0' AND B( 0)='1' )then
          cVar2S27S90N062P065P037nsss(0) <='1';
          else
          cVar2S27S90N062P065P037nsss(0) <='0';
          end if;
        if(cVar1S28S90N017P068P064N019(0)='1' AND  A( 2)='1' AND B(10)='0' AND E( 9)='1' )then
          cVar2S28S90P015P034P065nsss(0) <='1';
          else
          cVar2S28S90P015P034P065nsss(0) <='0';
          end if;
        if(cVar1S29S90N017P068P064N019(0)='1' AND  A( 2)='0' AND E(11)='0' AND D( 3)='1' )then
          cVar2S29S90N015N057P054nsss(0) <='1';
          else
          cVar2S29S90N015N057P054nsss(0) <='0';
          end if;
        if(cVar1S0S91P017P068P010P004(0)='1' AND  B( 6)='1' AND D( 5)='1' )then
          cVar2S0S91P025P046nsss(0) <='1';
          else
          cVar2S0S91P025P046nsss(0) <='0';
          end if;
        if(cVar1S1S91P017P068P010P004(0)='1' AND  B( 6)='0' AND B( 1)='0' )then
          cVar2S1S91N025P035nsss(0) <='1';
          else
          cVar2S1S91N025P035nsss(0) <='0';
          end if;
        if(cVar1S2S91P017P068P010P004(0)='1' AND  B( 6)='0' AND B( 1)='1' AND A(11)='1' )then
          cVar2S2S91N025P035P016nsss(0) <='1';
          else
          cVar2S2S91N025P035P016nsss(0) <='0';
          end if;
        if(cVar1S3S91P017P068P010N004(0)='1' AND  A(16)='1' AND B( 5)='1' )then
          cVar2S3S91P006P027nsss(0) <='1';
          else
          cVar2S3S91P006P027nsss(0) <='0';
          end if;
        if(cVar1S4S91P017P068P010N004(0)='1' AND  A(16)='1' AND B( 5)='0' AND D(13)='1' )then
          cVar2S4S91P006N027P047nsss(0) <='1';
          else
          cVar2S4S91P006N027P047nsss(0) <='0';
          end if;
        if(cVar1S5S91P017P068P010N004(0)='1' AND  A(16)='0' )then
          cVar2S5S91N006psss(0) <='1';
          else
          cVar2S5S91N006psss(0) <='0';
          end if;
        if(cVar1S6S91P017P068P010P021(0)='1' AND  A(19)='0' AND B(17)='0' AND A(15)='0' )then
          cVar2S6S91P000P020P008nsss(0) <='1';
          else
          cVar2S6S91P000P020P008nsss(0) <='0';
          end if;
        if(cVar1S7S91P017P068P010P021(0)='1' AND  A( 2)='1' AND A( 0)='0' )then
          cVar2S7S91P015P019nsss(0) <='1';
          else
          cVar2S7S91P015P019nsss(0) <='0';
          end if;
        if(cVar1S8S91P017P068P010P021(0)='1' AND  A( 2)='0' AND A( 5)='0' AND A( 8)='1' )then
          cVar2S8S91N015P009P003nsss(0) <='1';
          else
          cVar2S8S91N015P009P003nsss(0) <='0';
          end if;
        if(cVar1S9S91P017P068P064P062(0)='1' AND  D( 2)='0' )then
          cVar2S9S91P058nsss(0) <='1';
          else
          cVar2S9S91P058nsss(0) <='0';
          end if;
        if(cVar1S10S91P017P068P064P062(0)='1' AND  D( 2)='1' AND D( 0)='1' AND E(10)='0' )then
          cVar2S10S91P058P066P061nsss(0) <='1';
          else
          cVar2S10S91P058P066P061nsss(0) <='0';
          end if;
        if(cVar1S11S91P017P068P064P062(0)='1' AND  D( 2)='1' AND D( 0)='0' AND A(10)='0' )then
          cVar2S11S91P058N066P018nsss(0) <='1';
          else
          cVar2S11S91P058N066P018nsss(0) <='0';
          end if;
        if(cVar1S12S91P017P068P064P062(0)='1' AND  E( 2)='1' AND E( 8)='0' AND A( 3)='0' )then
          cVar2S12S91P060P069P013nsss(0) <='1';
          else
          cVar2S12S91P060P069P013nsss(0) <='0';
          end if;
        if(cVar1S13S91P017P068P064P062(0)='1' AND  E( 2)='1' AND E( 8)='1' AND A(12)='0' )then
          cVar2S13S91P060P069P014nsss(0) <='1';
          else
          cVar2S13S91P060P069P014nsss(0) <='0';
          end if;
        if(cVar1S14S91P017P068P064P062(0)='1' AND  E( 2)='0' AND A(15)='1' AND B( 0)='1' )then
          cVar2S14S91N060P008P037nsss(0) <='1';
          else
          cVar2S14S91N060P008P037nsss(0) <='0';
          end if;
        if(cVar1S15S91P017P068P064P062(0)='1' AND  E( 2)='0' AND A(15)='0' AND A( 5)='1' )then
          cVar2S15S91N060N008P009nsss(0) <='1';
          else
          cVar2S15S91N060N008P009nsss(0) <='0';
          end if;
        if(cVar1S16S91P017P068P064P019(0)='1' AND  D( 1)='1' AND D( 0)='1' AND B( 0)='0' )then
          cVar2S16S91P062P066P037nsss(0) <='1';
          else
          cVar2S16S91P062P066P037nsss(0) <='0';
          end if;
        if(cVar1S17S91P017P068P064P019(0)='1' AND  D( 1)='0' AND A(12)='1' AND A(10)='0' )then
          cVar2S17S91N062P014P018nsss(0) <='1';
          else
          cVar2S17S91N062P014P018nsss(0) <='0';
          end if;
        if(cVar1S18S91P017P068P064N019(0)='1' AND  A( 2)='1' AND B(10)='0' AND E( 8)='1' )then
          cVar2S18S91P015P034P069nsss(0) <='1';
          else
          cVar2S18S91P015P034P069nsss(0) <='0';
          end if;
        if(cVar1S19S91P017P068P064N019(0)='1' AND  A( 2)='0' AND E(11)='0' AND D( 3)='1' )then
          cVar2S19S91N015N057P054nsss(0) <='1';
          else
          cVar2S19S91N015N057P054nsss(0) <='0';
          end if;
        if(cVar1S20S91P017P044P060P010(0)='1' AND  D( 4)='0' )then
          cVar2S20S91P050nsss(0) <='1';
          else
          cVar2S20S91P050nsss(0) <='0';
          end if;
        if(cVar1S21S91P017P044P060P010(0)='1' AND  A( 2)='1' )then
          cVar2S21S91P015nsss(0) <='1';
          else
          cVar2S21S91P015nsss(0) <='0';
          end if;
        if(cVar1S22S91P017N044P023P042(0)='1' AND  A(18)='0' AND D( 7)='0' AND E(10)='1' )then
          cVar2S22S91P002P038P061nsss(0) <='1';
          else
          cVar2S22S91P002P038P061nsss(0) <='0';
          end if;
        if(cVar1S23S91P017N044P023P042(0)='1' AND  A(18)='0' AND D( 7)='1' AND A(17)='1' )then
          cVar2S23S91P002P038P004nsss(0) <='1';
          else
          cVar2S23S91P002P038P004nsss(0) <='0';
          end if;
        if(cVar1S24S91P017N044P023P042(0)='1' AND  A(18)='1' AND A( 3)='1' AND B( 9)='1' )then
          cVar2S24S91P002P013P036nsss(0) <='1';
          else
          cVar2S24S91P002P013P036nsss(0) <='0';
          end if;
        if(cVar1S25S91P017N044P023P042(0)='1' AND  A(18)='1' AND A( 3)='0' AND D( 7)='1' )then
          cVar2S25S91P002N013P038nsss(0) <='1';
          else
          cVar2S25S91P002N013P038nsss(0) <='0';
          end if;
        if(cVar1S26S91P017N044P023P042(0)='1' AND  A(17)='1' )then
          cVar2S26S91P004nsss(0) <='1';
          else
          cVar2S26S91P004nsss(0) <='0';
          end if;
        if(cVar1S27S91P017N044P023P042(0)='1' AND  A(17)='0' AND A( 0)='0' AND B( 1)='1' )then
          cVar2S27S91N004P019P035nsss(0) <='1';
          else
          cVar2S27S91N004P019P035nsss(0) <='0';
          end if;
        if(cVar1S29S91P017N044P023N065(0)='1' AND  A(14)='0' AND B(16)='0' AND A(11)='1' )then
          cVar2S29S91P010P022P016nsss(0) <='1';
          else
          cVar2S29S91P010P022P016nsss(0) <='0';
          end if;
        if(cVar1S0S92P017P059P061P013(0)='1' AND  A(18)='0' AND E(15)='0' )then
          cVar2S0S92P002P041nsss(0) <='1';
          else
          cVar2S0S92P002P041nsss(0) <='0';
          end if;
        if(cVar1S1S92P017P059P061P013(0)='1' AND  A(18)='0' AND E(15)='1' AND A(15)='1' )then
          cVar2S1S92P002P041P008nsss(0) <='1';
          else
          cVar2S1S92P002P041P008nsss(0) <='0';
          end if;
        if(cVar1S2S92P017P059P061P013(0)='1' AND  A(18)='1' AND E( 7)='1' )then
          cVar2S2S92P002P040nsss(0) <='1';
          else
          cVar2S2S92P002P040nsss(0) <='0';
          end if;
        if(cVar1S3S92P017P059P061P013(0)='1' AND  A(18)='1' AND E( 7)='0' AND E( 1)='1' )then
          cVar2S3S92P002N040P064nsss(0) <='1';
          else
          cVar2S3S92P002N040P064nsss(0) <='0';
          end if;
        if(cVar1S4S92P017P059P061P013(0)='1' AND  D( 2)='1' AND D( 0)='0' )then
          cVar2S4S92P058P066nsss(0) <='1';
          else
          cVar2S4S92P058P066nsss(0) <='0';
          end if;
        if(cVar1S5S92P017P059P061P013(0)='1' AND  D( 2)='1' AND D( 0)='1' AND B( 9)='1' )then
          cVar2S5S92P058P066P036nsss(0) <='1';
          else
          cVar2S5S92P058P066P036nsss(0) <='0';
          end if;
        if(cVar1S6S92P017P059P061P013(0)='1' AND  D( 2)='0' AND A(18)='1' AND A(11)='0' )then
          cVar2S6S92N058P002P016nsss(0) <='1';
          else
          cVar2S6S92N058P002P016nsss(0) <='0';
          end if;
        if(cVar1S7S92P017P059P061P013(0)='1' AND  D( 2)='0' AND A(18)='0' AND E( 4)='1' )then
          cVar2S7S92N058N002P052nsss(0) <='1';
          else
          cVar2S7S92N058N002P052nsss(0) <='0';
          end if;
        if(cVar1S8S92P017P059P061P066(0)='1' AND  A( 0)='0' )then
          cVar2S8S92P019nsss(0) <='1';
          else
          cVar2S8S92P019nsss(0) <='0';
          end if;
        if(cVar1S9S92P017P059P061P066(0)='1' AND  A( 0)='1' AND A(11)='1' )then
          cVar2S9S92P019P016nsss(0) <='1';
          else
          cVar2S9S92P019P016nsss(0) <='0';
          end if;
        if(cVar1S10S92P017P059P061N066(0)='1' AND  B(10)='1' AND A(10)='0' )then
          cVar2S10S92P034P018nsss(0) <='1';
          else
          cVar2S10S92P034P018nsss(0) <='0';
          end if;
        if(cVar1S11S92P017P059P030P012(0)='1' AND  E(11)='1' )then
          cVar2S11S92P057nsss(0) <='1';
          else
          cVar2S11S92P057nsss(0) <='0';
          end if;
        if(cVar1S12S92P017P059P030P012(0)='1' AND  E(11)='0' AND A(10)='0' )then
          cVar2S12S92N057P018nsss(0) <='1';
          else
          cVar2S12S92N057P018nsss(0) <='0';
          end if;
        if(cVar1S13S92P017P059P030P012(0)='1' AND  A( 0)='1' )then
          cVar2S13S92P019nsss(0) <='1';
          else
          cVar2S13S92P019nsss(0) <='0';
          end if;
        if(cVar1S14S92P017P059N030P055(0)='1' AND  E(10)='1' AND D( 2)='0' AND B(10)='1' )then
          cVar2S14S92P061P058P034nsss(0) <='1';
          else
          cVar2S14S92P061P058P034nsss(0) <='0';
          end if;
        if(cVar1S15S92P017P059N030P055(0)='1' AND  E(10)='1' AND D( 2)='1' AND A(12)='0' )then
          cVar2S15S92P061P058P014nsss(0) <='1';
          else
          cVar2S15S92P061P058P014nsss(0) <='0';
          end if;
        if(cVar1S16S92P017P059N030P055(0)='1' AND  E(10)='0' AND D( 1)='1' AND A( 0)='0' )then
          cVar2S16S92N061P062P019nsss(0) <='1';
          else
          cVar2S16S92N061P062P019nsss(0) <='0';
          end if;
        if(cVar1S17S92P017P059N030P055(0)='1' AND  E(10)='0' AND D( 1)='0' AND E( 3)='1' )then
          cVar2S17S92N061N062P056nsss(0) <='1';
          else
          cVar2S17S92N061N062P056nsss(0) <='0';
          end if;
        if(cVar1S18S92P017P059N030P055(0)='1' AND  E(10)='0' )then
          cVar2S18S92P061nsss(0) <='1';
          else
          cVar2S18S92P061nsss(0) <='0';
          end if;
        if(cVar1S20S92N017P006P027N048(0)='1' AND  E( 4)='1' )then
          cVar2S20S92P052nsss(0) <='1';
          else
          cVar2S20S92P052nsss(0) <='0';
          end if;
        if(cVar1S21S92N017P006P027N048(0)='1' AND  E( 4)='0' AND A( 4)='1' )then
          cVar2S21S92N052P011nsss(0) <='1';
          else
          cVar2S21S92N052P011nsss(0) <='0';
          end if;
        if(cVar1S22S92N017P006N027P015(0)='1' AND  D( 9)='0' )then
          cVar2S22S92P063nsss(0) <='1';
          else
          cVar2S22S92P063nsss(0) <='0';
          end if;
        if(cVar1S23S92N017P006N027P015(0)='1' AND  D( 9)='1' AND B( 0)='0' AND E( 9)='1' )then
          cVar2S23S92P063P037P065nsss(0) <='1';
          else
          cVar2S23S92P063P037P065nsss(0) <='0';
          end if;
        if(cVar1S24S92N017P006N027N015(0)='1' AND  D( 3)='0' AND A(14)='0' AND D(13)='1' )then
          cVar2S24S92P054P010P047nsss(0) <='1';
          else
          cVar2S24S92P054P010P047nsss(0) <='0';
          end if;
        if(cVar1S25S92N017P006N027N015(0)='1' AND  D( 3)='0' AND A(14)='1' AND D(14)='1' )then
          cVar2S25S92P054P010P043nsss(0) <='1';
          else
          cVar2S25S92P054P010P043nsss(0) <='0';
          end if;
        if(cVar1S26S92N017N006P030P028(0)='1' AND  E(10)='1' AND A( 3)='1' )then
          cVar2S26S92P061P013nsss(0) <='1';
          else
          cVar2S26S92P061P013nsss(0) <='0';
          end if;
        if(cVar1S27S92N017N006P030P028(0)='1' AND  E(10)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar2S27S92P061N013P011nsss(0) <='1';
          else
          cVar2S27S92P061N013P011nsss(0) <='0';
          end if;
        if(cVar1S28S92N017N006P030P028(0)='1' AND  E(10)='0' AND B(11)='0' )then
          cVar2S28S92N061P032nsss(0) <='1';
          else
          cVar2S28S92N061P032nsss(0) <='0';
          end if;
        if(cVar1S29S92N017N006P030P028(0)='1' AND  E(12)='1' )then
          cVar2S29S92P053nsss(0) <='1';
          else
          cVar2S29S92P053nsss(0) <='0';
          end if;
        if(cVar1S30S92N017N006P030P028(0)='1' AND  E(12)='0' AND A( 3)='0' AND A(10)='0' )then
          cVar2S30S92N053P013P018nsss(0) <='1';
          else
          cVar2S30S92N053P013P018nsss(0) <='0';
          end if;
        if(cVar1S31S92N017N006N030P014(0)='1' AND  B( 8)='0' AND B( 9)='1' AND E(10)='0' )then
          cVar2S31S92P021P036P061nsss(0) <='1';
          else
          cVar2S31S92P021P036P061nsss(0) <='0';
          end if;
        if(cVar1S32S92N017N006N030P014(0)='1' AND  B( 8)='0' AND B( 9)='0' AND E(10)='1' )then
          cVar2S32S92P021N036P061nsss(0) <='1';
          else
          cVar2S32S92P021N036P061nsss(0) <='0';
          end if;
        if(cVar1S33S92N017N006N030P014(0)='1' AND  B( 8)='1' AND A(13)='0' AND B( 9)='1' )then
          cVar2S33S92P021P012P036nsss(0) <='1';
          else
          cVar2S33S92P021P012P036nsss(0) <='0';
          end if;
        if(cVar1S34S92N017N006N030N014(0)='1' AND  E(15)='1' AND A( 7)='1' )then
          cVar2S34S92P041P005nsss(0) <='1';
          else
          cVar2S34S92P041P005nsss(0) <='0';
          end if;
        if(cVar1S35S92N017N006N030N014(0)='1' AND  E(15)='1' AND A( 7)='0' AND E( 8)='1' )then
          cVar2S35S92P041N005P069nsss(0) <='1';
          else
          cVar2S35S92P041N005P069nsss(0) <='0';
          end if;
        if(cVar1S0S93P017P030P014P010(0)='1' AND  A(16)='1' AND A( 3)='1' )then
          cVar2S0S93P006P013nsss(0) <='1';
          else
          cVar2S0S93P006P013nsss(0) <='0';
          end if;
        if(cVar1S1S93P017P030P014P010(0)='1' AND  A(16)='1' AND A( 3)='0' AND E( 0)='0' )then
          cVar2S1S93P006N013P068nsss(0) <='1';
          else
          cVar2S1S93P006N013P068nsss(0) <='0';
          end if;
        if(cVar1S2S93P017P030P014P010(0)='1' AND  A(16)='0' AND D( 3)='0' AND A( 3)='0' )then
          cVar2S2S93N006P054P013nsss(0) <='1';
          else
          cVar2S2S93N006P054P013nsss(0) <='0';
          end if;
        if(cVar1S3S93P017P030P014P010(0)='1' AND  A(16)='0' AND D( 3)='1' AND A( 3)='1' )then
          cVar2S3S93N006P054P013nsss(0) <='1';
          else
          cVar2S3S93N006P054P013nsss(0) <='0';
          end if;
        if(cVar1S4S93P017P030P014P010(0)='1' AND  D( 3)='1' AND D( 4)='0' )then
          cVar2S4S93P054P050nsss(0) <='1';
          else
          cVar2S4S93P054P050nsss(0) <='0';
          end if;
        if(cVar1S5S93P017P030P014P010(0)='1' AND  D( 3)='0' AND D( 4)='1' )then
          cVar2S5S93N054P050nsss(0) <='1';
          else
          cVar2S5S93N054P050nsss(0) <='0';
          end if;
        if(cVar1S6S93P017P030P014P010(0)='1' AND  D( 3)='0' AND D( 4)='0' AND B(13)='1' )then
          cVar2S6S93N054N050P028nsss(0) <='1';
          else
          cVar2S6S93N054N050P028nsss(0) <='0';
          end if;
        if(cVar1S7S93P017P030P014P021(0)='1' AND  B( 0)='1' AND D(12)='1' AND A(13)='0' )then
          cVar2S7S93P037P051P012nsss(0) <='1';
          else
          cVar2S7S93P037P051P012nsss(0) <='0';
          end if;
        if(cVar1S8S93P017P030P014P021(0)='1' AND  B( 0)='1' AND D(12)='0' AND D(14)='0' )then
          cVar2S8S93P037N051P043nsss(0) <='1';
          else
          cVar2S8S93P037N051P043nsss(0) <='0';
          end if;
        if(cVar1S9S93P017P030P014P021(0)='1' AND  B( 0)='0' AND E( 0)='0' AND E(10)='0' )then
          cVar2S9S93N037P068P061nsss(0) <='1';
          else
          cVar2S9S93N037P068P061nsss(0) <='0';
          end if;
        if(cVar1S10S93P017P030P014P021(0)='1' AND  B( 0)='0' AND E( 0)='1' AND A( 7)='1' )then
          cVar2S10S93N037P068P005nsss(0) <='1';
          else
          cVar2S10S93N037P068P005nsss(0) <='0';
          end if;
        if(cVar1S11S93P017P030P014P021(0)='1' AND  A( 3)='0' AND B( 0)='1' AND A( 0)='1' )then
          cVar2S11S93P013P037P019nsss(0) <='1';
          else
          cVar2S11S93P013P037P019nsss(0) <='0';
          end if;
        if(cVar1S13S93P017P030P061N013(0)='1' AND  A(11)='0' AND D(11)='1' )then
          cVar2S13S93P016P055nsss(0) <='1';
          else
          cVar2S13S93P016P055nsss(0) <='0';
          end if;
        if(cVar1S14S93P017P030P061N013(0)='1' AND  A(11)='0' AND D(11)='0' AND B( 0)='1' )then
          cVar2S14S93P016N055P037nsss(0) <='1';
          else
          cVar2S14S93P016N055P037nsss(0) <='0';
          end if;
        if(cVar1S15S93P017P030N061P032(0)='1' AND  B( 3)='0' AND E( 5)='1' )then
          cVar2S15S93P031P048nsss(0) <='1';
          else
          cVar2S15S93P031P048nsss(0) <='0';
          end if;
        if(cVar1S16S93P017P030N061P032(0)='1' AND  B( 3)='1' AND B( 1)='0' AND E( 8)='1' )then
          cVar2S16S93P031P035P069nsss(0) <='1';
          else
          cVar2S16S93P031P035P069nsss(0) <='0';
          end if;
        if(cVar1S17S93P017P030N061P032(0)='1' AND  A(13)='0' AND A(12)='0' )then
          cVar2S17S93P012P014nsss(0) <='1';
          else
          cVar2S17S93P012P014nsss(0) <='0';
          end if;
        if(cVar1S18S93P017P013P003P008(0)='1' AND  E(11)='1' AND B( 3)='1' )then
          cVar2S18S93P057P031nsss(0) <='1';
          else
          cVar2S18S93P057P031nsss(0) <='0';
          end if;
        if(cVar1S19S93P017P013P003P008(0)='1' AND  E(11)='1' AND B( 3)='0' AND B(12)='1' )then
          cVar2S19S93P057N031P030nsss(0) <='1';
          else
          cVar2S19S93P057N031P030nsss(0) <='0';
          end if;
        if(cVar1S20S93P017P013P003P008(0)='1' AND  E(11)='0' AND B( 2)='1' AND B( 3)='0' )then
          cVar2S20S93N057P033P031nsss(0) <='1';
          else
          cVar2S20S93N057P033P031nsss(0) <='0';
          end if;
        if(cVar1S21S93P017P013P003P008(0)='1' AND  E(11)='0' AND B( 2)='0' AND B(11)='1' )then
          cVar2S21S93N057N033P032nsss(0) <='1';
          else
          cVar2S21S93N057N033P032nsss(0) <='0';
          end if;
        if(cVar1S22S93P017P013P003P008(0)='1' AND  E( 4)='1' )then
          cVar2S22S93P052nsss(0) <='1';
          else
          cVar2S22S93P052nsss(0) <='0';
          end if;
        if(cVar1S23S93P017P013P003P008(0)='1' AND  E( 4)='0' AND B( 5)='1' )then
          cVar2S23S93N052P027nsss(0) <='1';
          else
          cVar2S23S93N052P027nsss(0) <='0';
          end if;
        if(cVar1S24S93P017P013P003P053(0)='1' AND  B(14)='0' AND D( 4)='1' )then
          cVar2S24S93P026P050nsss(0) <='1';
          else
          cVar2S24S93P026P050nsss(0) <='0';
          end if;
        if(cVar1S25S93P017P013P003P053(0)='1' AND  B(14)='0' AND D( 4)='0' AND E(14)='1' )then
          cVar2S25S93P026N050P045nsss(0) <='1';
          else
          cVar2S25S93P026N050P045nsss(0) <='0';
          end if;
        if(cVar1S26S93P017N013P003P068(0)='1' AND  A(15)='1' )then
          cVar2S26S93P008nsss(0) <='1';
          else
          cVar2S26S93P008nsss(0) <='0';
          end if;
        if(cVar1S27S93P017N013P003P068(0)='1' AND  A(15)='0' AND A( 7)='1' )then
          cVar2S27S93N008P005nsss(0) <='1';
          else
          cVar2S27S93N008P005nsss(0) <='0';
          end if;
        if(cVar1S28S93P017N013P003P068(0)='1' AND  A(15)='0' AND A( 7)='0' AND A( 6)='1' )then
          cVar2S28S93N008N005P007nsss(0) <='1';
          else
          cVar2S28S93N008N005P007nsss(0) <='0';
          end if;
        if(cVar1S29S93P017N013P003N068(0)='1' AND  A(15)='0' AND B( 1)='1' AND E( 1)='1' )then
          cVar2S29S93P008P035P064nsss(0) <='1';
          else
          cVar2S29S93P008P035P064nsss(0) <='0';
          end if;
        if(cVar1S30S93P017N013P003N068(0)='1' AND  A(15)='1' AND D( 8)='0' AND A(10)='0' )then
          cVar2S30S93P008P067P018nsss(0) <='1';
          else
          cVar2S30S93P008P067P018nsss(0) <='0';
          end if;
        if(cVar1S31S93P017N013N003P002(0)='1' AND  E( 0)='0' AND B(16)='1' AND A( 2)='0' )then
          cVar2S31S93P068P022P015nsss(0) <='1';
          else
          cVar2S31S93P068P022P015nsss(0) <='0';
          end if;
        if(cVar1S32S93P017N013N003P002(0)='1' AND  E( 0)='1' AND B(16)='0' AND A(10)='0' )then
          cVar2S32S93P068P022P018nsss(0) <='1';
          else
          cVar2S32S93P068P022P018nsss(0) <='0';
          end if;
        if(cVar1S33S93P017N013N003P002(0)='1' AND  E( 7)='1' )then
          cVar2S33S93P040nsss(0) <='1';
          else
          cVar2S33S93P040nsss(0) <='0';
          end if;
        if(cVar1S34S93P017N013N003P002(0)='1' AND  E( 7)='0' AND B( 0)='1' AND B( 9)='1' )then
          cVar2S34S93N040P037P036nsss(0) <='1';
          else
          cVar2S34S93N040P037P036nsss(0) <='0';
          end if;
        if(cVar1S35S93P017N013N003P002(0)='1' AND  E( 7)='0' AND B( 0)='0' AND B( 1)='1' )then
          cVar2S35S93N040N037P035nsss(0) <='1';
          else
          cVar2S35S93N040N037P035nsss(0) <='0';
          end if;
        if(cVar1S0S94P013P032P033P007(0)='1' AND  D(14)='0' AND E(10)='1' )then
          cVar2S0S94P043P061nsss(0) <='1';
          else
          cVar2S0S94P043P061nsss(0) <='0';
          end if;
        if(cVar1S1S94P013P032P033P007(0)='1' AND  D(14)='0' AND E(10)='0' AND A(14)='0' )then
          cVar2S1S94P043N061P010nsss(0) <='1';
          else
          cVar2S1S94P043N061P010nsss(0) <='0';
          end if;
        if(cVar1S2S94P013P032P033P007(0)='1' AND  A( 2)='0' AND E( 0)='1' )then
          cVar2S2S94P015P068nsss(0) <='1';
          else
          cVar2S2S94P015P068nsss(0) <='0';
          end if;
        if(cVar1S3S94P013P032P033P007(0)='1' AND  A( 2)='0' AND E( 0)='0' AND A( 1)='1' )then
          cVar2S3S94P015N068P017nsss(0) <='1';
          else
          cVar2S3S94P015N068P017nsss(0) <='0';
          end if;
        if(cVar1S4S94P013P032N033P031(0)='1' AND  E( 9)='0' AND B(12)='0' )then
          cVar2S4S94P065P030nsss(0) <='1';
          else
          cVar2S4S94P065P030nsss(0) <='0';
          end if;
        if(cVar1S5S94P013P032N033P031(0)='1' AND  E( 9)='1' AND A(13)='1' )then
          cVar2S5S94P065P012nsss(0) <='1';
          else
          cVar2S5S94P065P012nsss(0) <='0';
          end if;
        if(cVar1S6S94P013P032N033N031(0)='1' AND  B( 0)='1' AND E(11)='1' AND A( 0)='0' )then
          cVar2S6S94P037P057P019nsss(0) <='1';
          else
          cVar2S6S94P037P057P019nsss(0) <='0';
          end if;
        if(cVar1S7S94P013P032N033N031(0)='1' AND  B( 0)='1' AND E(11)='0' AND D( 0)='1' )then
          cVar2S7S94P037N057P066nsss(0) <='1';
          else
          cVar2S7S94P037N057P066nsss(0) <='0';
          end if;
        if(cVar1S8S94P013P032N033N031(0)='1' AND  B( 0)='0' AND E(12)='1' )then
          cVar2S8S94N037P053nsss(0) <='1';
          else
          cVar2S8S94N037P053nsss(0) <='0';
          end if;
        if(cVar1S9S94P013P032P061P067(0)='1' AND  D( 0)='1' )then
          cVar2S9S94P066nsss(0) <='1';
          else
          cVar2S9S94P066nsss(0) <='0';
          end if;
        if(cVar1S10S94P013P032P061P067(0)='1' AND  D( 0)='0' AND B( 9)='0' )then
          cVar2S10S94N066P036nsss(0) <='1';
          else
          cVar2S10S94N066P036nsss(0) <='0';
          end if;
        if(cVar1S11S94P013P032P061N067(0)='1' AND  A( 2)='0' AND A(12)='0' AND A(10)='0' )then
          cVar2S11S94P015P014P018nsss(0) <='1';
          else
          cVar2S11S94P015P014P018nsss(0) <='0';
          end if;
        if(cVar1S12S94P013P032P061N067(0)='1' AND  A( 2)='0' AND A(12)='1' AND A(10)='1' )then
          cVar2S12S94P015P014P018nsss(0) <='1';
          else
          cVar2S12S94P015P014P018nsss(0) <='0';
          end if;
        if(cVar1S13S94P013P032P061N067(0)='1' AND  A( 2)='1' AND A( 4)='1' )then
          cVar2S13S94P015P011nsss(0) <='1';
          else
          cVar2S13S94P015P011nsss(0) <='0';
          end if;
        if(cVar1S14S94P013P032N061P063(0)='1' AND  A(12)='0' )then
          cVar2S14S94P014nsss(0) <='1';
          else
          cVar2S14S94P014nsss(0) <='0';
          end if;
        if(cVar1S15S94P013P032N061N063(0)='1' AND  A(12)='1' AND D( 2)='1' )then
          cVar2S15S94P014P058nsss(0) <='1';
          else
          cVar2S15S94P014P058nsss(0) <='0';
          end if;
        if(cVar1S16S94P013P032N061N063(0)='1' AND  A(12)='0' AND D( 8)='1' AND B( 9)='0' )then
          cVar2S16S94N014P067P036nsss(0) <='1';
          else
          cVar2S16S94N014P067P036nsss(0) <='0';
          end if;
        if(cVar1S17S94N013P017P068P018(0)='1' AND  A(15)='1' AND D( 0)='0' )then
          cVar2S17S94P008P066nsss(0) <='1';
          else
          cVar2S17S94P008P066nsss(0) <='0';
          end if;
        if(cVar1S18S94N013P017P068P018(0)='1' AND  A(15)='0' AND E( 5)='0' AND B(14)='0' )then
          cVar2S18S94N008P048P026nsss(0) <='1';
          else
          cVar2S18S94N008P048P026nsss(0) <='0';
          end if;
        if(cVar1S19S94N013P017P068P018(0)='1' AND  A(15)='0' AND E( 5)='1' AND D( 4)='1' )then
          cVar2S19S94N008P048P050nsss(0) <='1';
          else
          cVar2S19S94N008P048P050nsss(0) <='0';
          end if;
        if(cVar1S20S94N013P017P068N018(0)='1' AND  D( 2)='0' AND D( 0)='1' )then
          cVar2S20S94P058P066nsss(0) <='1';
          else
          cVar2S20S94P058P066nsss(0) <='0';
          end if;
        if(cVar1S21S94N013P017P068N018(0)='1' AND  D( 2)='0' AND D( 0)='0' AND B( 0)='0' )then
          cVar2S21S94P058N066P037nsss(0) <='1';
          else
          cVar2S21S94P058N066P037nsss(0) <='0';
          end if;
        if(cVar1S22S94N013P017P068N018(0)='1' AND  D( 2)='1' AND E(10)='0' AND E( 2)='1' )then
          cVar2S22S94P058P061P060nsss(0) <='1';
          else
          cVar2S22S94P058P061P060nsss(0) <='0';
          end if;
        if(cVar1S23S94N013P017P068P003(0)='1' AND  E( 8)='1' )then
          cVar2S23S94P069nsss(0) <='1';
          else
          cVar2S23S94P069nsss(0) <='0';
          end if;
        if(cVar1S24S94N013P017P068P003(0)='1' AND  E( 8)='0' AND A(10)='0' )then
          cVar2S24S94N069P018nsss(0) <='1';
          else
          cVar2S24S94N069P018nsss(0) <='0';
          end if;
        if(cVar1S25S94N013P017P068P003(0)='1' AND  E( 8)='0' AND A(10)='1' AND A( 4)='1' )then
          cVar2S25S94N069P018P011nsss(0) <='1';
          else
          cVar2S25S94N069P018P011nsss(0) <='0';
          end if;
        if(cVar1S26S94N013P017P068N003(0)='1' AND  B(16)='0' AND A(11)='0' AND D( 6)='0' )then
          cVar2S26S94P022P016P042nsss(0) <='1';
          else
          cVar2S26S94P022P016P042nsss(0) <='0';
          end if;
        if(cVar1S27S94N013N017P015P036(0)='1' AND  B( 3)='0' )then
          cVar2S27S94P031nsss(0) <='1';
          else
          cVar2S27S94P031nsss(0) <='0';
          end if;
        if(cVar1S28S94N013N017P015P036(0)='1' AND  B( 3)='1' AND D( 3)='1' AND A(10)='1' )then
          cVar2S28S94P031P054P018nsss(0) <='1';
          else
          cVar2S28S94P031P054P018nsss(0) <='0';
          end if;
        if(cVar1S29S94N013N017P015P036(0)='1' AND  B( 3)='1' AND D( 3)='0' AND D( 2)='1' )then
          cVar2S29S94P031N054P058nsss(0) <='1';
          else
          cVar2S29S94P031N054P058nsss(0) <='0';
          end if;
        if(cVar1S30S94N013N017P015P036(0)='1' AND  B(10)='1' AND D( 2)='0' )then
          cVar2S30S94P034P058nsss(0) <='1';
          else
          cVar2S30S94P034P058nsss(0) <='0';
          end if;
        if(cVar1S31S94N013N017P015P036(0)='1' AND  B(10)='0' AND A(17)='1' AND E( 8)='1' )then
          cVar2S31S94N034P004P069nsss(0) <='1';
          else
          cVar2S31S94N034P004P069nsss(0) <='0';
          end if;
        if(cVar1S32S94N013N017P015P036(0)='1' AND  B(10)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S32S94N034N004P005nsss(0) <='1';
          else
          cVar2S32S94N034N004P005nsss(0) <='0';
          end if;
        if(cVar1S33S94N013N017N015P019(0)='1' AND  E(10)='0' AND A(19)='1' )then
          cVar2S33S94P061P000nsss(0) <='1';
          else
          cVar2S33S94P061P000nsss(0) <='0';
          end if;
        if(cVar1S34S94N013N017N015P019(0)='1' AND  E(10)='0' AND A(19)='0' AND D(14)='0' )then
          cVar2S34S94P061N000P043nsss(0) <='1';
          else
          cVar2S34S94P061N000P043nsss(0) <='0';
          end if;
        if(cVar1S35S94N013N017N015P019(0)='1' AND  E(10)='1' AND D( 8)='1' AND E( 2)='0' )then
          cVar2S35S94P061P067P060nsss(0) <='1';
          else
          cVar2S35S94P061P067P060nsss(0) <='0';
          end if;
        if(cVar1S36S94N013N017N015N019(0)='1' AND  A(19)='0' AND B( 0)='0' AND A( 4)='1' )then
          cVar2S36S94P000P037P011nsss(0) <='1';
          else
          cVar2S36S94P000P037P011nsss(0) <='0';
          end if;
        if(cVar1S37S94N013N017N015N019(0)='1' AND  A(19)='1' AND B( 2)='0' AND D(15)='1' )then
          cVar2S37S94P000P033P039nsss(0) <='1';
          else
          cVar2S37S94P000P033P039nsss(0) <='0';
          end if;
        if(cVar1S0S95P013P032P011P003(0)='1' AND  B( 6)='1' AND D( 5)='1' )then
          cVar2S0S95P025P046nsss(0) <='1';
          else
          cVar2S0S95P025P046nsss(0) <='0';
          end if;
        if(cVar1S1S95P013P032P011P003(0)='1' AND  B( 6)='1' AND D( 5)='0' AND D( 0)='1' )then
          cVar2S1S95P025N046P066nsss(0) <='1';
          else
          cVar2S1S95P025N046P066nsss(0) <='0';
          end if;
        if(cVar1S2S95P013P032P011P003(0)='1' AND  B( 6)='0' AND D(12)='1' AND E(12)='1' )then
          cVar2S2S95N025P051P053nsss(0) <='1';
          else
          cVar2S2S95N025P051P053nsss(0) <='0';
          end if;
        if(cVar1S3S95P013P032P011P003(0)='1' AND  B( 6)='0' AND D(12)='0' AND B(13)='0' )then
          cVar2S3S95N025N051P028nsss(0) <='1';
          else
          cVar2S3S95N025N051P028nsss(0) <='0';
          end if;
        if(cVar1S4S95P013P032P011P003(0)='1' AND  E(11)='1' )then
          cVar2S4S95P057nsss(0) <='1';
          else
          cVar2S4S95P057nsss(0) <='0';
          end if;
        if(cVar1S5S95P013P032P011P003(0)='1' AND  E(11)='0' AND A( 0)='1' AND E(10)='0' )then
          cVar2S5S95N057P019P061nsss(0) <='1';
          else
          cVar2S5S95N057P019P061nsss(0) <='0';
          end if;
        if(cVar1S6S95P013P032P011P036(0)='1' AND  A(18)='1' )then
          cVar2S6S95P002nsss(0) <='1';
          else
          cVar2S6S95P002nsss(0) <='0';
          end if;
        if(cVar1S7S95P013P032P011P036(0)='1' AND  A(18)='0' AND B( 2)='1' AND A( 2)='0' )then
          cVar2S7S95N002P033P015nsss(0) <='1';
          else
          cVar2S7S95N002P033P015nsss(0) <='0';
          end if;
        if(cVar1S8S95P013P032P011P036(0)='1' AND  A(18)='0' AND B( 2)='0' AND A( 5)='0' )then
          cVar2S8S95N002N033P009nsss(0) <='1';
          else
          cVar2S8S95N002N033P009nsss(0) <='0';
          end if;
        if(cVar1S9S95P013P032P011N036(0)='1' AND  A(19)='1' AND B( 0)='1' AND A( 0)='1' )then
          cVar2S9S95P000P037P019nsss(0) <='1';
          else
          cVar2S9S95P000P037P019nsss(0) <='0';
          end if;
        if(cVar1S10S95P013P032P011N036(0)='1' AND  A(19)='1' AND B( 0)='0' AND A(11)='0' )then
          cVar2S10S95P000N037P016nsss(0) <='1';
          else
          cVar2S10S95P000N037P016nsss(0) <='0';
          end if;
        if(cVar1S11S95P013P032P011N036(0)='1' AND  A(19)='0' AND E( 4)='1' AND B( 4)='1' )then
          cVar2S11S95N000P052P029nsss(0) <='1';
          else
          cVar2S11S95N000P052P029nsss(0) <='0';
          end if;
        if(cVar1S12S95P013P032P011N036(0)='1' AND  A(19)='0' AND E( 4)='0' AND E(14)='1' )then
          cVar2S12S95N000N052P045nsss(0) <='1';
          else
          cVar2S12S95N000N052P045nsss(0) <='0';
          end if;
        if(cVar1S14S95P013P032P061N067(0)='1' AND  A( 2)='0' AND B( 2)='1' )then
          cVar2S14S95P015P033nsss(0) <='1';
          else
          cVar2S14S95P015P033nsss(0) <='0';
          end if;
        if(cVar1S15S95P013P032P061N067(0)='1' AND  A( 2)='0' AND B( 2)='0' AND A(12)='0' )then
          cVar2S15S95P015N033P014nsss(0) <='1';
          else
          cVar2S15S95P015N033P014nsss(0) <='0';
          end if;
        if(cVar1S16S95P013P032P061N067(0)='1' AND  A( 2)='1' AND A( 4)='1' )then
          cVar2S16S95P015P011nsss(0) <='1';
          else
          cVar2S16S95P015P011nsss(0) <='0';
          end if;
        if(cVar1S17S95P013P032P061N067(0)='1' AND  A( 2)='1' AND A( 4)='0' AND B( 0)='1' )then
          cVar2S17S95P015N011P037nsss(0) <='1';
          else
          cVar2S17S95P015N011P037nsss(0) <='0';
          end if;
        if(cVar1S18S95P013P032N061P063(0)='1' AND  A( 2)='0' )then
          cVar2S18S95P015nsss(0) <='1';
          else
          cVar2S18S95P015nsss(0) <='0';
          end if;
        if(cVar1S19S95P013P032N061N063(0)='1' AND  A(12)='1' AND D( 2)='1' )then
          cVar2S19S95P014P058nsss(0) <='1';
          else
          cVar2S19S95P014P058nsss(0) <='0';
          end if;
        if(cVar1S20S95P013P032N061N063(0)='1' AND  A(12)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar2S20S95P014N058P011nsss(0) <='1';
          else
          cVar2S20S95P014N058P011nsss(0) <='0';
          end if;
        if(cVar1S21S95N013P019P041P004(0)='1' AND  B(16)='1' )then
          cVar2S21S95P022nsss(0) <='1';
          else
          cVar2S21S95P022nsss(0) <='0';
          end if;
        if(cVar1S22S95N013P019P041P004(0)='1' AND  B(16)='0' AND B(17)='1' )then
          cVar2S22S95N022P020nsss(0) <='1';
          else
          cVar2S22S95N022P020nsss(0) <='0';
          end if;
        if(cVar1S23S95N013P019P041N004(0)='1' AND  D( 0)='0' AND E( 7)='0' AND D( 9)='0' )then
          cVar2S23S95P066P040P063nsss(0) <='1';
          else
          cVar2S23S95P066P040P063nsss(0) <='0';
          end if;
        if(cVar1S24S95N013P019P041N004(0)='1' AND  D( 0)='0' AND E( 7)='1' AND D(15)='0' )then
          cVar2S24S95P066P040P039nsss(0) <='1';
          else
          cVar2S24S95P066P040P039nsss(0) <='0';
          end if;
        if(cVar1S25S95N013P019P041N004(0)='1' AND  D( 0)='1' AND A(12)='0' AND E( 0)='1' )then
          cVar2S25S95P066P014P068nsss(0) <='1';
          else
          cVar2S25S95P066P014P068nsss(0) <='0';
          end if;
        if(cVar1S26S95N013P019N041P020(0)='1' AND  A(13)='1' AND A(14)='0' )then
          cVar2S26S95P012P010nsss(0) <='1';
          else
          cVar2S26S95P012P010nsss(0) <='0';
          end if;
        if(cVar1S27S95N013P019N041P020(0)='1' AND  A(13)='0' AND B( 7)='1' AND B(14)='0' )then
          cVar2S27S95N012P023P026nsss(0) <='1';
          else
          cVar2S27S95N012P023P026nsss(0) <='0';
          end if;
        if(cVar1S28S95N013P019N041P020(0)='1' AND  B( 2)='0' AND B(14)='1' )then
          cVar2S28S95P033P026nsss(0) <='1';
          else
          cVar2S28S95P033P026nsss(0) <='0';
          end if;
        if(cVar1S29S95N013P019N041P020(0)='1' AND  B( 2)='0' AND B(14)='0' AND B(11)='1' )then
          cVar2S29S95P033N026P032nsss(0) <='1';
          else
          cVar2S29S95P033N026P032nsss(0) <='0';
          end if;
        if(cVar1S30S95N013P019P017P066(0)='1' AND  B( 5)='1' AND A(10)='0' )then
          cVar2S30S95P027P018nsss(0) <='1';
          else
          cVar2S30S95P027P018nsss(0) <='0';
          end if;
        if(cVar1S31S95N013P019P017P066(0)='1' AND  B( 5)='1' AND A(10)='1' AND A(12)='0' )then
          cVar2S31S95P027P018P014nsss(0) <='1';
          else
          cVar2S31S95P027P018P014nsss(0) <='0';
          end if;
        if(cVar1S32S95N013P019P017P066(0)='1' AND  B( 5)='0' AND A(18)='0' )then
          cVar2S32S95N027P002nsss(0) <='1';
          else
          cVar2S32S95N027P002nsss(0) <='0';
          end if;
        if(cVar1S33S95N013P019P017P066(0)='1' AND  B( 5)='0' AND A(18)='1' AND A( 5)='1' )then
          cVar2S33S95N027P002P009nsss(0) <='1';
          else
          cVar2S33S95N027P002P009nsss(0) <='0';
          end if;
        if(cVar1S34S95N013P019P017P066(0)='1' AND  A(19)='0' AND D( 9)='1' )then
          cVar2S34S95P000P063nsss(0) <='1';
          else
          cVar2S34S95P000P063nsss(0) <='0';
          end if;
        if(cVar1S35S95N013P019N017P048(0)='1' AND  E(13)='1' )then
          cVar2S35S95P049nsss(0) <='1';
          else
          cVar2S35S95P049nsss(0) <='0';
          end if;
        if(cVar1S36S95N013P019N017P048(0)='1' AND  E(13)='0' AND A(14)='1' )then
          cVar2S36S95N049P010nsss(0) <='1';
          else
          cVar2S36S95N049P010nsss(0) <='0';
          end if;
        if(cVar1S37S95N013P019N017P048(0)='1' AND  E(13)='0' AND A(14)='0' AND A( 5)='1' )then
          cVar2S37S95N049N010P009nsss(0) <='1';
          else
          cVar2S37S95N049N010P009nsss(0) <='0';
          end if;
        if(cVar1S38S95N013P019N017N048(0)='1' AND  A( 9)='1' AND A(11)='0' )then
          cVar2S38S95P001P016nsss(0) <='1';
          else
          cVar2S38S95P001P016nsss(0) <='0';
          end if;
        if(cVar1S39S95N013P019N017N048(0)='1' AND  A( 9)='1' AND A(11)='1' AND B( 9)='0' )then
          cVar2S39S95P001P016P036nsss(0) <='1';
          else
          cVar2S39S95P001P016P036nsss(0) <='0';
          end if;
        if(cVar1S40S95N013P019N017N048(0)='1' AND  A( 9)='0' AND B(13)='1' AND D(11)='1' )then
          cVar2S40S95N001P028P055nsss(0) <='1';
          else
          cVar2S40S95N001P028P055nsss(0) <='0';
          end if;
        if(cVar1S0S96P019P012P058P011(0)='1' AND  A(12)='1' )then
          cVar2S0S96P014nsss(0) <='1';
          else
          cVar2S0S96P014nsss(0) <='0';
          end if;
        if(cVar1S1S96P019P012P058P011(0)='1' AND  A(12)='0' AND E( 2)='0' AND E( 3)='0' )then
          cVar2S1S96N014P060P056nsss(0) <='1';
          else
          cVar2S1S96N014P060P056nsss(0) <='0';
          end if;
        if(cVar1S2S96P019P012P058P011(0)='1' AND  A(12)='0' AND E( 2)='1' AND E( 0)='1' )then
          cVar2S2S96N014P060P068nsss(0) <='1';
          else
          cVar2S2S96N014P060P068nsss(0) <='0';
          end if;
        if(cVar1S3S96P019P012P058P011(0)='1' AND  B(16)='1' AND A( 2)='1' )then
          cVar2S3S96P022P015nsss(0) <='1';
          else
          cVar2S3S96P022P015nsss(0) <='0';
          end if;
        if(cVar1S4S96P019P012P058P011(0)='1' AND  B(16)='1' AND A( 2)='0' AND A(11)='0' )then
          cVar2S4S96P022N015P016nsss(0) <='1';
          else
          cVar2S4S96P022N015P016nsss(0) <='0';
          end if;
        if(cVar1S5S96P019P012P058P011(0)='1' AND  B(16)='0' AND E(13)='1' AND A( 2)='0' )then
          cVar2S5S96N022P049P015nsss(0) <='1';
          else
          cVar2S5S96N022P049P015nsss(0) <='0';
          end if;
        if(cVar1S6S96P019P012P058P011(0)='1' AND  B(16)='0' AND E(13)='0' AND B( 4)='1' )then
          cVar2S6S96N022N049P029nsss(0) <='1';
          else
          cVar2S6S96N022N049P029nsss(0) <='0';
          end if;
        if(cVar1S7S96P019P012P058P068(0)='1' AND  A(10)='1' AND E(10)='1' )then
          cVar2S7S96P018P061nsss(0) <='1';
          else
          cVar2S7S96P018P061nsss(0) <='0';
          end if;
        if(cVar1S8S96P019P012P058P068(0)='1' AND  A(10)='1' AND E(10)='0' AND A(12)='1' )then
          cVar2S8S96P018N061P014nsss(0) <='1';
          else
          cVar2S8S96P018N061P014nsss(0) <='0';
          end if;
        if(cVar1S9S96P019P012P058P068(0)='1' AND  A(10)='0' AND B(12)='1' )then
          cVar2S9S96N018P030nsss(0) <='1';
          else
          cVar2S9S96N018P030nsss(0) <='0';
          end if;
        if(cVar1S10S96P019P012P058P068(0)='1' AND  A(10)='0' AND B(12)='0' AND B( 2)='0' )then
          cVar2S10S96N018N030P033nsss(0) <='1';
          else
          cVar2S10S96N018N030P033nsss(0) <='0';
          end if;
        if(cVar1S11S96P019P012P058P068(0)='1' AND  B( 1)='0' AND A(17)='1' )then
          cVar2S11S96P035P004nsss(0) <='1';
          else
          cVar2S11S96P035P004nsss(0) <='0';
          end if;
        if(cVar1S12S96P019P012P058P068(0)='1' AND  B( 1)='1' AND A( 1)='1' AND E( 1)='0' )then
          cVar2S12S96P035P017P064nsss(0) <='1';
          else
          cVar2S12S96P035P017P064nsss(0) <='0';
          end if;
        if(cVar1S13S96P019P012P043P056(0)='1' AND  D( 1)='0' AND A( 1)='1' )then
          cVar2S13S96P062P017nsss(0) <='1';
          else
          cVar2S13S96P062P017nsss(0) <='0';
          end if;
        if(cVar1S14S96P019P012P043P056(0)='1' AND  D( 1)='0' AND A( 1)='0' AND A(12)='1' )then
          cVar2S14S96P062N017P014nsss(0) <='1';
          else
          cVar2S14S96P062N017P014nsss(0) <='0';
          end if;
        if(cVar1S15S96P019P012P043P056(0)='1' AND  D( 1)='1' AND D( 9)='0' AND A(12)='0' )then
          cVar2S15S96P062P063P014nsss(0) <='1';
          else
          cVar2S15S96P062P063P014nsss(0) <='0';
          end if;
        if(cVar1S16S96P019P012P043N056(0)='1' AND  A( 6)='0' AND B( 3)='1' AND E( 2)='1' )then
          cVar2S16S96P007P031P060nsss(0) <='1';
          else
          cVar2S16S96P007P031P060nsss(0) <='0';
          end if;
        if(cVar1S17S96P019P012P043N056(0)='1' AND  A( 6)='1' AND D(13)='1' )then
          cVar2S17S96P007P047nsss(0) <='1';
          else
          cVar2S17S96P007P047nsss(0) <='0';
          end if;
        if(cVar1S18S96P019P012P043N056(0)='1' AND  A( 6)='1' AND D(13)='0' AND D( 4)='1' )then
          cVar2S18S96P007N047P050nsss(0) <='1';
          else
          cVar2S18S96P007N047P050nsss(0) <='0';
          end if;
        if(cVar1S20S96P019P003P057P015(0)='1' AND  A(10)='0' )then
          cVar2S20S96P018nsss(0) <='1';
          else
          cVar2S20S96P018nsss(0) <='0';
          end if;
        if(cVar1S21S96P019P003N057P068(0)='1' AND  D(10)='1' )then
          cVar2S21S96P059nsss(0) <='1';
          else
          cVar2S21S96P059nsss(0) <='0';
          end if;
        if(cVar1S22S96P019P003N057P068(0)='1' AND  D(10)='0' AND B(11)='0' )then
          cVar2S22S96N059P032nsss(0) <='1';
          else
          cVar2S22S96N059P032nsss(0) <='0';
          end if;
        if(cVar1S23S96P019P003N057N068(0)='1' AND  D( 8)='1' AND A(12)='1' AND E( 8)='1' )then
          cVar2S23S96P067P014P069nsss(0) <='1';
          else
          cVar2S23S96P067P014P069nsss(0) <='0';
          end if;
        if(cVar1S24S96P019P003N057N068(0)='1' AND  D( 8)='1' AND A(12)='0' AND A( 1)='0' )then
          cVar2S24S96P067N014P017nsss(0) <='1';
          else
          cVar2S24S96P067N014P017nsss(0) <='0';
          end if;
        if(cVar1S25S96P019P003N057N068(0)='1' AND  D( 8)='0' AND A( 5)='1' AND A( 1)='1' )then
          cVar2S25S96N067P009P017nsss(0) <='1';
          else
          cVar2S25S96N067P009P017nsss(0) <='0';
          end if;
        if(cVar1S26S96P019N003P057P025(0)='1' AND  D( 4)='0' AND A( 3)='1' AND A(12)='0' )then
          cVar2S26S96P050P013P014nsss(0) <='1';
          else
          cVar2S26S96P050P013P014nsss(0) <='0';
          end if;
        if(cVar1S27S96P019N003P057P025(0)='1' AND  D( 4)='0' AND A( 3)='0' AND A(14)='0' )then
          cVar2S27S96P050N013P010nsss(0) <='1';
          else
          cVar2S27S96P050N013P010nsss(0) <='0';
          end if;
        if(cVar1S28S96P019N003P057N025(0)='1' AND  A(14)='1' AND E( 5)='1' AND A(10)='0' )then
          cVar2S28S96P010P048P018nsss(0) <='1';
          else
          cVar2S28S96P010P048P018nsss(0) <='0';
          end if;
        if(cVar1S29S96P019N003P057N025(0)='1' AND  A(14)='1' AND E( 5)='0' AND D( 0)='1' )then
          cVar2S29S96P010N048P066nsss(0) <='1';
          else
          cVar2S29S96P010N048P066nsss(0) <='0';
          end if;
        if(cVar1S30S96P019N003P057N025(0)='1' AND  A(14)='0' AND D(13)='0' AND A(18)='1' )then
          cVar2S30S96N010P047P002nsss(0) <='1';
          else
          cVar2S30S96N010P047P002nsss(0) <='0';
          end if;
        if(cVar1S31S96P019N003P057N025(0)='1' AND  A(14)='0' AND D(13)='1' AND B(15)='1' )then
          cVar2S31S96N010P047P024nsss(0) <='1';
          else
          cVar2S31S96N010P047P024nsss(0) <='0';
          end if;
        if(cVar1S32S96P019N003P057P066(0)='1' AND  B( 9)='0' AND D( 3)='0' AND A( 6)='0' )then
          cVar2S32S96P036P054P007nsss(0) <='1';
          else
          cVar2S32S96P036P054P007nsss(0) <='0';
          end if;
        if(cVar1S33S96P019N003P057P066(0)='1' AND  B( 9)='0' AND D( 3)='1' AND A( 1)='1' )then
          cVar2S33S96P036P054P017nsss(0) <='1';
          else
          cVar2S33S96P036P054P017nsss(0) <='0';
          end if;
        if(cVar1S34S96P019N003P057P066(0)='1' AND  B( 9)='1' AND A( 4)='1' )then
          cVar2S34S96P036P011nsss(0) <='1';
          else
          cVar2S34S96P036P011nsss(0) <='0';
          end if;
        if(cVar1S35S96P019N003P057P066(0)='1' AND  E( 9)='1' )then
          cVar2S35S96P065nsss(0) <='1';
          else
          cVar2S35S96P065nsss(0) <='0';
          end if;
        if(cVar1S36S96P019N003P057P066(0)='1' AND  E( 9)='0' AND B(12)='1' AND A( 2)='1' )then
          cVar2S36S96N065P030P015nsss(0) <='1';
          else
          cVar2S36S96N065P030P015nsss(0) <='0';
          end if;
        if(cVar1S0S97P019P057P069P007(0)='1' AND  A(15)='0' )then
          cVar2S0S97P008nsss(0) <='1';
          else
          cVar2S0S97P008nsss(0) <='0';
          end if;
        if(cVar1S1S97P019P057P069P007(0)='1' AND  A(15)='1' AND A( 4)='0' )then
          cVar2S1S97P008P011nsss(0) <='1';
          else
          cVar2S1S97P008P011nsss(0) <='0';
          end if;
        if(cVar1S2S97P019P057P069N007(0)='1' AND  A( 3)='1' AND B( 1)='0' )then
          cVar2S2S97P013P035nsss(0) <='1';
          else
          cVar2S2S97P013P035nsss(0) <='0';
          end if;
        if(cVar1S3S97P019P057P069N007(0)='1' AND  A( 3)='1' AND B( 1)='1' AND A(12)='1' )then
          cVar2S3S97P013P035P014nsss(0) <='1';
          else
          cVar2S3S97P013P035P014nsss(0) <='0';
          end if;
        if(cVar1S4S97P019P057P069N007(0)='1' AND  A( 3)='0' )then
          cVar2S4S97N013psss(0) <='1';
          else
          cVar2S4S97N013psss(0) <='0';
          end if;
        if(cVar1S5S97P019P057N069P038(0)='1' AND  D(11)='0' AND D( 2)='1' AND B(17)='0' )then
          cVar2S5S97P055P058P020nsss(0) <='1';
          else
          cVar2S5S97P055P058P020nsss(0) <='0';
          end if;
        if(cVar1S6S97P019P057N069P038(0)='1' AND  D(11)='0' AND D( 2)='0' )then
          cVar2S6S97P055N058psss(0) <='1';
          else
          cVar2S6S97P055N058psss(0) <='0';
          end if;
        if(cVar1S7S97P019P057N069P038(0)='1' AND  D(11)='1' AND D( 9)='1' )then
          cVar2S7S97P055P063nsss(0) <='1';
          else
          cVar2S7S97P055P063nsss(0) <='0';
          end if;
        if(cVar1S8S97P019P057N069P038(0)='1' AND  B( 8)='1' )then
          cVar2S8S97P021nsss(0) <='1';
          else
          cVar2S8S97P021nsss(0) <='0';
          end if;
        if(cVar1S10S97P019P057P003P015(0)='1' AND  A( 3)='0' )then
          cVar2S10S97P013nsss(0) <='1';
          else
          cVar2S10S97P013nsss(0) <='0';
          end if;
        if(cVar1S11S97P019P057N003P011(0)='1' AND  A( 3)='0' AND D(11)='1' )then
          cVar2S11S97P013P055nsss(0) <='1';
          else
          cVar2S11S97P013P055nsss(0) <='0';
          end if;
        if(cVar1S12S97P019P057N003P011(0)='1' AND  A( 3)='1' AND D( 1)='1' )then
          cVar2S12S97P013P062nsss(0) <='1';
          else
          cVar2S12S97P013P062nsss(0) <='0';
          end if;
        if(cVar1S13S97P019P057N003N011(0)='1' AND  D( 0)='0' AND B( 9)='0' )then
          cVar2S13S97P066P036nsss(0) <='1';
          else
          cVar2S13S97P066P036nsss(0) <='0';
          end if;
        if(cVar1S14S97P019P057N003N011(0)='1' AND  D( 0)='1' AND A( 3)='1' AND A(12)='1' )then
          cVar2S14S97P066P013P014nsss(0) <='1';
          else
          cVar2S14S97P066P013P014nsss(0) <='0';
          end if;
        if(cVar1S15S97P019P057N003N011(0)='1' AND  D( 0)='1' AND A( 3)='0' AND D( 9)='1' )then
          cVar2S15S97P066N013P063nsss(0) <='1';
          else
          cVar2S15S97P066N013P063nsss(0) <='0';
          end if;
        if(cVar1S16S97N019P060P021P055(0)='1' AND  B(13)='0' AND A(14)='1' AND B( 2)='1' )then
          cVar2S16S97P028P010P033nsss(0) <='1';
          else
          cVar2S16S97P028P010P033nsss(0) <='0';
          end if;
        if(cVar1S17S97N019P060P021P055(0)='1' AND  B(13)='0' AND A(14)='0' )then
          cVar2S17S97P028N010psss(0) <='1';
          else
          cVar2S17S97P028N010psss(0) <='0';
          end if;
        if(cVar1S18S97N019P060P021P055(0)='1' AND  B(13)='1' AND D( 1)='1' )then
          cVar2S18S97P028P062nsss(0) <='1';
          else
          cVar2S18S97P028P062nsss(0) <='0';
          end if;
        if(cVar1S19S97N019P060P021P055(0)='1' AND  E( 1)='0' AND B( 2)='0' AND B( 1)='0' )then
          cVar2S19S97P064P033P035nsss(0) <='1';
          else
          cVar2S19S97P064P033P035nsss(0) <='0';
          end if;
        if(cVar1S20S97N019P060P021P055(0)='1' AND  E( 1)='0' AND B( 2)='1' AND A(13)='0' )then
          cVar2S20S97P064P033P012nsss(0) <='1';
          else
          cVar2S20S97P064P033P012nsss(0) <='0';
          end if;
        if(cVar1S22S97N019N060P068P036(0)='1' AND  D( 7)='0' AND E( 1)='1' )then
          cVar2S22S97P038P064nsss(0) <='1';
          else
          cVar2S22S97P038P064nsss(0) <='0';
          end if;
        if(cVar1S23S97N019N060P068P036(0)='1' AND  D( 7)='0' AND E( 1)='0' AND A(10)='1' )then
          cVar2S23S97P038N064P018nsss(0) <='1';
          else
          cVar2S23S97P038N064P018nsss(0) <='0';
          end if;
        if(cVar1S24S97N019N060P068N036(0)='1' AND  E( 3)='1' AND E( 9)='0' AND A( 9)='0' )then
          cVar2S24S97P056P065P001nsss(0) <='1';
          else
          cVar2S24S97P056P065P001nsss(0) <='0';
          end if;
        if(cVar1S25S97N019N060P068N036(0)='1' AND  E( 3)='1' AND E( 9)='1' AND B( 4)='1' )then
          cVar2S25S97P056P065P029nsss(0) <='1';
          else
          cVar2S25S97P056P065P029nsss(0) <='0';
          end if;
        if(cVar1S26S97N019N060P068N036(0)='1' AND  E( 3)='0' AND B( 8)='1' )then
          cVar2S26S97N056P021nsss(0) <='1';
          else
          cVar2S26S97N056P021nsss(0) <='0';
          end if;
        if(cVar1S27S97N019N060P068P023(0)='1' AND  A( 1)='0' AND E( 1)='0' AND B(10)='1' )then
          cVar2S27S97P017P064P034nsss(0) <='1';
          else
          cVar2S27S97P017P064P034nsss(0) <='0';
          end if;
        if(cVar1S28S97N019N060P068P023(0)='1' AND  A( 1)='0' AND E( 1)='1' AND A( 2)='1' )then
          cVar2S28S97P017P064P015nsss(0) <='1';
          else
          cVar2S28S97P017P064P015nsss(0) <='0';
          end if;
        if(cVar1S29S97N019N060P068P023(0)='1' AND  A( 1)='1' AND E(11)='1' )then
          cVar2S29S97P017P057nsss(0) <='1';
          else
          cVar2S29S97P017P057nsss(0) <='0';
          end if;
        if(cVar1S30S97N019N060P068P023(0)='1' AND  A( 1)='1' AND E(11)='0' AND B( 1)='1' )then
          cVar2S30S97P017N057P035nsss(0) <='1';
          else
          cVar2S30S97P017N057P035nsss(0) <='0';
          end if;
        if(cVar1S31S97N019N060P068P023(0)='1' AND  B( 0)='1' AND A(10)='1' )then
          cVar2S31S97P037P018nsss(0) <='1';
          else
          cVar2S31S97P037P018nsss(0) <='0';
          end if;
        if(cVar1S0S98P019P060P033P003(0)='1' AND  A(10)='1' AND E( 9)='1' )then
          cVar2S0S98P018P065nsss(0) <='1';
          else
          cVar2S0S98P018P065nsss(0) <='0';
          end if;
        if(cVar1S1S98P019P060P033P003(0)='1' AND  A(10)='1' AND E( 9)='0' AND D( 9)='0' )then
          cVar2S1S98P018N065P063nsss(0) <='1';
          else
          cVar2S1S98P018N065P063nsss(0) <='0';
          end if;
        if(cVar1S2S98P019P060P033P003(0)='1' AND  A(10)='0' AND D(10)='1' )then
          cVar2S2S98N018P059nsss(0) <='1';
          else
          cVar2S2S98N018P059nsss(0) <='0';
          end if;
        if(cVar1S3S98P019P060P033P003(0)='1' AND  A(10)='0' AND D(10)='0' AND D(11)='1' )then
          cVar2S3S98N018N059P055nsss(0) <='1';
          else
          cVar2S3S98N018N059P055nsss(0) <='0';
          end if;
        if(cVar1S4S98P019P060P033P003(0)='1' AND  D( 0)='0' AND E( 8)='0' AND A( 2)='1' )then
          cVar2S4S98P066P069P015nsss(0) <='1';
          else
          cVar2S4S98P066P069P015nsss(0) <='0';
          end if;
        if(cVar1S5S98P019P060N033P058(0)='1' AND  D(12)='1' AND E( 5)='0' )then
          cVar2S5S98P051P048nsss(0) <='1';
          else
          cVar2S5S98P051P048nsss(0) <='0';
          end if;
        if(cVar1S6S98P019P060N033P058(0)='1' AND  D(12)='0' )then
          cVar2S6S98N051psss(0) <='1';
          else
          cVar2S6S98N051psss(0) <='0';
          end if;
        if(cVar1S7S98P019P060N033P058(0)='1' AND  B(12)='1' AND D(11)='0' )then
          cVar2S7S98P030P055nsss(0) <='1';
          else
          cVar2S7S98P030P055nsss(0) <='0';
          end if;
        if(cVar1S8S98P019P060N033P058(0)='1' AND  B(12)='0' AND B(10)='1' AND A( 1)='1' )then
          cVar2S8S98N030P034P017nsss(0) <='1';
          else
          cVar2S8S98N030P034P017nsss(0) <='0';
          end if;
        if(cVar1S9S98P019P060P021P010(0)='1' AND  A(12)='1' AND B( 0)='0' )then
          cVar2S9S98P014P037nsss(0) <='1';
          else
          cVar2S9S98P014P037nsss(0) <='0';
          end if;
        if(cVar1S10S98P019P060P021P010(0)='1' AND  A(12)='0' AND D( 3)='1' AND B( 2)='1' )then
          cVar2S10S98N014P054P033nsss(0) <='1';
          else
          cVar2S10S98N014P054P033nsss(0) <='0';
          end if;
        if(cVar1S11S98P019P060P021P010(0)='1' AND  A(12)='0' AND D( 3)='0' AND B(11)='1' )then
          cVar2S11S98N014N054P032nsss(0) <='1';
          else
          cVar2S11S98N014N054P032nsss(0) <='0';
          end if;
        if(cVar1S12S98P019P060P021N010(0)='1' AND  B( 2)='0' AND A(13)='1' )then
          cVar2S12S98P033P012nsss(0) <='1';
          else
          cVar2S12S98P033P012nsss(0) <='0';
          end if;
        if(cVar1S13S98P019P060P021N010(0)='1' AND  B( 2)='0' AND A(13)='0' AND D( 0)='1' )then
          cVar2S13S98P033N012P066nsss(0) <='1';
          else
          cVar2S13S98P033N012P066nsss(0) <='0';
          end if;
        if(cVar1S15S98P019P069P013P017(0)='1' AND  D( 2)='1' )then
          cVar2S15S98P058nsss(0) <='1';
          else
          cVar2S15S98P058nsss(0) <='0';
          end if;
        if(cVar1S16S98P019P069P013P017(0)='1' AND  D( 2)='0' AND A(16)='0' AND A(14)='0' )then
          cVar2S16S98N058P006P010nsss(0) <='1';
          else
          cVar2S16S98N058P006P010nsss(0) <='0';
          end if;
        if(cVar1S17S98P019P069P013P017(0)='1' AND  A(12)='1' AND B(10)='0' )then
          cVar2S17S98P014P034nsss(0) <='1';
          else
          cVar2S17S98P014P034nsss(0) <='0';
          end if;
        if(cVar1S18S98P019P069P013P017(0)='1' AND  A(12)='0' AND A( 8)='0' AND B( 0)='0' )then
          cVar2S18S98N014P003P037nsss(0) <='1';
          else
          cVar2S18S98N014P003P037nsss(0) <='0';
          end if;
        if(cVar1S20S98P019P069N013N022(0)='1' AND  A( 6)='1' AND E( 1)='1' )then
          cVar2S20S98P007P064nsss(0) <='1';
          else
          cVar2S20S98P007P064nsss(0) <='0';
          end if;
        if(cVar1S21S98P019P069N013N022(0)='1' AND  A( 6)='1' AND E( 1)='0' AND A( 2)='1' )then
          cVar2S21S98P007N064P015nsss(0) <='1';
          else
          cVar2S21S98P007N064P015nsss(0) <='0';
          end if;
        if(cVar1S22S98P019P069N013N022(0)='1' AND  A( 6)='0' AND D(14)='1' )then
          cVar2S22S98N007P043nsss(0) <='1';
          else
          cVar2S22S98N007P043nsss(0) <='0';
          end if;
        if(cVar1S23S98P019N069P058P063(0)='1' AND  D( 1)='1' )then
          cVar2S23S98P062nsss(0) <='1';
          else
          cVar2S23S98P062nsss(0) <='0';
          end if;
        if(cVar1S24S98P019N069P058P063(0)='1' AND  D( 1)='0' AND E(10)='0' )then
          cVar2S24S98N062P061nsss(0) <='1';
          else
          cVar2S24S98N062P061nsss(0) <='0';
          end if;
        if(cVar1S25S98P019N069P058N063(0)='1' AND  A( 6)='0' AND B( 0)='0' AND B( 2)='1' )then
          cVar2S25S98P007P037P033nsss(0) <='1';
          else
          cVar2S25S98P007P037P033nsss(0) <='0';
          end if;
        if(cVar1S26S98P019N069P058N063(0)='1' AND  A( 6)='1' AND B( 1)='1' )then
          cVar2S26S98P007P035nsss(0) <='1';
          else
          cVar2S26S98P007P035nsss(0) <='0';
          end if;
        if(cVar1S27S98P019N069N058P060(0)='1' AND  D( 3)='1' AND E(11)='0' AND A( 3)='0' )then
          cVar2S27S98P054P057P013nsss(0) <='1';
          else
          cVar2S27S98P054P057P013nsss(0) <='0';
          end if;
        if(cVar1S28S98P019N069N058P060(0)='1' AND  D( 3)='1' AND E(11)='1' AND A( 1)='1' )then
          cVar2S28S98P054P057P017nsss(0) <='1';
          else
          cVar2S28S98P054P057P017nsss(0) <='0';
          end if;
        if(cVar1S29S98P019N069N058P060(0)='1' AND  D( 3)='0' AND B( 3)='1' AND E(11)='1' )then
          cVar2S29S98N054P031P057nsss(0) <='1';
          else
          cVar2S29S98N054P031P057nsss(0) <='0';
          end if;
        if(cVar1S30S98P019N069N058P060(0)='1' AND  B(14)='0' AND D( 0)='1' AND E(10)='0' )then
          cVar2S30S98P026P066P061nsss(0) <='1';
          else
          cVar2S30S98P026P066P061nsss(0) <='0';
          end if;
        if(cVar1S1S99P019P069P006N027(0)='1' AND  E( 6)='1' )then
          cVar2S1S99P044nsss(0) <='1';
          else
          cVar2S1S99P044nsss(0) <='0';
          end if;
        if(cVar1S2S99P019P069P006N027(0)='1' AND  E( 6)='0' AND D(13)='1' )then
          cVar2S2S99N044P047nsss(0) <='1';
          else
          cVar2S2S99N044P047nsss(0) <='0';
          end if;
        if(cVar1S3S99P019P069P006N027(0)='1' AND  E( 6)='0' AND D(13)='0' AND A(15)='1' )then
          cVar2S3S99N044N047P008nsss(0) <='1';
          else
          cVar2S3S99N044N047P008nsss(0) <='0';
          end if;
        if(cVar1S4S99P019P069N006P047(0)='1' AND  B( 6)='1' AND D( 0)='1' )then
          cVar2S4S99P025P066nsss(0) <='1';
          else
          cVar2S4S99P025P066nsss(0) <='0';
          end if;
        if(cVar1S5S99P019P069N006P047(0)='1' AND  B( 6)='1' AND D( 0)='0' AND A(10)='0' )then
          cVar2S5S99P025N066P018nsss(0) <='1';
          else
          cVar2S5S99P025N066P018nsss(0) <='0';
          end if;
        if(cVar1S6S99P019P069N006P047(0)='1' AND  B( 6)='0' AND A(15)='0' )then
          cVar2S6S99N025P008nsss(0) <='1';
          else
          cVar2S6S99N025P008nsss(0) <='0';
          end if;
        if(cVar1S7S99P019P069N006P047(0)='1' AND  E(13)='1' AND B(14)='1' )then
          cVar2S7S99P049P026nsss(0) <='1';
          else
          cVar2S7S99P049P026nsss(0) <='0';
          end if;
        if(cVar1S8S99P019N069P060P016(0)='1' AND  D( 1)='1' AND E(11)='1' )then
          cVar2S8S99P062P057nsss(0) <='1';
          else
          cVar2S8S99P062P057nsss(0) <='0';
          end if;
        if(cVar1S9S99P019N069P060P016(0)='1' AND  D( 1)='1' AND E(11)='0' AND A(10)='0' )then
          cVar2S9S99P062N057P018nsss(0) <='1';
          else
          cVar2S9S99P062N057P018nsss(0) <='0';
          end if;
        if(cVar1S10S99P019N069P060P016(0)='1' AND  D( 1)='0' AND B(10)='0' AND E( 3)='0' )then
          cVar2S10S99N062P034P056nsss(0) <='1';
          else
          cVar2S10S99N062P034P056nsss(0) <='0';
          end if;
        if(cVar1S11S99P019N069P060P016(0)='1' AND  D( 1)='0' AND B(10)='1' AND B(17)='1' )then
          cVar2S11S99N062P034P020nsss(0) <='1';
          else
          cVar2S11S99N062P034P020nsss(0) <='0';
          end if;
        if(cVar1S12S99P019N069P060N016(0)='1' AND  A( 9)='1' AND A( 4)='0' AND A( 7)='0' )then
          cVar2S12S99P001P011P005nsss(0) <='1';
          else
          cVar2S12S99P001P011P005nsss(0) <='0';
          end if;
        if(cVar1S13S99P019N069P060N016(0)='1' AND  A( 9)='1' AND A( 4)='1' AND A(12)='1' )then
          cVar2S13S99P001P011P014nsss(0) <='1';
          else
          cVar2S13S99P001P011P014nsss(0) <='0';
          end if;
        if(cVar1S14S99P019N069P060N016(0)='1' AND  A( 9)='0' AND D(10)='1' )then
          cVar2S14S99N001P059nsss(0) <='1';
          else
          cVar2S14S99N001P059nsss(0) <='0';
          end if;
        if(cVar1S15S99P019N069P060N016(0)='1' AND  A( 9)='0' AND D(10)='0' AND B( 2)='0' )then
          cVar2S15S99N001N059P033nsss(0) <='1';
          else
          cVar2S15S99N001N059P033nsss(0) <='0';
          end if;
        if(cVar1S16S99P019N069P060P058(0)='1' AND  B(17)='0' AND A(18)='0' AND D( 9)='1' )then
          cVar2S16S99P020P002P063nsss(0) <='1';
          else
          cVar2S16S99P020P002P063nsss(0) <='0';
          end if;
        if(cVar1S17S99P019N069P060N058(0)='1' AND  B(14)='0' AND D( 1)='1' AND D( 0)='1' )then
          cVar2S17S99P026P062P066nsss(0) <='1';
          else
          cVar2S17S99P026P062P066nsss(0) <='0';
          end if;
        if(cVar1S18S99P019N069P060N058(0)='1' AND  B(14)='0' AND D( 1)='0' AND E( 9)='1' )then
          cVar2S18S99P026N062P065nsss(0) <='1';
          else
          cVar2S18S99P026N062P065nsss(0) <='0';
          end if;
        if(cVar1S19S99N019P033P030P003(0)='1' AND  B(17)='0' AND E( 2)='0' )then
          cVar2S19S99P020P060nsss(0) <='1';
          else
          cVar2S19S99P020P060nsss(0) <='0';
          end if;
        if(cVar1S20S99N019P033P030P003(0)='1' AND  B(17)='0' AND E( 2)='1' AND D(10)='0' )then
          cVar2S20S99P020P060P059nsss(0) <='1';
          else
          cVar2S20S99P020P060P059nsss(0) <='0';
          end if;
        if(cVar1S21S99N019P033P030P003(0)='1' AND  B(17)='1' AND B( 0)='1' )then
          cVar2S21S99P020P037nsss(0) <='1';
          else
          cVar2S21S99P020P037nsss(0) <='0';
          end if;
        if(cVar1S22S99N019P033P030P003(0)='1' AND  E( 8)='0' AND A(13)='1' AND A( 1)='1' )then
          cVar2S22S99P069P012P017nsss(0) <='1';
          else
          cVar2S22S99P069P012P017nsss(0) <='0';
          end if;
        if(cVar1S23S99N019P033P030P012(0)='1' AND  A( 3)='1' )then
          cVar2S23S99P013nsss(0) <='1';
          else
          cVar2S23S99P013nsss(0) <='0';
          end if;
        if(cVar1S24S99N019P033P030P012(0)='1' AND  A( 3)='0' AND A(14)='1' )then
          cVar2S24S99N013P010nsss(0) <='1';
          else
          cVar2S24S99N013P010nsss(0) <='0';
          end if;
        if(cVar1S25S99N019P033P030P012(0)='1' AND  A( 3)='0' AND A(14)='0' AND A( 4)='1' )then
          cVar2S25S99N013N010P011nsss(0) <='1';
          else
          cVar2S25S99N013N010P011nsss(0) <='0';
          end if;
        if(cVar1S26S99N019P033P030P012(0)='1' AND  B( 0)='1' )then
          cVar2S26S99P037nsss(0) <='1';
          else
          cVar2S26S99P037nsss(0) <='0';
          end if;
        if(cVar1S27S99N019N033P036P027(0)='1' AND  B( 6)='0' AND E(11)='1' AND A( 5)='0' )then
          cVar2S27S99P025P057P009nsss(0) <='1';
          else
          cVar2S27S99P025P057P009nsss(0) <='0';
          end if;
        if(cVar1S28S99N019N033P036P027(0)='1' AND  B( 6)='0' AND E(11)='0' AND B( 3)='0' )then
          cVar2S28S99P025N057P031nsss(0) <='1';
          else
          cVar2S28S99P025N057P031nsss(0) <='0';
          end if;
        if(cVar1S29S99N019N033P036P027(0)='1' AND  B( 6)='1' AND D( 5)='0' )then
          cVar2S29S99P025P046nsss(0) <='1';
          else
          cVar2S29S99P025P046nsss(0) <='0';
          end if;
        if(cVar1S30S99N019N033P036N027(0)='1' AND  B( 6)='1' AND A(17)='1' AND D( 5)='1' )then
          cVar2S30S99P025P004P046nsss(0) <='1';
          else
          cVar2S30S99P025P004P046nsss(0) <='0';
          end if;
        if(cVar1S31S99N019N033P036N027(0)='1' AND  B( 6)='1' AND A(17)='0' AND B(13)='0' )then
          cVar2S31S99P025N004P028nsss(0) <='1';
          else
          cVar2S31S99P025N004P028nsss(0) <='0';
          end if;
        if(cVar1S32S99N019N033P036N027(0)='1' AND  B( 6)='0' AND A(13)='1' AND A( 6)='0' )then
          cVar2S32S99N025P012P007nsss(0) <='1';
          else
          cVar2S32S99N025P012P007nsss(0) <='0';
          end if;
        if(cVar1S33S99N019N033P036P021(0)='1' AND  E(11)='0' AND A( 1)='0' AND A( 7)='0' )then
          cVar2S33S99P057P017P005nsss(0) <='1';
          else
          cVar2S33S99P057P017P005nsss(0) <='0';
          end if;
        if(cVar1S34S99N019N033P036P021(0)='1' AND  E(11)='1' AND B(12)='1' AND A( 2)='1' )then
          cVar2S34S99P057P030P015nsss(0) <='1';
          else
          cVar2S34S99P057P030P015nsss(0) <='0';
          end if;
        if(cVar1S35S99N019N033P036P021(0)='1' AND  A( 2)='1' AND A(10)='0' )then
          cVar2S35S99P015P018nsss(0) <='1';
          else
          cVar2S35S99P015P018nsss(0) <='0';
          end if;
        if(cVar1S36S99N019N033P036P021(0)='1' AND  A( 2)='0' AND D( 8)='0' AND D( 9)='0' )then
          cVar2S36S99N015P067P063nsss(0) <='1';
          else
          cVar2S36S99N015P067P063nsss(0) <='0';
          end if;
        if(cVar1S0S100P036P012P019P014(0)='1' AND  E( 1)='0' AND A( 7)='0' AND A( 3)='0' )then
          cVar2S0S100P064P005P013nsss(0) <='1';
          else
          cVar2S0S100P064P005P013nsss(0) <='0';
          end if;
        if(cVar1S1S100P036P012P019P014(0)='1' AND  E( 1)='0' AND A( 7)='1' AND D( 2)='1' )then
          cVar2S1S100P064P005P058nsss(0) <='1';
          else
          cVar2S1S100P064P005P058nsss(0) <='0';
          end if;
        if(cVar1S2S100P036P012P019P014(0)='1' AND  E( 1)='1' AND E( 0)='0' AND E(10)='0' )then
          cVar2S2S100P064P068P061nsss(0) <='1';
          else
          cVar2S2S100P064P068P061nsss(0) <='0';
          end if;
        if(cVar1S3S100P036P012P019N014(0)='1' AND  E( 6)='1' AND B( 1)='1' )then
          cVar2S3S100P044P035nsss(0) <='1';
          else
          cVar2S3S100P044P035nsss(0) <='0';
          end if;
        if(cVar1S4S100P036P012P019N014(0)='1' AND  E( 6)='1' AND B( 1)='0' AND B(11)='0' )then
          cVar2S4S100P044N035P032nsss(0) <='1';
          else
          cVar2S4S100P044N035P032nsss(0) <='0';
          end if;
        if(cVar1S5S100P036P012P019N014(0)='1' AND  E( 6)='0' AND D( 7)='1' AND D(15)='0' )then
          cVar2S5S100N044P038P039nsss(0) <='1';
          else
          cVar2S5S100N044P038P039nsss(0) <='0';
          end if;
        if(cVar1S6S100P036P012P019N014(0)='1' AND  E( 6)='0' AND D( 7)='0' )then
          cVar2S6S100N044N038psss(0) <='1';
          else
          cVar2S6S100N044N038psss(0) <='0';
          end if;
        if(cVar1S7S100P036P012P019P016(0)='1' AND  B( 4)='1' AND B( 0)='1' )then
          cVar2S7S100P029P037nsss(0) <='1';
          else
          cVar2S7S100P029P037nsss(0) <='0';
          end if;
        if(cVar1S8S100P036P012P019P016(0)='1' AND  B( 4)='1' AND B( 0)='0' AND B(10)='0' )then
          cVar2S8S100P029N037P034nsss(0) <='1';
          else
          cVar2S8S100P029N037P034nsss(0) <='0';
          end if;
        if(cVar1S9S100P036P012P019P016(0)='1' AND  B( 4)='0' AND B(10)='0' AND A( 8)='0' )then
          cVar2S9S100N029P034P003nsss(0) <='1';
          else
          cVar2S9S100N029P034P003nsss(0) <='0';
          end if;
        if(cVar1S10S100P036P012P019P016(0)='1' AND  B( 4)='0' AND B(10)='1' AND E( 0)='0' )then
          cVar2S10S100N029P034P068nsss(0) <='1';
          else
          cVar2S10S100N029P034P068nsss(0) <='0';
          end if;
        if(cVar1S11S100P036P012P019N016(0)='1' AND  E( 1)='0' AND E( 2)='0' )then
          cVar2S11S100P064P060nsss(0) <='1';
          else
          cVar2S11S100P064P060nsss(0) <='0';
          end if;
        if(cVar1S12S100P036P012P019N016(0)='1' AND  E( 1)='0' AND E( 2)='1' AND A(12)='1' )then
          cVar2S12S100P064P060P014nsss(0) <='1';
          else
          cVar2S12S100P064P060P014nsss(0) <='0';
          end if;
        if(cVar1S13S100P036P012P019N016(0)='1' AND  E( 1)='1' AND B( 0)='1' AND E( 8)='1' )then
          cVar2S13S100P064P037P069nsss(0) <='1';
          else
          cVar2S13S100P064P037P069nsss(0) <='0';
          end if;
        if(cVar1S14S100P036P012P018P066(0)='1' AND  E(10)='1' AND A( 1)='0' )then
          cVar2S14S100P061P017nsss(0) <='1';
          else
          cVar2S14S100P061P017nsss(0) <='0';
          end if;
        if(cVar1S15S100P036P012P018P066(0)='1' AND  E(10)='1' AND A( 1)='1' AND A( 2)='1' )then
          cVar2S15S100P061P017P015nsss(0) <='1';
          else
          cVar2S15S100P061P017P015nsss(0) <='0';
          end if;
        if(cVar1S16S100P036P012P018P066(0)='1' AND  E(10)='0' AND E( 9)='1' AND A( 1)='1' )then
          cVar2S16S100N061P065P017nsss(0) <='1';
          else
          cVar2S16S100N061P065P017nsss(0) <='0';
          end if;
        if(cVar1S17S100P036P012P018P066(0)='1' AND  E(10)='0' AND E( 9)='0' AND A( 9)='1' )then
          cVar2S17S100N061N065P001nsss(0) <='1';
          else
          cVar2S17S100N061N065P001nsss(0) <='0';
          end if;
        if(cVar1S18S100P036P012P018N066(0)='1' AND  E( 4)='1' AND D( 4)='0' )then
          cVar2S18S100P052P050nsss(0) <='1';
          else
          cVar2S18S100P052P050nsss(0) <='0';
          end if;
        if(cVar1S19S100P036P012P018N066(0)='1' AND  E( 4)='1' AND D( 4)='1' AND A( 2)='0' )then
          cVar2S19S100P052P050P015nsss(0) <='1';
          else
          cVar2S19S100P052P050P015nsss(0) <='0';
          end if;
        if(cVar1S20S100P036P012P018N066(0)='1' AND  E( 4)='0' AND D(11)='1' )then
          cVar2S20S100N052P055nsss(0) <='1';
          else
          cVar2S20S100N052P055nsss(0) <='0';
          end if;
        if(cVar1S21S100P036P012N018P043(0)='1' AND  D( 2)='1' AND A( 9)='1' )then
          cVar2S21S100P058P001nsss(0) <='1';
          else
          cVar2S21S100P058P001nsss(0) <='0';
          end if;
        if(cVar1S22S100P036P012N018P043(0)='1' AND  D( 2)='1' AND A( 9)='0' AND A(16)='0' )then
          cVar2S22S100P058N001P006nsss(0) <='1';
          else
          cVar2S22S100P058N001P006nsss(0) <='0';
          end if;
        if(cVar1S23S100P036P012N018P043(0)='1' AND  D( 2)='0' AND E(11)='1' AND A( 2)='1' )then
          cVar2S23S100N058P057P015nsss(0) <='1';
          else
          cVar2S23S100N058P057P015nsss(0) <='0';
          end if;
        if(cVar1S24S100P036P012N018P043(0)='1' AND  D( 1)='0' AND A( 3)='0' AND A( 2)='0' )then
          cVar2S24S100P062P013P015nsss(0) <='1';
          else
          cVar2S24S100P062P013P015nsss(0) <='0';
          end if;
        if(cVar1S25S100P036P006P053P033(0)='1' AND  B( 5)='1' )then
          cVar2S25S100P027nsss(0) <='1';
          else
          cVar2S25S100P027nsss(0) <='0';
          end if;
        if(cVar1S26S100P036P006P053P033(0)='1' AND  B( 5)='0' AND B( 0)='1' )then
          cVar2S26S100N027P037nsss(0) <='1';
          else
          cVar2S26S100N027P037nsss(0) <='0';
          end if;
        if(cVar1S27S100P036P006P053P033(0)='1' AND  B( 5)='0' AND B( 0)='0' AND E(11)='0' )then
          cVar2S27S100N027N037P057nsss(0) <='1';
          else
          cVar2S27S100N027N037P057nsss(0) <='0';
          end if;
        if(cVar1S28S100P036P006P053P033(0)='1' AND  A( 1)='0' AND B( 0)='0' )then
          cVar2S28S100P017P037nsss(0) <='1';
          else
          cVar2S28S100P017P037nsss(0) <='0';
          end if;
        if(cVar1S29S100P036N006P008P026(0)='1' AND  A(13)='0' )then
          cVar2S29S100P012nsss(0) <='1';
          else
          cVar2S29S100P012nsss(0) <='0';
          end if;
        if(cVar1S30S100P036N006P008N026(0)='1' AND  E( 4)='1' AND B( 4)='1' )then
          cVar2S30S100P052P029nsss(0) <='1';
          else
          cVar2S30S100P052P029nsss(0) <='0';
          end if;
        if(cVar1S31S100P036N006P008N026(0)='1' AND  E( 4)='1' AND B( 4)='0' AND A( 0)='0' )then
          cVar2S31S100P052N029P019nsss(0) <='1';
          else
          cVar2S31S100P052N029P019nsss(0) <='0';
          end if;
        if(cVar1S32S100P036N006P008N026(0)='1' AND  E( 4)='0' AND B( 4)='0' AND A(19)='1' )then
          cVar2S32S100N052P029P000nsss(0) <='1';
          else
          cVar2S32S100N052P029P000nsss(0) <='0';
          end if;
        if(cVar1S33S100P036N006N008P047(0)='1' AND  B( 7)='0' AND A( 7)='0' AND A( 4)='1' )then
          cVar2S33S100P023P005P011nsss(0) <='1';
          else
          cVar2S33S100P023P005P011nsss(0) <='0';
          end if;
        if(cVar1S34S100P036N006N008P047(0)='1' AND  B( 7)='0' AND A( 7)='1' AND E( 8)='1' )then
          cVar2S34S100P023P005P069nsss(0) <='1';
          else
          cVar2S34S100P023P005P069nsss(0) <='0';
          end if;
        if(cVar1S35S100P036N006N008P047(0)='1' AND  B( 7)='1' AND D( 6)='1' AND E( 8)='0' )then
          cVar2S35S100P023P042P069nsss(0) <='1';
          else
          cVar2S35S100P023P042P069nsss(0) <='0';
          end if;
        if(cVar1S36S100P036N006N008P047(0)='1' AND  A(13)='0' AND E( 1)='1' )then
          cVar2S36S100P012P064nsss(0) <='1';
          else
          cVar2S36S100P012P064nsss(0) <='0';
          end if;
        if(cVar1S0S101P036P005P023P029(0)='1' AND  A(19)='1' AND E( 8)='1' )then
          cVar2S0S101P000P069nsss(0) <='1';
          else
          cVar2S0S101P000P069nsss(0) <='0';
          end if;
        if(cVar1S1S101P036P005P023P029(0)='1' AND  A(19)='1' AND E( 8)='0' AND A(10)='1' )then
          cVar2S1S101P000N069P018nsss(0) <='1';
          else
          cVar2S1S101P000N069P018nsss(0) <='0';
          end if;
        if(cVar1S2S101P036P005P023P029(0)='1' AND  A(19)='0' AND E(11)='0' )then
          cVar2S2S101N000P057nsss(0) <='1';
          else
          cVar2S2S101N000P057nsss(0) <='0';
          end if;
        if(cVar1S3S101P036P005P023P029(0)='1' AND  A(19)='0' AND E(11)='1' AND D( 2)='1' )then
          cVar2S3S101N000P057P058nsss(0) <='1';
          else
          cVar2S3S101N000P057P058nsss(0) <='0';
          end if;
        if(cVar1S4S101P036P005P023P029(0)='1' AND  B( 5)='0' AND E( 2)='1' )then
          cVar2S4S101P027P060nsss(0) <='1';
          else
          cVar2S4S101P027P060nsss(0) <='0';
          end if;
        if(cVar1S5S101P036P005P023P029(0)='1' AND  B( 5)='0' AND E( 2)='0' AND D( 8)='0' )then
          cVar2S5S101P027N060P067nsss(0) <='1';
          else
          cVar2S5S101P027N060P067nsss(0) <='0';
          end if;
        if(cVar1S7S101P036P005P023N004(0)='1' AND  E( 9)='1' )then
          cVar2S7S101P065nsss(0) <='1';
          else
          cVar2S7S101P065nsss(0) <='0';
          end if;
        if(cVar1S8S101P036P005P069P013(0)='1' AND  B( 2)='0' AND A( 8)='1' )then
          cVar2S8S101P033P003nsss(0) <='1';
          else
          cVar2S8S101P033P003nsss(0) <='0';
          end if;
        if(cVar1S9S101P036P005P069P013(0)='1' AND  B( 2)='0' AND A( 8)='0' AND D( 0)='1' )then
          cVar2S9S101P033N003P066nsss(0) <='1';
          else
          cVar2S9S101P033N003P066nsss(0) <='0';
          end if;
        if(cVar1S11S101P036P005N069N032(0)='1' AND  D( 2)='0' AND A(14)='1' AND A( 1)='0' )then
          cVar2S11S101P058P010P017nsss(0) <='1';
          else
          cVar2S11S101P058P010P017nsss(0) <='0';
          end if;
        if(cVar1S12S101N036P014P061P069(0)='1' AND  A( 2)='1' )then
          cVar2S12S101P015nsss(0) <='1';
          else
          cVar2S12S101P015nsss(0) <='0';
          end if;
        if(cVar1S13S101N036P014P061P069(0)='1' AND  A( 2)='0' AND A( 1)='1' )then
          cVar2S13S101N015P017nsss(0) <='1';
          else
          cVar2S13S101N015P017nsss(0) <='0';
          end if;
        if(cVar1S14S101N036P014P061P069(0)='1' AND  A( 2)='0' AND A( 1)='0' AND D( 2)='0' )then
          cVar2S14S101N015N017P058nsss(0) <='1';
          else
          cVar2S14S101N015N017P058nsss(0) <='0';
          end if;
        if(cVar1S15S101N036P014P061N069(0)='1' AND  B( 4)='0' AND D( 1)='0' AND B(14)='0' )then
          cVar2S15S101P029P062P026nsss(0) <='1';
          else
          cVar2S15S101P029P062P026nsss(0) <='0';
          end if;
        if(cVar1S16S101N036P014P061N069(0)='1' AND  B( 4)='0' AND D( 1)='1' AND A(11)='1' )then
          cVar2S16S101P029P062P016nsss(0) <='1';
          else
          cVar2S16S101P029P062P016nsss(0) <='0';
          end if;
        if(cVar1S17S101N036P014P061N069(0)='1' AND  B( 4)='1' AND D( 3)='0' AND A( 4)='0' )then
          cVar2S17S101P029P054P011nsss(0) <='1';
          else
          cVar2S17S101P029P054P011nsss(0) <='0';
          end if;
        if(cVar1S18S101N036P014N061P069(0)='1' AND  D( 1)='1' AND B( 2)='1' AND D( 0)='0' )then
          cVar2S18S101P062P033P066nsss(0) <='1';
          else
          cVar2S18S101P062P033P066nsss(0) <='0';
          end if;
        if(cVar1S19S101N036P014N061P069(0)='1' AND  D( 1)='1' AND B( 2)='0' AND E( 0)='1' )then
          cVar2S19S101P062N033P068nsss(0) <='1';
          else
          cVar2S19S101P062N033P068nsss(0) <='0';
          end if;
        if(cVar1S20S101N036P014N061P069(0)='1' AND  D( 1)='0' AND D(14)='1' )then
          cVar2S20S101N062P043nsss(0) <='1';
          else
          cVar2S20S101N062P043nsss(0) <='0';
          end if;
        if(cVar1S21S101N036P014N061P069(0)='1' AND  B( 8)='0' AND A(16)='1' AND B( 0)='1' )then
          cVar2S21S101P021P006P037nsss(0) <='1';
          else
          cVar2S21S101P021P006P037nsss(0) <='0';
          end if;
        if(cVar1S22S101N036P014N061P069(0)='1' AND  B( 8)='0' AND A(16)='0' AND E(11)='1' )then
          cVar2S22S101P021N006P057nsss(0) <='1';
          else
          cVar2S22S101P021N006P057nsss(0) <='0';
          end if;
        if(cVar1S23S101N036N014P012P023(0)='1' AND  A(10)='1' AND E( 1)='1' AND A( 2)='0' )then
          cVar2S23S101P018P064P015nsss(0) <='1';
          else
          cVar2S23S101P018P064P015nsss(0) <='0';
          end if;
        if(cVar1S24S101N036N014P012P023(0)='1' AND  A(10)='1' AND E( 1)='0' AND E( 8)='1' )then
          cVar2S24S101P018N064P069nsss(0) <='1';
          else
          cVar2S24S101P018N064P069nsss(0) <='0';
          end if;
        if(cVar1S25S101N036N014P012P023(0)='1' AND  A(10)='0' AND B( 2)='1' )then
          cVar2S25S101N018P033nsss(0) <='1';
          else
          cVar2S25S101N018P033nsss(0) <='0';
          end if;
        if(cVar1S26S101N036N014P012P023(0)='1' AND  A(10)='0' AND B( 2)='0' AND A( 4)='1' )then
          cVar2S26S101N018N033P011nsss(0) <='1';
          else
          cVar2S26S101N018N033P011nsss(0) <='0';
          end if;
        if(cVar1S27S101N036N014P012P023(0)='1' AND  A(14)='0' AND A(11)='1' )then
          cVar2S27S101P010P016nsss(0) <='1';
          else
          cVar2S27S101P010P016nsss(0) <='0';
          end if;
        if(cVar1S28S101N036N014N012P015(0)='1' AND  D( 2)='0' AND A(11)='1' )then
          cVar2S28S101P058P016nsss(0) <='1';
          else
          cVar2S28S101P058P016nsss(0) <='0';
          end if;
        if(cVar1S29S101N036N014N012P015(0)='1' AND  D( 2)='0' AND A(11)='0' AND B( 3)='1' )then
          cVar2S29S101P058N016P031nsss(0) <='1';
          else
          cVar2S29S101P058N016P031nsss(0) <='0';
          end if;
        if(cVar1S30S101N036N014N012P015(0)='1' AND  D( 2)='1' AND E(10)='1' AND A(11)='1' )then
          cVar2S30S101P058P061P016nsss(0) <='1';
          else
          cVar2S30S101P058P061P016nsss(0) <='0';
          end if;
        if(cVar1S31S101N036N014N012P015(0)='1' AND  E( 6)='1' )then
          cVar2S31S101P044nsss(0) <='1';
          else
          cVar2S31S101P044nsss(0) <='0';
          end if;
        if(cVar1S0S102P036P016P030P031(0)='1' AND  D(10)='1' )then
          cVar2S0S102P059nsss(0) <='1';
          else
          cVar2S0S102P059nsss(0) <='0';
          end if;
        if(cVar1S1S102P036P016P030P031(0)='1' AND  D(10)='0' AND E( 9)='0' AND B( 2)='0' )then
          cVar2S1S102N059P065P033nsss(0) <='1';
          else
          cVar2S1S102N059P065P033nsss(0) <='0';
          end if;
        if(cVar1S2S102P036P016P030P031(0)='1' AND  D(10)='0' AND E( 9)='1' AND D( 3)='0' )then
          cVar2S2S102N059P065P054nsss(0) <='1';
          else
          cVar2S2S102N059P065P054nsss(0) <='0';
          end if;
        if(cVar1S3S102P036P016P030P031(0)='1' AND  A( 5)='0' AND E( 0)='0' AND A( 2)='1' )then
          cVar2S3S102P009P068P015nsss(0) <='1';
          else
          cVar2S3S102P009P068P015nsss(0) <='0';
          end if;
        if(cVar1S4S102P036P016N030P028(0)='1' AND  D(11)='1' AND E( 3)='0' AND B( 1)='0' )then
          cVar2S4S102P055P056P035nsss(0) <='1';
          else
          cVar2S4S102P055P056P035nsss(0) <='0';
          end if;
        if(cVar1S5S102P036P016N030P028(0)='1' AND  D(11)='1' AND E( 3)='1' AND A(14)='0' )then
          cVar2S5S102P055P056P010nsss(0) <='1';
          else
          cVar2S5S102P055P056P010nsss(0) <='0';
          end if;
        if(cVar1S6S102P036P016N030P028(0)='1' AND  D(11)='0' AND A( 3)='1' AND A( 8)='0' )then
          cVar2S6S102N055P013P003nsss(0) <='1';
          else
          cVar2S6S102N055P013P003nsss(0) <='0';
          end if;
        if(cVar1S7S102P036P016N030P028(0)='1' AND  D(11)='0' AND A( 3)='0' AND E(14)='1' )then
          cVar2S7S102N055N013P045nsss(0) <='1';
          else
          cVar2S7S102N055N013P045nsss(0) <='0';
          end if;
        if(cVar1S8S102P036P016N030N028(0)='1' AND  A( 4)='0' AND A( 3)='0' AND D(11)='0' )then
          cVar2S8S102P011P013P055nsss(0) <='1';
          else
          cVar2S8S102P011P013P055nsss(0) <='0';
          end if;
        if(cVar1S9S102P036P016N030N028(0)='1' AND  A( 4)='0' AND A( 3)='1' AND A(13)='1' )then
          cVar2S9S102P011P013P012nsss(0) <='1';
          else
          cVar2S9S102P011P013P012nsss(0) <='0';
          end if;
        if(cVar1S10S102P036P016N030N028(0)='1' AND  A( 4)='1' AND A( 8)='1' AND A( 1)='1' )then
          cVar2S10S102P011P003P017nsss(0) <='1';
          else
          cVar2S10S102P011P003P017nsss(0) <='0';
          end if;
        if(cVar1S11S102P036P016P014P039(0)='1' AND  A( 1)='1' AND D( 9)='1' )then
          cVar2S11S102P017P063nsss(0) <='1';
          else
          cVar2S11S102P017P063nsss(0) <='0';
          end if;
        if(cVar1S12S102P036P016P014P039(0)='1' AND  A( 1)='1' AND D( 9)='0' AND E( 8)='1' )then
          cVar2S12S102P017N063P069nsss(0) <='1';
          else
          cVar2S12S102P017N063P069nsss(0) <='0';
          end if;
        if(cVar1S13S102P036P016P014P039(0)='1' AND  A( 1)='0' AND E( 8)='0' )then
          cVar2S13S102N017P069nsss(0) <='1';
          else
          cVar2S13S102N017P069nsss(0) <='0';
          end if;
        if(cVar1S14S102P036P016P014P039(0)='1' AND  A( 1)='0' AND E( 8)='1' AND B( 2)='1' )then
          cVar2S14S102N017P069P033nsss(0) <='1';
          else
          cVar2S14S102N017P069P033nsss(0) <='0';
          end if;
        if(cVar1S15S102P036P016N014P037(0)='1' AND  B(12)='1' AND E(11)='1' )then
          cVar2S15S102P030P057nsss(0) <='1';
          else
          cVar2S15S102P030P057nsss(0) <='0';
          end if;
        if(cVar1S16S102P036P016N014P037(0)='1' AND  B(12)='1' AND E(11)='0' AND A( 3)='0' )then
          cVar2S16S102P030N057P013nsss(0) <='1';
          else
          cVar2S16S102P030N057P013nsss(0) <='0';
          end if;
        if(cVar1S17S102P036P016N014P037(0)='1' AND  B(12)='0' AND E( 3)='0' AND A( 2)='1' )then
          cVar2S17S102N030P056P015nsss(0) <='1';
          else
          cVar2S17S102N030P056P015nsss(0) <='0';
          end if;
        if(cVar1S18S102P036P016N014N037(0)='1' AND  E( 3)='1' AND A(13)='1' )then
          cVar2S18S102P056P012nsss(0) <='1';
          else
          cVar2S18S102P056P012nsss(0) <='0';
          end if;
        if(cVar1S19S102P036P016N014N037(0)='1' AND  E( 3)='1' AND A(13)='0' AND A( 3)='1' )then
          cVar2S19S102P056N012P013nsss(0) <='1';
          else
          cVar2S19S102P056N012P013nsss(0) <='0';
          end if;
        if(cVar1S20S102P036P016N014N037(0)='1' AND  E( 3)='0' AND E( 6)='1' AND A( 3)='0' )then
          cVar2S20S102N056P044P013nsss(0) <='1';
          else
          cVar2S20S102N056P044P013nsss(0) <='0';
          end if;
        if(cVar1S22S102P036P000N069P013(0)='1' AND  D( 1)='1' )then
          cVar2S22S102P062nsss(0) <='1';
          else
          cVar2S22S102P062nsss(0) <='0';
          end if;
        if(cVar1S23S102P036P000N069P013(0)='1' AND  D( 1)='0' AND A(10)='1' AND A( 2)='1' )then
          cVar2S23S102N062P018P015nsss(0) <='1';
          else
          cVar2S23S102N062P018P015nsss(0) <='0';
          end if;
        if(cVar1S24S102P036N000P030P037(0)='1' AND  B(10)='0' AND B(11)='0' )then
          cVar2S24S102P034P032nsss(0) <='1';
          else
          cVar2S24S102P034P032nsss(0) <='0';
          end if;
        if(cVar1S25S102P036N000P030P037(0)='1' AND  E( 9)='1' )then
          cVar2S25S102P065nsss(0) <='1';
          else
          cVar2S25S102P065nsss(0) <='0';
          end if;
        if(cVar1S26S102P036N000P030P037(0)='1' AND  E( 9)='0' AND E(11)='1' )then
          cVar2S26S102N065P057nsss(0) <='1';
          else
          cVar2S26S102N065P057nsss(0) <='0';
          end if;
        if(cVar1S27S102P036N000N030P057(0)='1' AND  A(15)='1' AND B(14)='1' )then
          cVar2S27S102P008P026nsss(0) <='1';
          else
          cVar2S27S102P008P026nsss(0) <='0';
          end if;
        if(cVar1S28S102P036N000N030P057(0)='1' AND  A(15)='1' AND B(14)='0' AND B( 3)='0' )then
          cVar2S28S102P008N026P031nsss(0) <='1';
          else
          cVar2S28S102P008N026P031nsss(0) <='0';
          end if;
        if(cVar1S29S102P036N000N030P057(0)='1' AND  A(15)='0' AND A( 4)='1' AND A( 5)='1' )then
          cVar2S29S102N008P011P009nsss(0) <='1';
          else
          cVar2S29S102N008P011P009nsss(0) <='0';
          end if;
        if(cVar1S30S102P036N000N030P057(0)='1' AND  D( 2)='1' AND A(10)='0' )then
          cVar2S30S102P058P018nsss(0) <='1';
          else
          cVar2S30S102P058P018nsss(0) <='0';
          end if;
        if(cVar1S31S102P036N000N030P057(0)='1' AND  D( 2)='0' AND B( 3)='1' AND D( 8)='0' )then
          cVar2S31S102N058P031P067nsss(0) <='1';
          else
          cVar2S31S102N058P031P067nsss(0) <='0';
          end if;
        if(cVar1S0S103P036P001P023P043(0)='1' AND  A( 1)='0' AND A(13)='0' )then
          cVar2S0S103P017P012nsss(0) <='1';
          else
          cVar2S0S103P017P012nsss(0) <='0';
          end if;
        if(cVar1S1S103P036P001P023P043(0)='1' AND  A( 1)='1' AND A( 0)='1' )then
          cVar2S1S103P017P019nsss(0) <='1';
          else
          cVar2S1S103P017P019nsss(0) <='0';
          end if;
        if(cVar1S2S103P036P001P023N043(0)='1' AND  E(14)='0' AND D( 7)='0' )then
          cVar2S2S103P045P038nsss(0) <='1';
          else
          cVar2S2S103P045P038nsss(0) <='0';
          end if;
        if(cVar1S3S103P036P001P023N043(0)='1' AND  E(14)='0' AND D( 7)='1' AND A( 0)='1' )then
          cVar2S3S103P045P038P019nsss(0) <='1';
          else
          cVar2S3S103P045P038P019nsss(0) <='0';
          end if;
        if(cVar1S4S103P036P001P023N043(0)='1' AND  E(14)='1' AND A(11)='1' AND A(10)='0' )then
          cVar2S4S103P045P016P018nsss(0) <='1';
          else
          cVar2S4S103P045P016P018nsss(0) <='0';
          end if;
        if(cVar1S5S103P036P001P023P042(0)='1' AND  E( 8)='0' )then
          cVar2S5S103P069nsss(0) <='1';
          else
          cVar2S5S103P069nsss(0) <='0';
          end if;
        if(cVar1S8S103P036P001N034N033(0)='1' AND  E( 0)='1' AND B( 0)='0' AND D( 8)='0' )then
          cVar2S8S103P068P037P067nsss(0) <='1';
          else
          cVar2S8S103P068P037P067nsss(0) <='0';
          end if;
        if(cVar1S9S103N036P011P040P010(0)='1' AND  A( 6)='0' AND D( 4)='1' )then
          cVar2S9S103P007P050nsss(0) <='1';
          else
          cVar2S9S103P007P050nsss(0) <='0';
          end if;
        if(cVar1S10S103N036P011P040P010(0)='1' AND  A( 6)='0' AND D( 4)='0' AND E( 4)='0' )then
          cVar2S10S103P007N050P052nsss(0) <='1';
          else
          cVar2S10S103P007N050P052nsss(0) <='0';
          end if;
        if(cVar1S11S103N036P011P040P010(0)='1' AND  A( 6)='1' AND A(10)='1' AND E( 0)='1' )then
          cVar2S11S103P007P018P068nsss(0) <='1';
          else
          cVar2S11S103P007P018P068nsss(0) <='0';
          end if;
        if(cVar1S12S103N036P011P040P010(0)='1' AND  A( 6)='1' AND A(10)='0' AND D( 1)='1' )then
          cVar2S12S103P007N018P062nsss(0) <='1';
          else
          cVar2S12S103P007N018P062nsss(0) <='0';
          end if;
        if(cVar1S13S103N036P011P040P010(0)='1' AND  E( 4)='1' AND A( 0)='0' )then
          cVar2S13S103P052P019nsss(0) <='1';
          else
          cVar2S13S103P052P019nsss(0) <='0';
          end if;
        if(cVar1S14S103N036P011P040P010(0)='1' AND  E( 4)='0' AND D( 9)='1' AND A( 2)='0' )then
          cVar2S14S103N052P063P015nsss(0) <='1';
          else
          cVar2S14S103N052P063P015nsss(0) <='0';
          end if;
        if(cVar1S16S103N036P011P040N038(0)='1' AND  A(14)='1' )then
          cVar2S16S103P010nsss(0) <='1';
          else
          cVar2S16S103P010nsss(0) <='0';
          end if;
        if(cVar1S17S103N036N011P016P055(0)='1' AND  A(13)='1' AND A( 3)='0' )then
          cVar2S17S103P012P013nsss(0) <='1';
          else
          cVar2S17S103P012P013nsss(0) <='0';
          end if;
        if(cVar1S18S103N036N011P016P055(0)='1' AND  A(13)='1' AND A( 3)='1' AND A( 1)='1' )then
          cVar2S18S103P012P013P017nsss(0) <='1';
          else
          cVar2S18S103P012P013P017nsss(0) <='0';
          end if;
        if(cVar1S19S103N036N011P016P055(0)='1' AND  A(13)='0' AND A( 1)='1' )then
          cVar2S19S103N012P017nsss(0) <='1';
          else
          cVar2S19S103N012P017nsss(0) <='0';
          end if;
        if(cVar1S20S103N036N011P016P055(0)='1' AND  A(13)='0' AND A( 1)='0' AND A( 3)='1' )then
          cVar2S20S103N012N017P013nsss(0) <='1';
          else
          cVar2S20S103N012N017P013nsss(0) <='0';
          end if;
        if(cVar1S21S103N036N011P016P055(0)='1' AND  A(14)='0' AND A(10)='0' AND A( 1)='1' )then
          cVar2S21S103P010P018P017nsss(0) <='1';
          else
          cVar2S21S103P010P018P017nsss(0) <='0';
          end if;
        if(cVar1S22S103N036N011P016P055(0)='1' AND  A(14)='0' AND A(10)='1' AND B( 2)='1' )then
          cVar2S22S103P010P018P033nsss(0) <='1';
          else
          cVar2S22S103P010P018P033nsss(0) <='0';
          end if;
        if(cVar1S23S103N036N011N016P013(0)='1' AND  D( 8)='0' AND B(11)='0' )then
          cVar2S23S103P067P032nsss(0) <='1';
          else
          cVar2S23S103P067P032nsss(0) <='0';
          end if;
        if(cVar1S24S103N036N011N016P013(0)='1' AND  D( 8)='0' AND B(11)='1' AND B( 1)='1' )then
          cVar2S24S103P067P032P035nsss(0) <='1';
          else
          cVar2S24S103P067P032P035nsss(0) <='0';
          end if;
        if(cVar1S25S103N036N011N016P013(0)='1' AND  D( 8)='1' AND D(10)='1' )then
          cVar2S25S103P067P059nsss(0) <='1';
          else
          cVar2S25S103P067P059nsss(0) <='0';
          end if;
        if(cVar1S26S103N036N011N016P013(0)='1' AND  D( 8)='1' AND D(10)='0' AND E( 5)='1' )then
          cVar2S26S103P067N059P048nsss(0) <='1';
          else
          cVar2S26S103P067N059P048nsss(0) <='0';
          end if;
        if(cVar1S27S103N036N011N016N013(0)='1' AND  B( 3)='0' AND A( 6)='1' AND E(13)='1' )then
          cVar2S27S103P031P007P049nsss(0) <='1';
          else
          cVar2S27S103P031P007P049nsss(0) <='0';
          end if;
        if(cVar1S28S103N036N011N016N013(0)='1' AND  B( 3)='0' AND A( 6)='0' AND A( 9)='1' )then
          cVar2S28S103P031N007P001nsss(0) <='1';
          else
          cVar2S28S103P031N007P001nsss(0) <='0';
          end if;
        if(cVar1S29S103N036N011N016N013(0)='1' AND  B( 3)='1' AND A(14)='1' AND D( 8)='0' )then
          cVar2S29S103P031P010P067nsss(0) <='1';
          else
          cVar2S29S103P031P010P067nsss(0) <='0';
          end if;
        if(cVar1S0S104P036P051P026P048(0)='1' AND  A( 5)='1' )then
          cVar2S0S104P009nsss(0) <='1';
          else
          cVar2S0S104P009nsss(0) <='0';
          end if;
        if(cVar1S1S104P036P051P026P048(0)='1' AND  A( 5)='0' AND D( 4)='0' )then
          cVar2S1S104N009P050nsss(0) <='1';
          else
          cVar2S1S104N009P050nsss(0) <='0';
          end if;
        if(cVar1S2S104P036P051N026P028(0)='1' AND  A( 3)='1' )then
          cVar2S2S104P013nsss(0) <='1';
          else
          cVar2S2S104P013nsss(0) <='0';
          end if;
        if(cVar1S3S104P036P051N026P028(0)='1' AND  A( 3)='0' AND B(10)='1' )then
          cVar2S3S104N013P034nsss(0) <='1';
          else
          cVar2S3S104N013P034nsss(0) <='0';
          end if;
        if(cVar1S4S104P036P051N026P028(0)='1' AND  A( 3)='0' AND B(10)='0' AND D(10)='0' )then
          cVar2S4S104N013N034P059nsss(0) <='1';
          else
          cVar2S4S104N013N034P059nsss(0) <='0';
          end if;
        if(cVar1S5S104P036P051N026N028(0)='1' AND  E(11)='0' AND B( 3)='0' AND B( 5)='1' )then
          cVar2S5S104P057P031P027nsss(0) <='1';
          else
          cVar2S5S104P057P031P027nsss(0) <='0';
          end if;
        if(cVar1S6S104P036N051P053P009(0)='1' AND  E(13)='0' AND B(14)='0' AND A( 3)='0' )then
          cVar2S6S104P049P026P013nsss(0) <='1';
          else
          cVar2S6S104P049P026P013nsss(0) <='0';
          end if;
        if(cVar1S7S104P036N051P053P009(0)='1' AND  E(13)='0' AND B(14)='1' AND D( 4)='1' )then
          cVar2S7S104P049P026P050nsss(0) <='1';
          else
          cVar2S7S104P049P026P050nsss(0) <='0';
          end if;
        if(cVar1S8S104P036N051P053P009(0)='1' AND  E(13)='1' AND A( 6)='1' AND D( 5)='0' )then
          cVar2S8S104P049P007P046nsss(0) <='1';
          else
          cVar2S8S104P049P007P046nsss(0) <='0';
          end if;
        if(cVar1S9S104P036N051P053P009(0)='1' AND  E(13)='1' AND A( 6)='0' AND A( 7)='1' )then
          cVar2S9S104P049N007P005nsss(0) <='1';
          else
          cVar2S9S104P049N007P005nsss(0) <='0';
          end if;
        if(cVar1S10S104P036N051P053P009(0)='1' AND  D(13)='1' )then
          cVar2S10S104P047nsss(0) <='1';
          else
          cVar2S10S104P047nsss(0) <='0';
          end if;
        if(cVar1S11S104P036N051P053P009(0)='1' AND  D(13)='0' AND D( 4)='1' )then
          cVar2S11S104N047P050nsss(0) <='1';
          else
          cVar2S11S104N047P050nsss(0) <='0';
          end if;
        if(cVar1S12S104P036N051P053P026(0)='1' AND  E(11)='0' AND A(10)='0' )then
          cVar2S12S104P057P018nsss(0) <='1';
          else
          cVar2S12S104P057P018nsss(0) <='0';
          end if;
        if(cVar1S13S104P036N051P053P026(0)='1' AND  E(11)='0' AND A(10)='1' AND A(13)='1' )then
          cVar2S13S104P057P018P012nsss(0) <='1';
          else
          cVar2S13S104P057P018P012nsss(0) <='0';
          end if;
        if(cVar1S14S104P036N051P053P026(0)='1' AND  E(11)='1' AND A( 0)='0' AND A( 3)='1' )then
          cVar2S14S104P057P019P013nsss(0) <='1';
          else
          cVar2S14S104P057P019P013nsss(0) <='0';
          end if;
        if(cVar1S17S104P036P043N022N024(0)='1' AND  D( 1)='1' )then
          cVar2S17S104P062nsss(0) <='1';
          else
          cVar2S17S104P062nsss(0) <='0';
          end if;
        if(cVar1S18S104P036P043N022N024(0)='1' AND  D( 1)='0' AND A(11)='0' AND E( 8)='0' )then
          cVar2S18S104N062P016P069nsss(0) <='1';
          else
          cVar2S18S104N062P016P069nsss(0) <='0';
          end if;
        if(cVar1S19S104P036N043P045P038(0)='1' AND  A( 7)='0' AND A( 8)='1' AND E(13)='1' )then
          cVar2S19S104P005P003P049nsss(0) <='1';
          else
          cVar2S19S104P005P003P049nsss(0) <='0';
          end if;
        if(cVar1S20S104P036N043P045P038(0)='1' AND  A( 7)='1' AND B( 3)='0' AND E( 8)='1' )then
          cVar2S20S104P005P031P069nsss(0) <='1';
          else
          cVar2S20S104P005P031P069nsss(0) <='0';
          end if;
        if(cVar1S21S104P036N043P045P038(0)='1' AND  E( 7)='1' AND A( 0)='1' )then
          cVar2S21S104P040P019nsss(0) <='1';
          else
          cVar2S21S104P040P019nsss(0) <='0';
          end if;
        if(cVar1S22S104P036N043P045P016(0)='1' AND  B( 0)='1' )then
          cVar2S22S104P037nsss(0) <='1';
          else
          cVar2S22S104P037nsss(0) <='0';
          end if;
        if(cVar1S23S104P036N043P045N016(0)='1' AND  D( 0)='0' AND A(13)='0' AND D( 8)='0' )then
          cVar2S23S104P066P012P067nsss(0) <='1';
          else
          cVar2S23S104P066P012P067nsss(0) <='0';
          end if;
        if(cVar1S0S105P013P061P016P030(0)='1' AND  B( 2)='0' )then
          cVar2S0S105P033nsss(0) <='1';
          else
          cVar2S0S105P033nsss(0) <='0';
          end if;
        if(cVar1S1S105P013P061P016N030(0)='1' AND  D(11)='0' )then
          cVar2S1S105P055nsss(0) <='1';
          else
          cVar2S1S105P055nsss(0) <='0';
          end if;
        if(cVar1S2S105P013P061P016N030(0)='1' AND  D(11)='1' AND B( 3)='1' )then
          cVar2S2S105P055P031nsss(0) <='1';
          else
          cVar2S2S105P055P031nsss(0) <='0';
          end if;
        if(cVar1S3S105P013P061P016P033(0)='1' AND  A(12)='0' )then
          cVar2S3S105P014nsss(0) <='1';
          else
          cVar2S3S105P014nsss(0) <='0';
          end if;
        if(cVar1S4S105P013P061P016N033(0)='1' AND  B( 3)='1' )then
          cVar2S4S105P031nsss(0) <='1';
          else
          cVar2S4S105P031nsss(0) <='0';
          end if;
        if(cVar1S5S105P013P061P016N033(0)='1' AND  B( 3)='0' AND B(11)='1' AND E( 0)='1' )then
          cVar2S5S105N031P032P068nsss(0) <='1';
          else
          cVar2S5S105N031P032P068nsss(0) <='0';
          end if;
        if(cVar1S6S105P013P061P016N033(0)='1' AND  B( 3)='0' AND B(11)='0' AND D( 1)='1' )then
          cVar2S6S105N031N032P062nsss(0) <='1';
          else
          cVar2S6S105N031N032P062nsss(0) <='0';
          end if;
        if(cVar1S7S105P013N061P032P051(0)='1' AND  B(13)='1' AND A(10)='0' )then
          cVar2S7S105P028P018nsss(0) <='1';
          else
          cVar2S7S105P028P018nsss(0) <='0';
          end if;
        if(cVar1S8S105P013N061P032P051(0)='1' AND  B(13)='1' AND A(10)='1' AND A( 0)='0' )then
          cVar2S8S105P028P018P019nsss(0) <='1';
          else
          cVar2S8S105P028P018P019nsss(0) <='0';
          end if;
        if(cVar1S9S105P013N061P032P051(0)='1' AND  B(13)='0' AND B(14)='1' AND E(12)='1' )then
          cVar2S9S105N028P026P053nsss(0) <='1';
          else
          cVar2S9S105N028P026P053nsss(0) <='0';
          end if;
        if(cVar1S10S105P013N061P032P051(0)='1' AND  B(13)='0' AND B(14)='0' AND B( 4)='1' )then
          cVar2S10S105N028N026P029nsss(0) <='1';
          else
          cVar2S10S105N028N026P029nsss(0) <='0';
          end if;
        if(cVar1S11S105P013N061P032N051(0)='1' AND  B(13)='0' AND E(11)='1' )then
          cVar2S11S105P028P057nsss(0) <='1';
          else
          cVar2S11S105P028P057nsss(0) <='0';
          end if;
        if(cVar1S12S105P013N061P032N051(0)='1' AND  B(13)='0' AND E(11)='0' AND B( 6)='1' )then
          cVar2S12S105P028N057P025nsss(0) <='1';
          else
          cVar2S12S105P028N057P025nsss(0) <='0';
          end if;
        if(cVar1S13S105P013N061P032N051(0)='1' AND  B(13)='1' AND B(12)='0' AND A(11)='0' )then
          cVar2S13S105P028P030P016nsss(0) <='1';
          else
          cVar2S13S105P028P030P016nsss(0) <='0';
          end if;
        if(cVar1S14S105P013N061P032P063(0)='1' AND  A(10)='1' )then
          cVar2S14S105P018nsss(0) <='1';
          else
          cVar2S14S105P018nsss(0) <='0';
          end if;
        if(cVar1S15S105P013N061P032N063(0)='1' AND  A(12)='1' AND D( 2)='1' )then
          cVar2S15S105P014P058nsss(0) <='1';
          else
          cVar2S15S105P014P058nsss(0) <='0';
          end if;
        if(cVar1S16S105N013P036P002P011(0)='1' AND  D(12)='0' AND D( 7)='0' )then
          cVar2S16S105P051P038nsss(0) <='1';
          else
          cVar2S16S105P051P038nsss(0) <='0';
          end if;
        if(cVar1S17S105N013P036P002P011(0)='1' AND  D(12)='1' AND A(15)='1' )then
          cVar2S17S105P051P008nsss(0) <='1';
          else
          cVar2S17S105P051P008nsss(0) <='0';
          end if;
        if(cVar1S18S105N013P036P002P011(0)='1' AND  A( 8)='0' AND A( 1)='1' )then
          cVar2S18S105P003P017nsss(0) <='1';
          else
          cVar2S18S105P003P017nsss(0) <='0';
          end if;
        if(cVar1S19S105N013P036P002P011(0)='1' AND  A( 8)='0' AND A( 1)='0' AND D(12)='1' )then
          cVar2S19S105P003N017P051nsss(0) <='1';
          else
          cVar2S19S105P003N017P051nsss(0) <='0';
          end if;
        if(cVar1S20S105N013P036P002P011(0)='1' AND  A( 8)='1' AND A( 7)='1' )then
          cVar2S20S105P003P005nsss(0) <='1';
          else
          cVar2S20S105P003P005nsss(0) <='0';
          end if;
        if(cVar1S21S105N013P036P002P011(0)='1' AND  A( 8)='1' AND A( 7)='0' AND B(10)='1' )then
          cVar2S21S105P003N005P034nsss(0) <='1';
          else
          cVar2S21S105P003N005P034nsss(0) <='0';
          end if;
        if(cVar1S22S105N013P036P002P068(0)='1' AND  A(17)='0' AND B(10)='0' )then
          cVar2S22S105P004P034nsss(0) <='1';
          else
          cVar2S22S105P004P034nsss(0) <='0';
          end if;
        if(cVar1S23S105N013N036P028P055(0)='1' AND  D( 8)='1' )then
          cVar2S23S105P067nsss(0) <='1';
          else
          cVar2S23S105P067nsss(0) <='0';
          end if;
        if(cVar1S24S105N013N036P028P055(0)='1' AND  D( 8)='0' AND B( 1)='0' )then
          cVar2S24S105N067P035nsss(0) <='1';
          else
          cVar2S24S105N067P035nsss(0) <='0';
          end if;
        if(cVar1S25S105N013N036P028N055(0)='1' AND  D( 4)='1' AND B( 4)='0' )then
          cVar2S25S105P050P029nsss(0) <='1';
          else
          cVar2S25S105P050P029nsss(0) <='0';
          end if;
        if(cVar1S26S105N013N036P028N055(0)='1' AND  D( 4)='0' AND B(16)='1' )then
          cVar2S26S105N050P022nsss(0) <='1';
          else
          cVar2S26S105N050P022nsss(0) <='0';
          end if;
        if(cVar1S27S105N013N036N028P026(0)='1' AND  B( 8)='0' AND D( 6)='0' )then
          cVar2S27S105P021P042nsss(0) <='1';
          else
          cVar2S27S105P021P042nsss(0) <='0';
          end if;
        if(cVar1S28S105N013N036N028N026(0)='1' AND  B( 3)='0' AND B( 4)='1' AND A(10)='1' )then
          cVar2S28S105P031P029P018nsss(0) <='1';
          else
          cVar2S28S105P031P029P018nsss(0) <='0';
          end if;
        if(cVar1S29S105N013N036N028N026(0)='1' AND  B( 3)='1' AND D( 3)='1' AND A( 1)='1' )then
          cVar2S29S105P031P054P017nsss(0) <='1';
          else
          cVar2S29S105P031P054P017nsss(0) <='0';
          end if;
        if(cVar1S30S105N013N036N028N026(0)='1' AND  B( 3)='1' AND D( 3)='0' AND D( 2)='1' )then
          cVar2S30S105P031N054P058nsss(0) <='1';
          else
          cVar2S30S105P031N054P058nsss(0) <='0';
          end if;
        if(cVar1S0S106P036P064P002P048(0)='1' AND  A(15)='1' AND B( 0)='1' AND B(14)='0' )then
          cVar2S0S106P008P037P026nsss(0) <='1';
          else
          cVar2S0S106P008P037P026nsss(0) <='0';
          end if;
        if(cVar1S1S106P036P064P002P048(0)='1' AND  A(15)='1' AND B( 0)='0' AND E(12)='1' )then
          cVar2S1S106P008N037P053nsss(0) <='1';
          else
          cVar2S1S106P008N037P053nsss(0) <='0';
          end if;
        if(cVar1S2S106P036P064P002P048(0)='1' AND  A(15)='0' AND A( 0)='1' AND A( 2)='0' )then
          cVar2S2S106N008P019P015nsss(0) <='1';
          else
          cVar2S2S106N008P019P015nsss(0) <='0';
          end if;
        if(cVar1S3S106P036P064P002P048(0)='1' AND  A(15)='0' AND A( 0)='0' AND A(16)='0' )then
          cVar2S3S106N008N019P006nsss(0) <='1';
          else
          cVar2S3S106N008N019P006nsss(0) <='0';
          end if;
        if(cVar1S4S106P036P064P002P048(0)='1' AND  B(15)='1' )then
          cVar2S4S106P024nsss(0) <='1';
          else
          cVar2S4S106P024nsss(0) <='0';
          end if;
        if(cVar1S5S106P036P064P002P048(0)='1' AND  B(15)='0' AND B(14)='0' AND D( 9)='0' )then
          cVar2S5S106N024P026P063nsss(0) <='1';
          else
          cVar2S5S106N024P026P063nsss(0) <='0';
          end if;
        if(cVar1S6S106P036P064P002P012(0)='1' AND  A(14)='0' AND A( 1)='0' AND A(11)='1' )then
          cVar2S6S106P010P017P016nsss(0) <='1';
          else
          cVar2S6S106P010P017P016nsss(0) <='0';
          end if;
        if(cVar1S7S106P036P064P002P012(0)='1' AND  A(14)='0' AND A( 1)='1' AND D( 0)='1' )then
          cVar2S7S106P010P017P066nsss(0) <='1';
          else
          cVar2S7S106P010P017P066nsss(0) <='0';
          end if;
        if(cVar1S8S106P036N064P062P015(0)='1' AND  D(12)='1' AND D( 4)='0' )then
          cVar2S8S106P051P050nsss(0) <='1';
          else
          cVar2S8S106P051P050nsss(0) <='0';
          end if;
        if(cVar1S9S106P036N064P062P015(0)='1' AND  D(12)='0' AND E(12)='0' )then
          cVar2S9S106N051P053nsss(0) <='1';
          else
          cVar2S9S106N051P053nsss(0) <='0';
          end if;
        if(cVar1S10S106P036N064P062N015(0)='1' AND  B( 7)='1' AND A(16)='1' )then
          cVar2S10S106P023P006nsss(0) <='1';
          else
          cVar2S10S106P023P006nsss(0) <='0';
          end if;
        if(cVar1S11S106P036N064P062N015(0)='1' AND  B( 7)='1' AND A(16)='0' AND A(10)='1' )then
          cVar2S11S106P023N006P018nsss(0) <='1';
          else
          cVar2S11S106P023N006P018nsss(0) <='0';
          end if;
        if(cVar1S12S106P036N064P062N015(0)='1' AND  B( 7)='0' AND D( 6)='0' )then
          cVar2S12S106N023P042nsss(0) <='1';
          else
          cVar2S12S106N023P042nsss(0) <='0';
          end if;
        if(cVar1S13S106P036N064P062N015(0)='1' AND  B( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar2S13S106N023P042P021nsss(0) <='1';
          else
          cVar2S13S106N023P042P021nsss(0) <='0';
          end if;
        if(cVar1S14S106P036N064P062P042(0)='1' AND  E( 2)='1' AND D( 9)='0' AND A( 1)='0' )then
          cVar2S14S106P060P063P017nsss(0) <='1';
          else
          cVar2S14S106P060P063P017nsss(0) <='0';
          end if;
        if(cVar1S15S106P036N064P062P042(0)='1' AND  E( 2)='1' AND D( 9)='1' AND A( 1)='1' )then
          cVar2S15S106P060P063P017nsss(0) <='1';
          else
          cVar2S15S106P060P063P017nsss(0) <='0';
          end if;
        if(cVar1S16S106P036N064P062P042(0)='1' AND  E( 2)='0' AND E( 9)='1' AND B( 0)='1' )then
          cVar2S16S106N060P065P037nsss(0) <='1';
          else
          cVar2S16S106N060P065P037nsss(0) <='0';
          end if;
        if(cVar1S17S106P036N064P062P042(0)='1' AND  E( 2)='0' AND E( 9)='0' AND D(12)='1' )then
          cVar2S17S106N060N065P051nsss(0) <='1';
          else
          cVar2S17S106N060N065P051nsss(0) <='0';
          end if;
        if(cVar1S18S106P036P005P013P008(0)='1' AND  A(18)='1' AND A( 4)='1' )then
          cVar2S18S106P002P011nsss(0) <='1';
          else
          cVar2S18S106P002P011nsss(0) <='0';
          end if;
        if(cVar1S19S106P036P005P013P008(0)='1' AND  A(18)='1' AND A( 4)='0' AND A(10)='0' )then
          cVar2S19S106P002N011P018nsss(0) <='1';
          else
          cVar2S19S106P002N011P018nsss(0) <='0';
          end if;
        if(cVar1S20S106P036P005P013P008(0)='1' AND  A(18)='0' AND B( 2)='1' AND A( 6)='0' )then
          cVar2S20S106N002P033P007nsss(0) <='1';
          else
          cVar2S20S106N002P033P007nsss(0) <='0';
          end if;
        if(cVar1S21S106P036P005P013P008(0)='1' AND  A(18)='0' AND B( 2)='0' AND D(13)='0' )then
          cVar2S21S106N002N033P047nsss(0) <='1';
          else
          cVar2S21S106N002N033P047nsss(0) <='0';
          end if;
        if(cVar1S22S106P036P005P013P008(0)='1' AND  B( 2)='1' AND D( 8)='0' )then
          cVar2S22S106P033P067nsss(0) <='1';
          else
          cVar2S22S106P033P067nsss(0) <='0';
          end if;
        if(cVar1S23S106P036P005N013P061(0)='1' AND  D(10)='0' AND D( 2)='1' )then
          cVar2S23S106P059P058nsss(0) <='1';
          else
          cVar2S23S106P059P058nsss(0) <='0';
          end if;
        if(cVar1S24S106P036P005N013P061(0)='1' AND  D(10)='1' AND E( 2)='1' )then
          cVar2S24S106P059P060nsss(0) <='1';
          else
          cVar2S24S106P059P060nsss(0) <='0';
          end if;
        if(cVar1S25S106P036P005N013P061(0)='1' AND  D( 2)='0' AND D(10)='1' AND B( 1)='1' )then
          cVar2S25S106P058P059P035nsss(0) <='1';
          else
          cVar2S25S106P058P059P035nsss(0) <='0';
          end if;
        if(cVar1S26S106P036P005N013P061(0)='1' AND  D( 2)='0' AND D(10)='0' AND A( 4)='1' )then
          cVar2S26S106P058N059P011nsss(0) <='1';
          else
          cVar2S26S106P058N059P011nsss(0) <='0';
          end if;
        if(cVar1S27S106P036P005N013P061(0)='1' AND  D( 2)='1' AND A(12)='0' AND D( 9)='1' )then
          cVar2S27S106P058P014P063nsss(0) <='1';
          else
          cVar2S27S106P058P014P063nsss(0) <='0';
          end if;
        if(cVar1S29S106P036P005P031N020(0)='1' AND  E( 8)='1' AND E( 2)='1' )then
          cVar2S29S106P069P060nsss(0) <='1';
          else
          cVar2S29S106P069P060nsss(0) <='0';
          end if;
        if(cVar1S30S106P036P005P031N020(0)='1' AND  E( 8)='0' AND E(10)='1' )then
          cVar2S30S106N069P061nsss(0) <='1';
          else
          cVar2S30S106N069P061nsss(0) <='0';
          end if;
        if(cVar1S31S106P036P005P031N020(0)='1' AND  E( 8)='0' AND E(10)='0' AND B(14)='1' )then
          cVar2S31S106N069N061P026nsss(0) <='1';
          else
          cVar2S31S106N069N061P026nsss(0) <='0';
          end if;
        if(cVar1S0S107P036P005P019P047(0)='1' AND  E(10)='0' AND B( 0)='0' AND D(10)='0' )then
          cVar2S0S107P061P037P059nsss(0) <='1';
          else
          cVar2S0S107P061P037P059nsss(0) <='0';
          end if;
        if(cVar1S1S107P036P005P019P047(0)='1' AND  E(10)='0' AND B( 0)='1' AND D( 0)='0' )then
          cVar2S1S107P061P037P066nsss(0) <='1';
          else
          cVar2S1S107P061P037P066nsss(0) <='0';
          end if;
        if(cVar1S2S107P036P005P019P047(0)='1' AND  E(10)='1' AND B( 0)='1' )then
          cVar2S2S107P061P037nsss(0) <='1';
          else
          cVar2S2S107P061P037nsss(0) <='0';
          end if;
        if(cVar1S3S107P036P005P019P047(0)='1' AND  E(13)='1' AND E( 8)='1' )then
          cVar2S3S107P049P069nsss(0) <='1';
          else
          cVar2S3S107P049P069nsss(0) <='0';
          end if;
        if(cVar1S4S107P036P005N019P048(0)='1' AND  A(13)='0' AND B(11)='0' AND E(12)='1' )then
          cVar2S4S107P012P032P053nsss(0) <='1';
          else
          cVar2S4S107P012P032P053nsss(0) <='0';
          end if;
        if(cVar1S5S107P036P005N019P048(0)='1' AND  A(13)='0' AND B(11)='1' AND A(10)='1' )then
          cVar2S5S107P012P032P018nsss(0) <='1';
          else
          cVar2S5S107P012P032P018nsss(0) <='0';
          end if;
        if(cVar1S6S107P036P005N019P048(0)='1' AND  A(13)='1' AND E( 3)='1' )then
          cVar2S6S107P012P056nsss(0) <='1';
          else
          cVar2S6S107P012P056nsss(0) <='0';
          end if;
        if(cVar1S7S107P036P005N019P048(0)='1' AND  A(13)='1' AND E( 3)='0' AND B(11)='1' )then
          cVar2S7S107P012N056P032nsss(0) <='1';
          else
          cVar2S7S107P012N056P032nsss(0) <='0';
          end if;
        if(cVar1S8S107P036P005N019P048(0)='1' AND  B(14)='1' )then
          cVar2S8S107P026nsss(0) <='1';
          else
          cVar2S8S107P026nsss(0) <='0';
          end if;
        if(cVar1S9S107P036P005N019P048(0)='1' AND  B(14)='0' AND A( 5)='1' AND B( 5)='0' )then
          cVar2S9S107N026P009P027nsss(0) <='1';
          else
          cVar2S9S107N026P009P027nsss(0) <='0';
          end if;
        if(cVar1S10S107P036P005P031P069(0)='1' AND  B( 2)='0' AND A( 8)='1' )then
          cVar2S10S107P033P003nsss(0) <='1';
          else
          cVar2S10S107P033P003nsss(0) <='0';
          end if;
        if(cVar1S11S107P036P005P031P069(0)='1' AND  B( 2)='0' AND A( 8)='0' AND A(11)='0' )then
          cVar2S11S107P033N003P016nsss(0) <='1';
          else
          cVar2S11S107P033N003P016nsss(0) <='0';
          end if;
        if(cVar1S12S107P036P005P031N069(0)='1' AND  B(11)='1' )then
          cVar2S12S107P032nsss(0) <='1';
          else
          cVar2S12S107P032nsss(0) <='0';
          end if;
        if(cVar1S13S107P036P005P031N069(0)='1' AND  B(11)='0' AND D( 2)='0' AND A(14)='1' )then
          cVar2S13S107N032P058P010nsss(0) <='1';
          else
          cVar2S13S107N032P058P010nsss(0) <='0';
          end if;
        if(cVar1S14S107N036P064P019P059(0)='1' AND  A(14)='0' AND A( 3)='0' )then
          cVar2S14S107P010P013nsss(0) <='1';
          else
          cVar2S14S107P010P013nsss(0) <='0';
          end if;
        if(cVar1S15S107N036P064P019P059(0)='1' AND  A(14)='0' AND A( 3)='1' AND B(11)='1' )then
          cVar2S15S107P010P013P032nsss(0) <='1';
          else
          cVar2S15S107P010P013P032nsss(0) <='0';
          end if;
        if(cVar1S16S107N036P064P019N059(0)='1' AND  B(12)='1' AND D( 9)='0' )then
          cVar2S16S107P030P063nsss(0) <='1';
          else
          cVar2S16S107P030P063nsss(0) <='0';
          end if;
        if(cVar1S17S107N036P064P019N059(0)='1' AND  B(12)='0' AND A( 1)='0' )then
          cVar2S17S107N030P017nsss(0) <='1';
          else
          cVar2S17S107N030P017nsss(0) <='0';
          end if;
        if(cVar1S18S107N036P064P019N059(0)='1' AND  B(12)='0' AND A( 1)='1' AND A( 7)='1' )then
          cVar2S18S107N030P017P005nsss(0) <='1';
          else
          cVar2S18S107N030P017P005nsss(0) <='0';
          end if;
        if(cVar1S19S107N036P064N019P056(0)='1' AND  A( 8)='1' AND D( 1)='1' )then
          cVar2S19S107P003P062nsss(0) <='1';
          else
          cVar2S19S107P003P062nsss(0) <='0';
          end if;
        if(cVar1S20S107N036P064N019P056(0)='1' AND  A( 8)='0' AND A( 1)='1' )then
          cVar2S20S107N003P017nsss(0) <='1';
          else
          cVar2S20S107N003P017nsss(0) <='0';
          end if;
        if(cVar1S21S107N036P064N019P056(0)='1' AND  B( 1)='1' AND D(11)='1' )then
          cVar2S21S107P035P055nsss(0) <='1';
          else
          cVar2S21S107P035P055nsss(0) <='0';
          end if;
        if(cVar1S22S107N036P064N019P056(0)='1' AND  B( 1)='1' AND D(11)='0' AND D( 9)='0' )then
          cVar2S22S107P035N055P063nsss(0) <='1';
          else
          cVar2S22S107P035N055P063nsss(0) <='0';
          end if;
        if(cVar1S23S107N036P064N019P056(0)='1' AND  B( 1)='0' AND A( 5)='1' )then
          cVar2S23S107N035P009nsss(0) <='1';
          else
          cVar2S23S107N035P009nsss(0) <='0';
          end if;
        if(cVar1S24S107N036P064N019P056(0)='1' AND  B( 1)='0' AND A( 5)='0' AND A(12)='1' )then
          cVar2S24S107N035N009P014nsss(0) <='1';
          else
          cVar2S24S107N035N009P014nsss(0) <='0';
          end if;
        if(cVar1S25S107N036N064P051P057(0)='1' AND  D( 0)='1' AND D( 2)='0' )then
          cVar2S25S107P066P058nsss(0) <='1';
          else
          cVar2S25S107P066P058nsss(0) <='0';
          end if;
        if(cVar1S26S107N036N064P051P057(0)='1' AND  D( 0)='0' AND B(15)='1' )then
          cVar2S26S107N066P024nsss(0) <='1';
          else
          cVar2S26S107N066P024nsss(0) <='0';
          end if;
        if(cVar1S27S107N036N064P051P057(0)='1' AND  D( 0)='0' AND B(15)='0' AND A( 2)='1' )then
          cVar2S27S107N066N024P015nsss(0) <='1';
          else
          cVar2S27S107N066N024P015nsss(0) <='0';
          end if;
        if(cVar1S28S107N036N064P051P057(0)='1' AND  E(12)='1' AND B(12)='1' )then
          cVar2S28S107P053P030nsss(0) <='1';
          else
          cVar2S28S107P053P030nsss(0) <='0';
          end if;
        if(cVar1S29S107N036N064P051P057(0)='1' AND  E(12)='1' AND B(12)='0' AND A(14)='1' )then
          cVar2S29S107P053N030P010nsss(0) <='1';
          else
          cVar2S29S107P053N030P010nsss(0) <='0';
          end if;
        if(cVar1S30S107N036N064N051P053(0)='1' AND  B( 7)='1' AND A(16)='1' AND A(10)='0' )then
          cVar2S30S107P023P006P018nsss(0) <='1';
          else
          cVar2S30S107P023P006P018nsss(0) <='0';
          end if;
        if(cVar1S31S107N036N064N051P053(0)='1' AND  B( 7)='1' AND A(16)='0' AND D( 6)='1' )then
          cVar2S31S107P023N006P042nsss(0) <='1';
          else
          cVar2S31S107P023N006P042nsss(0) <='0';
          end if;
        if(cVar1S32S107N036N064N051P053(0)='1' AND  B( 7)='0' AND D(10)='1' AND B(12)='1' )then
          cVar2S32S107N023P059P030nsss(0) <='1';
          else
          cVar2S32S107N023P059P030nsss(0) <='0';
          end if;
        if(cVar1S33S107N036N064N051P053(0)='1' AND  B(14)='0' AND E(11)='0' AND A( 4)='1' )then
          cVar2S33S107P026P057P011nsss(0) <='1';
          else
          cVar2S33S107P026P057P011nsss(0) <='0';
          end if;
        if(cVar1S0S108P064P012P031P054(0)='1' AND  B(12)='0' AND E(11)='0' )then
          cVar2S0S108P030P057nsss(0) <='1';
          else
          cVar2S0S108P030P057nsss(0) <='0';
          end if;
        if(cVar1S1S108P064P012P031P054(0)='1' AND  B(12)='0' AND E(11)='1' AND E(10)='0' )then
          cVar2S1S108P030P057P061nsss(0) <='1';
          else
          cVar2S1S108P030P057P061nsss(0) <='0';
          end if;
        if(cVar1S2S108P064P012P031P054(0)='1' AND  B(12)='1' AND B( 4)='0' AND E(11)='1' )then
          cVar2S2S108P030P029P057nsss(0) <='1';
          else
          cVar2S2S108P030P029P057nsss(0) <='0';
          end if;
        if(cVar1S3S108P064P012P031P054(0)='1' AND  B( 4)='1' AND A(15)='1' )then
          cVar2S3S108P029P008nsss(0) <='1';
          else
          cVar2S3S108P029P008nsss(0) <='0';
          end if;
        if(cVar1S4S108P064P012P031P054(0)='1' AND  B( 4)='1' AND A(15)='0' AND A(14)='1' )then
          cVar2S4S108P029N008P010nsss(0) <='1';
          else
          cVar2S4S108P029N008P010nsss(0) <='0';
          end if;
        if(cVar1S5S108P064P012P031P054(0)='1' AND  B( 4)='0' AND E(10)='1' )then
          cVar2S5S108N029P061nsss(0) <='1';
          else
          cVar2S5S108N029P061nsss(0) <='0';
          end if;
        if(cVar1S6S108P064P012P031P054(0)='1' AND  B( 4)='0' AND E(10)='0' AND B(12)='1' )then
          cVar2S6S108N029N061P030nsss(0) <='1';
          else
          cVar2S6S108N029N061P030nsss(0) <='0';
          end if;
        if(cVar1S7S108P064P012P031P005(0)='1' AND  D( 3)='1' AND A( 2)='1' AND A( 1)='0' )then
          cVar2S7S108P054P015P017nsss(0) <='1';
          else
          cVar2S7S108P054P015P017nsss(0) <='0';
          end if;
        if(cVar1S8S108P064P012P031P005(0)='1' AND  D( 3)='1' AND A( 2)='0' AND D( 0)='1' )then
          cVar2S8S108P054N015P066nsss(0) <='1';
          else
          cVar2S8S108P054N015P066nsss(0) <='0';
          end if;
        if(cVar1S9S108P064P012P031P005(0)='1' AND  D( 3)='0' AND E(11)='1' AND B(12)='0' )then
          cVar2S9S108N054P057P030nsss(0) <='1';
          else
          cVar2S9S108N054P057P030nsss(0) <='0';
          end if;
        if(cVar1S10S108P064P012P031P005(0)='1' AND  E( 0)='1' )then
          cVar2S10S108P068nsss(0) <='1';
          else
          cVar2S10S108P068nsss(0) <='0';
          end if;
        if(cVar1S11S108P064P012P030P032(0)='1' AND  E( 3)='0' AND B( 2)='0' )then
          cVar2S11S108P056P033nsss(0) <='1';
          else
          cVar2S11S108P056P033nsss(0) <='0';
          end if;
        if(cVar1S12S108P064P012P030P032(0)='1' AND  E( 3)='0' AND B( 2)='1' AND A( 0)='1' )then
          cVar2S12S108P056P033P019nsss(0) <='1';
          else
          cVar2S12S108P056P033P019nsss(0) <='0';
          end if;
        if(cVar1S13S108P064P012P030P032(0)='1' AND  E( 3)='1' AND A(14)='0' AND A(10)='1' )then
          cVar2S13S108P056P010P018nsss(0) <='1';
          else
          cVar2S13S108P056P010P018nsss(0) <='0';
          end if;
        if(cVar1S14S108P064P012P030P032(0)='1' AND  E(10)='1' AND D(11)='0' )then
          cVar2S14S108P061P055nsss(0) <='1';
          else
          cVar2S14S108P061P055nsss(0) <='0';
          end if;
        if(cVar1S15S108P064P012P030P032(0)='1' AND  E(10)='0' AND A( 1)='1' )then
          cVar2S15S108N061P017nsss(0) <='1';
          else
          cVar2S15S108N061P017nsss(0) <='0';
          end if;
        if(cVar1S16S108P064P012N030P054(0)='1' AND  E( 2)='0' )then
          cVar2S16S108P060nsss(0) <='1';
          else
          cVar2S16S108P060nsss(0) <='0';
          end if;
        if(cVar1S17S108P064P012N030P054(0)='1' AND  E( 2)='1' AND D(10)='0' AND B( 2)='1' )then
          cVar2S17S108P060P059P033nsss(0) <='1';
          else
          cVar2S17S108P060P059P033nsss(0) <='0';
          end if;
        if(cVar1S18S108P064P012N030N054(0)='1' AND  E( 2)='1' AND A(17)='0' AND E( 3)='0' )then
          cVar2S18S108P060P004P056nsss(0) <='1';
          else
          cVar2S18S108P060P004P056nsss(0) <='0';
          end if;
        if(cVar1S19S108P064P012N030N054(0)='1' AND  E( 2)='0' AND E( 0)='1' AND A(10)='1' )then
          cVar2S19S108N060P068P018nsss(0) <='1';
          else
          cVar2S19S108N060P068P018nsss(0) <='0';
          end if;
        if(cVar1S20S108P064P068P062P066(0)='1' AND  E(10)='1' )then
          cVar2S20S108P061nsss(0) <='1';
          else
          cVar2S20S108P061nsss(0) <='0';
          end if;
        if(cVar1S21S108P064P068P062P066(0)='1' AND  E(10)='0' AND A(12)='0' AND A( 7)='0' )then
          cVar2S21S108N061P014P005nsss(0) <='1';
          else
          cVar2S21S108N061P014P005nsss(0) <='0';
          end if;
        if(cVar1S22S108P064P068P062P066(0)='1' AND  E(10)='0' AND A(12)='1' AND A( 3)='1' )then
          cVar2S22S108N061P014P013nsss(0) <='1';
          else
          cVar2S22S108N061P014P013nsss(0) <='0';
          end if;
        if(cVar1S23S108P064P068P062N066(0)='1' AND  E( 8)='1' AND B(10)='1' )then
          cVar2S23S108P069P034nsss(0) <='1';
          else
          cVar2S23S108P069P034nsss(0) <='0';
          end if;
        if(cVar1S24S108P064P068P062N066(0)='1' AND  E( 8)='1' AND B(10)='0' AND A( 0)='1' )then
          cVar2S24S108P069N034P019nsss(0) <='1';
          else
          cVar2S24S108P069N034P019nsss(0) <='0';
          end if;
        if(cVar1S25S108P064P068P062N066(0)='1' AND  E( 8)='0' AND D( 9)='1' AND A(12)='1' )then
          cVar2S25S108N069P063P014nsss(0) <='1';
          else
          cVar2S25S108N069P063P014nsss(0) <='0';
          end if;
        if(cVar1S26S108P064P068P062P045(0)='1' AND  A(11)='1' )then
          cVar2S26S108P016nsss(0) <='1';
          else
          cVar2S26S108P016nsss(0) <='0';
          end if;
        if(cVar1S27S108P064P068P062P045(0)='1' AND  A(11)='0' AND A( 2)='0' AND B(16)='1' )then
          cVar2S27S108N016P015P022nsss(0) <='1';
          else
          cVar2S27S108N016P015P022nsss(0) <='0';
          end if;
        if(cVar1S28S108P064P068P062N045(0)='1' AND  D(14)='0' AND A(15)='1' )then
          cVar2S28S108P043P008nsss(0) <='1';
          else
          cVar2S28S108P043P008nsss(0) <='0';
          end if;
        if(cVar1S29S108P064P068P062N045(0)='1' AND  D(14)='0' AND A(15)='0' AND B( 6)='1' )then
          cVar2S29S108P043N008P025nsss(0) <='1';
          else
          cVar2S29S108P043N008P025nsss(0) <='0';
          end if;
        if(cVar1S30S108P064P068P012P035(0)='1' AND  E( 9)='1' )then
          cVar2S30S108P065nsss(0) <='1';
          else
          cVar2S30S108P065nsss(0) <='0';
          end if;
        if(cVar1S31S108P064P068P012P035(0)='1' AND  E( 9)='0' AND A(10)='1' )then
          cVar2S31S108N065P018nsss(0) <='1';
          else
          cVar2S31S108N065P018nsss(0) <='0';
          end if;
        if(cVar1S32S108P064P068P012P035(0)='1' AND  E( 9)='0' AND A(10)='0' AND A( 4)='0' )then
          cVar2S32S108N065N018P011nsss(0) <='1';
          else
          cVar2S32S108N065N018P011nsss(0) <='0';
          end if;
        if(cVar1S33S108P064P068P012N035(0)='1' AND  E(11)='1' )then
          cVar2S33S108P057nsss(0) <='1';
          else
          cVar2S33S108P057nsss(0) <='0';
          end if;
        if(cVar1S34S108P064P068P012N035(0)='1' AND  E(11)='0' AND A( 3)='0' AND D( 0)='1' )then
          cVar2S34S108N057P013P066nsss(0) <='1';
          else
          cVar2S34S108N057P013P066nsss(0) <='0';
          end if;
        if(cVar1S35S108P064P068N012P019(0)='1' AND  B(12)='1' )then
          cVar2S35S108P030nsss(0) <='1';
          else
          cVar2S35S108P030nsss(0) <='0';
          end if;
        if(cVar1S36S108P064P068N012P019(0)='1' AND  B(12)='0' AND D(12)='0' AND A(16)='1' )then
          cVar2S36S108N030P051P006nsss(0) <='1';
          else
          cVar2S36S108N030P051P006nsss(0) <='0';
          end if;
        if(cVar1S37S108P064P068N012N019(0)='1' AND  A( 1)='1' AND A( 5)='1' )then
          cVar2S37S108P017P009nsss(0) <='1';
          else
          cVar2S37S108P017P009nsss(0) <='0';
          end if;
        if(cVar1S38S108P064P068N012N019(0)='1' AND  A( 1)='1' AND A( 5)='0' AND A(15)='1' )then
          cVar2S38S108P017N009P008nsss(0) <='1';
          else
          cVar2S38S108P017N009P008nsss(0) <='0';
          end if;
        if(cVar1S39S108P064P068N012N019(0)='1' AND  A( 1)='0' AND A( 2)='1' AND A( 4)='1' )then
          cVar2S39S108N017P015P011nsss(0) <='1';
          else
          cVar2S39S108N017P015P011nsss(0) <='0';
          end if;
        if(cVar1S0S109P064P068P055P056(0)='1' AND  E(11)='1' AND A(12)='1' )then
          cVar2S0S109P057P014nsss(0) <='1';
          else
          cVar2S0S109P057P014nsss(0) <='0';
          end if;
        if(cVar1S1S109P064P068P055P056(0)='1' AND  E(11)='1' AND A(12)='0' AND A(10)='1' )then
          cVar2S1S109P057N014P018nsss(0) <='1';
          else
          cVar2S1S109P057N014P018nsss(0) <='0';
          end if;
        if(cVar1S2S109P064P068P055P056(0)='1' AND  E(11)='0' AND E( 5)='0' )then
          cVar2S2S109N057P048nsss(0) <='1';
          else
          cVar2S2S109N057P048nsss(0) <='0';
          end if;
        if(cVar1S3S109P064P068P055P056(0)='1' AND  E(11)='0' AND E( 5)='1' AND B( 6)='1' )then
          cVar2S3S109N057P048P025nsss(0) <='1';
          else
          cVar2S3S109N057P048P025nsss(0) <='0';
          end if;
        if(cVar1S4S109P064P068P055P056(0)='1' AND  E( 4)='0' AND D( 8)='1' AND B( 1)='1' )then
          cVar2S4S109P052P067P035nsss(0) <='1';
          else
          cVar2S4S109P052P067P035nsss(0) <='0';
          end if;
        if(cVar1S5S109P064P068P055P060(0)='1' AND  B( 3)='1' AND A( 3)='1' )then
          cVar2S5S109P031P013nsss(0) <='1';
          else
          cVar2S5S109P031P013nsss(0) <='0';
          end if;
        if(cVar1S6S109P064P068P055P060(0)='1' AND  B( 3)='0' AND B( 4)='1' )then
          cVar2S6S109N031P029nsss(0) <='1';
          else
          cVar2S6S109N031P029nsss(0) <='0';
          end if;
        if(cVar1S7S109P064P068P055P060(0)='1' AND  B( 3)='0' AND B( 4)='0' AND A( 2)='1' )then
          cVar2S7S109N031N029P015nsss(0) <='1';
          else
          cVar2S7S109N031N029P015nsss(0) <='0';
          end if;
        if(cVar1S8S109P064P068P051P019(0)='1' AND  D(13)='0' )then
          cVar2S8S109P047nsss(0) <='1';
          else
          cVar2S8S109P047nsss(0) <='0';
          end if;
        if(cVar1S9S109P064P068P051N019(0)='1' AND  A( 5)='1' AND D( 9)='1' )then
          cVar2S9S109P009P063nsss(0) <='1';
          else
          cVar2S9S109P009P063nsss(0) <='0';
          end if;
        if(cVar1S10S109P064P068P051N019(0)='1' AND  A( 5)='1' AND D( 9)='0' AND D( 8)='1' )then
          cVar2S10S109P009N063P067nsss(0) <='1';
          else
          cVar2S10S109P009N063P067nsss(0) <='0';
          end if;
        if(cVar1S11S109P064P068P051N019(0)='1' AND  A( 5)='0' AND B( 9)='0' AND B( 0)='0' )then
          cVar2S11S109N009P036P037nsss(0) <='1';
          else
          cVar2S11S109N009P036P037nsss(0) <='0';
          end if;
        if(cVar1S13S109N064P054P040P015(0)='1' AND  A( 3)='1' AND D( 2)='1' )then
          cVar2S13S109P013P058nsss(0) <='1';
          else
          cVar2S13S109P013P058nsss(0) <='0';
          end if;
        if(cVar1S14S109N064P054P040P015(0)='1' AND  A( 3)='1' AND D( 2)='0' AND A(10)='0' )then
          cVar2S14S109P013N058P018nsss(0) <='1';
          else
          cVar2S14S109P013N058P018nsss(0) <='0';
          end if;
        if(cVar1S15S109N064P054P040P015(0)='1' AND  A( 3)='0' AND E( 4)='1' AND A(11)='0' )then
          cVar2S15S109N013P052P016nsss(0) <='1';
          else
          cVar2S15S109N013P052P016nsss(0) <='0';
          end if;
        if(cVar1S16S109N064P054P040P015(0)='1' AND  A( 3)='0' AND E( 4)='0' AND B(12)='1' )then
          cVar2S16S109N013N052P030nsss(0) <='1';
          else
          cVar2S16S109N013N052P030nsss(0) <='0';
          end if;
        if(cVar1S17S109N064P054P040N015(0)='1' AND  A(15)='1' AND A( 4)='0' )then
          cVar2S17S109P008P011nsss(0) <='1';
          else
          cVar2S17S109P008P011nsss(0) <='0';
          end if;
        if(cVar1S18S109N064P054P040N015(0)='1' AND  A(15)='1' AND A( 4)='1' AND E( 3)='0' )then
          cVar2S18S109P008P011P056nsss(0) <='1';
          else
          cVar2S18S109P008P011P056nsss(0) <='0';
          end if;
        if(cVar1S19S109N064P054P040N015(0)='1' AND  A(15)='0' AND A( 5)='1' )then
          cVar2S19S109N008P009nsss(0) <='1';
          else
          cVar2S19S109N008P009nsss(0) <='0';
          end if;
        if(cVar1S20S109N064N054P022P043(0)='1' AND  A( 8)='1' )then
          cVar2S20S109P003nsss(0) <='1';
          else
          cVar2S20S109P003nsss(0) <='0';
          end if;
        if(cVar1S21S109N064N054P022P043(0)='1' AND  A( 8)='0' AND A( 6)='1' )then
          cVar2S21S109N003P007nsss(0) <='1';
          else
          cVar2S21S109N003P007nsss(0) <='0';
          end if;
        if(cVar1S22S109N064N054P022P043(0)='1' AND  A( 8)='0' AND A( 6)='0' AND E(14)='0' )then
          cVar2S22S109N003N007P045nsss(0) <='1';
          else
          cVar2S22S109N003N007P045nsss(0) <='0';
          end if;
        if(cVar1S23S109N064N054P022N043(0)='1' AND  D( 6)='1' AND A(17)='1' )then
          cVar2S23S109P042P004nsss(0) <='1';
          else
          cVar2S23S109P042P004nsss(0) <='0';
          end if;
        if(cVar1S24S109N064N054P022N043(0)='1' AND  D( 6)='1' AND A(17)='0' AND A(16)='1' )then
          cVar2S24S109P042N004P006nsss(0) <='1';
          else
          cVar2S24S109P042N004P006nsss(0) <='0';
          end if;
        if(cVar1S25S109N064N054P022N043(0)='1' AND  D( 6)='0' AND A(16)='0' AND E( 4)='1' )then
          cVar2S25S109N042P006P052nsss(0) <='1';
          else
          cVar2S25S109N042P006P052nsss(0) <='0';
          end if;
        if(cVar1S26S109N064N054N022P043(0)='1' AND  D(13)='1' AND B(15)='1' AND B(14)='0' )then
          cVar2S26S109P047P024P026nsss(0) <='1';
          else
          cVar2S26S109P047P024P026nsss(0) <='0';
          end if;
        if(cVar1S27S109N064N054N022P043(0)='1' AND  D(13)='1' AND B(15)='0' AND B(14)='1' )then
          cVar2S27S109P047N024P026nsss(0) <='1';
          else
          cVar2S27S109P047N024P026nsss(0) <='0';
          end if;
        if(cVar1S28S109N064N054N022P043(0)='1' AND  D(13)='0' AND B(15)='1' AND A( 7)='1' )then
          cVar2S28S109N047P024P005nsss(0) <='1';
          else
          cVar2S28S109N047P024P005nsss(0) <='0';
          end if;
        if(cVar1S29S109N064N054N022P043(0)='1' AND  D(13)='0' AND A(16)='1' )then
          cVar2S29S109P047P006nsss(0) <='1';
          else
          cVar2S29S109P047P006nsss(0) <='0';
          end if;
        if(cVar1S0S110P064P056P052P027(0)='1' AND  D( 4)='0' AND D( 6)='0' )then
          cVar2S0S110P050P042nsss(0) <='1';
          else
          cVar2S0S110P050P042nsss(0) <='0';
          end if;
        if(cVar1S1S110P064P056P052P027(0)='1' AND  D( 4)='1' AND D( 2)='1' )then
          cVar2S1S110P050P058nsss(0) <='1';
          else
          cVar2S1S110P050P058nsss(0) <='0';
          end if;
        if(cVar1S2S110P064P056P052P027(0)='1' AND  B( 3)='1' )then
          cVar2S2S110P031nsss(0) <='1';
          else
          cVar2S2S110P031nsss(0) <='0';
          end if;
        if(cVar1S4S110P064P056P052N009(0)='1' AND  A( 2)='1' )then
          cVar2S4S110P015nsss(0) <='1';
          else
          cVar2S4S110P015nsss(0) <='0';
          end if;
        if(cVar1S5S110P064P056P052N009(0)='1' AND  A( 2)='0' AND B( 4)='0' AND D( 4)='0' )then
          cVar2S5S110N015P029P050nsss(0) <='1';
          else
          cVar2S5S110N015P029P050nsss(0) <='0';
          end if;
        if(cVar1S6S110P064N056P026P049(0)='1' AND  A(11)='1' AND E( 9)='1' )then
          cVar2S6S110P016P065nsss(0) <='1';
          else
          cVar2S6S110P016P065nsss(0) <='0';
          end if;
        if(cVar1S7S110P064N056P026P049(0)='1' AND  A(11)='1' AND E( 9)='0' AND E( 0)='1' )then
          cVar2S7S110P016N065P068nsss(0) <='1';
          else
          cVar2S7S110P016N065P068nsss(0) <='0';
          end if;
        if(cVar1S8S110P064N056P026P049(0)='1' AND  A(11)='0' AND D( 9)='0' AND B(10)='0' )then
          cVar2S8S110N016P063P034nsss(0) <='1';
          else
          cVar2S8S110N016P063P034nsss(0) <='0';
          end if;
        if(cVar1S9S110P064N056P026P049(0)='1' AND  A(11)='0' AND D( 9)='1' AND B(10)='1' )then
          cVar2S9S110N016P063P034nsss(0) <='1';
          else
          cVar2S9S110N016P063P034nsss(0) <='0';
          end if;
        if(cVar1S10S110P064N056P026P049(0)='1' AND  B(15)='1' AND E(14)='0' )then
          cVar2S10S110P024P045nsss(0) <='1';
          else
          cVar2S10S110P024P045nsss(0) <='0';
          end if;
        if(cVar1S11S110P064N056P026P049(0)='1' AND  B(15)='0' AND B( 5)='1' )then
          cVar2S11S110N024P027nsss(0) <='1';
          else
          cVar2S11S110N024P027nsss(0) <='0';
          end if;
        if(cVar1S12S110P064N056P026P049(0)='1' AND  B(15)='0' AND B( 5)='0' AND B( 2)='1' )then
          cVar2S12S110N024N027P033nsss(0) <='1';
          else
          cVar2S12S110N024N027P033nsss(0) <='0';
          end if;
        if(cVar1S13S110P064N056P026P050(0)='1' AND  B( 9)='1' )then
          cVar2S13S110P036nsss(0) <='1';
          else
          cVar2S13S110P036nsss(0) <='0';
          end if;
        if(cVar1S14S110P064N056P026P050(0)='1' AND  B( 9)='0' AND A(11)='0' )then
          cVar2S14S110N036P016nsss(0) <='1';
          else
          cVar2S14S110N036P016nsss(0) <='0';
          end if;
        if(cVar1S15S110P064N056P026P050(0)='1' AND  B( 9)='0' AND A(11)='1' AND A( 0)='1' )then
          cVar2S15S110N036P016P019nsss(0) <='1';
          else
          cVar2S15S110N036P016P019nsss(0) <='0';
          end if;
        if(cVar1S16S110P064N056P026N050(0)='1' AND  D(12)='1' AND A( 0)='1' )then
          cVar2S16S110P051P019nsss(0) <='1';
          else
          cVar2S16S110P051P019nsss(0) <='0';
          end if;
        if(cVar1S17S110P064N056P026N050(0)='1' AND  D(12)='1' AND A( 0)='0' AND E( 8)='0' )then
          cVar2S17S110P051N019P069nsss(0) <='1';
          else
          cVar2S17S110P051N019P069nsss(0) <='0';
          end if;
        if(cVar1S18S110P064N056P026N050(0)='1' AND  D(12)='0' AND D( 5)='1' AND A(14)='1' )then
          cVar2S18S110N051P046P010nsss(0) <='1';
          else
          cVar2S18S110N051P046P010nsss(0) <='0';
          end if;
        if(cVar1S19S110P064P013P047P026(0)='1' AND  A( 0)='0' AND B(13)='1' AND A(14)='0' )then
          cVar2S19S110P019P028P010nsss(0) <='1';
          else
          cVar2S19S110P019P028P010nsss(0) <='0';
          end if;
        if(cVar1S20S110P064P013P047P026(0)='1' AND  A( 0)='0' AND B(13)='0' )then
          cVar2S20S110P019N028psss(0) <='1';
          else
          cVar2S20S110P019N028psss(0) <='0';
          end if;
        if(cVar1S21S110P064P013P047P026(0)='1' AND  A( 0)='1' AND E( 0)='1' AND B( 0)='1' )then
          cVar2S21S110P019P068P037nsss(0) <='1';
          else
          cVar2S21S110P019P068P037nsss(0) <='0';
          end if;
        if(cVar1S22S110P064P013P047P026(0)='1' AND  A( 0)='1' AND E( 0)='0' AND D( 9)='1' )then
          cVar2S22S110P019N068P063nsss(0) <='1';
          else
          cVar2S22S110P019N068P063nsss(0) <='0';
          end if;
        if(cVar1S23S110P064P013P047P026(0)='1' AND  A( 5)='0' AND A(11)='1' )then
          cVar2S23S110P009P016nsss(0) <='1';
          else
          cVar2S23S110P009P016nsss(0) <='0';
          end if;
        if(cVar1S24S110P064N013P033P022(0)='1' AND  B( 7)='1' )then
          cVar2S24S110P023nsss(0) <='1';
          else
          cVar2S24S110P023nsss(0) <='0';
          end if;
        if(cVar1S25S110P064N013P033P022(0)='1' AND  B( 9)='0' AND A( 2)='0' AND A(11)='0' )then
          cVar2S25S110P036P015P016nsss(0) <='1';
          else
          cVar2S25S110P036P015P016nsss(0) <='0';
          end if;
        if(cVar1S26S110P064N013P033P050(0)='1' AND  B(10)='1' )then
          cVar2S26S110P034nsss(0) <='1';
          else
          cVar2S26S110P034nsss(0) <='0';
          end if;
        if(cVar1S27S110P064N013P033P050(0)='1' AND  B(10)='0' AND E( 5)='0' AND A(19)='1' )then
          cVar2S27S110N034P048P000nsss(0) <='1';
          else
          cVar2S27S110N034P048P000nsss(0) <='0';
          end if;
        if(cVar1S0S111P064P033P041P018(0)='1' AND  A( 2)='1' AND E(14)='0' )then
          cVar2S0S111P015P045nsss(0) <='1';
          else
          cVar2S0S111P015P045nsss(0) <='0';
          end if;
        if(cVar1S1S111P064P033P041P018(0)='1' AND  A( 2)='0' AND D( 2)='0' )then
          cVar2S1S111N015P058nsss(0) <='1';
          else
          cVar2S1S111N015P058nsss(0) <='0';
          end if;
        if(cVar1S2S111P064P033P041P018(0)='1' AND  A( 2)='0' AND D( 2)='1' AND B(11)='1' )then
          cVar2S2S111N015P058P032nsss(0) <='1';
          else
          cVar2S2S111N015P058P032nsss(0) <='0';
          end if;
        if(cVar1S3S111P064P033P041P018(0)='1' AND  E( 9)='1' )then
          cVar2S3S111P065nsss(0) <='1';
          else
          cVar2S3S111P065nsss(0) <='0';
          end if;
        if(cVar1S4S111P064P033P041P018(0)='1' AND  E( 9)='0' AND A( 4)='1' AND A( 2)='0' )then
          cVar2S4S111N065P011P015nsss(0) <='1';
          else
          cVar2S4S111N065P011P015nsss(0) <='0';
          end if;
        if(cVar1S6S111P064P033P048P050(0)='1' AND  B(10)='1' AND A( 8)='0' )then
          cVar2S6S111P034P003nsss(0) <='1';
          else
          cVar2S6S111P034P003nsss(0) <='0';
          end if;
        if(cVar1S7S111P064P033P048P050(0)='1' AND  B(10)='0' AND A( 8)='1' AND A( 0)='1' )then
          cVar2S7S111N034P003P019nsss(0) <='1';
          else
          cVar2S7S111N034P003P019nsss(0) <='0';
          end if;
        if(cVar1S8S111P064P033P048P050(0)='1' AND  B(10)='0' AND A( 8)='0' AND A(12)='0' )then
          cVar2S8S111N034N003P014nsss(0) <='1';
          else
          cVar2S8S111N034N003P014nsss(0) <='0';
          end if;
        if(cVar1S9S111N064P016P047P024(0)='1' AND  B(17)='0' AND E(11)='1' )then
          cVar2S9S111P020P057nsss(0) <='1';
          else
          cVar2S9S111P020P057nsss(0) <='0';
          end if;
        if(cVar1S10S111N064P016P047P024(0)='1' AND  B(17)='0' AND E(11)='0' AND A(19)='0' )then
          cVar2S10S111P020N057P000nsss(0) <='1';
          else
          cVar2S10S111P020N057P000nsss(0) <='0';
          end if;
        if(cVar1S11S111N064P016P047P024(0)='1' AND  B(17)='1' AND A( 2)='0' AND A(14)='0' )then
          cVar2S11S111P020P015P010nsss(0) <='1';
          else
          cVar2S11S111P020P015P010nsss(0) <='0';
          end if;
        if(cVar1S12S111N064P016P047P024(0)='1' AND  B(17)='1' AND A( 2)='1' AND A(13)='1' )then
          cVar2S12S111P020P015P012nsss(0) <='1';
          else
          cVar2S12S111P020P015P012nsss(0) <='0';
          end if;
        if(cVar1S13S111N064P016P047P024(0)='1' AND  A(16)='1' AND E( 0)='0' )then
          cVar2S13S111P006P068nsss(0) <='1';
          else
          cVar2S13S111P006P068nsss(0) <='0';
          end if;
        if(cVar1S14S111N064P016P047P024(0)='1' AND  A(16)='0' AND A( 9)='0' AND E( 8)='1' )then
          cVar2S14S111N006P001P069nsss(0) <='1';
          else
          cVar2S14S111N006P001P069nsss(0) <='0';
          end if;
        if(cVar1S15S111N064P016P047P034(0)='1' AND  A( 4)='0' )then
          cVar2S15S111P011nsss(0) <='1';
          else
          cVar2S15S111P011nsss(0) <='0';
          end if;
        if(cVar1S16S111N064P016P047N034(0)='1' AND  E( 9)='0' AND A(10)='1' AND E( 0)='0' )then
          cVar2S16S111P065P018P068nsss(0) <='1';
          else
          cVar2S16S111P065P018P068nsss(0) <='0';
          end if;
        if(cVar1S17S111N064P016P047N034(0)='1' AND  E( 9)='0' AND A(10)='0' AND A( 2)='1' )then
          cVar2S17S111P065N018P015nsss(0) <='1';
          else
          cVar2S17S111P065N018P015nsss(0) <='0';
          end if;
        if(cVar1S18S111N064N016P018P015(0)='1' AND  E(13)='1' AND D( 8)='1' )then
          cVar2S18S111P049P067nsss(0) <='1';
          else
          cVar2S18S111P049P067nsss(0) <='0';
          end if;
        if(cVar1S19S111N064N016P018P015(0)='1' AND  E(13)='1' AND D( 8)='0' AND A( 1)='1' )then
          cVar2S19S111P049N067P017nsss(0) <='1';
          else
          cVar2S19S111P049N067P017nsss(0) <='0';
          end if;
        if(cVar1S20S111N064N016P018P015(0)='1' AND  E(13)='0' AND A( 1)='1' AND E( 0)='1' )then
          cVar2S20S111N049P017P068nsss(0) <='1';
          else
          cVar2S20S111N049P017P068nsss(0) <='0';
          end if;
        if(cVar1S21S111N064N016P018P015(0)='1' AND  E(13)='0' AND A( 1)='0' AND A( 8)='1' )then
          cVar2S21S111N049N017P003nsss(0) <='1';
          else
          cVar2S21S111N049N017P003nsss(0) <='0';
          end if;
        if(cVar1S22S111N064N016P018N015(0)='1' AND  A(17)='1' AND A( 1)='1' )then
          cVar2S22S111P004P017nsss(0) <='1';
          else
          cVar2S22S111P004P017nsss(0) <='0';
          end if;
        if(cVar1S23S111N064N016P018N015(0)='1' AND  A(17)='1' AND A( 1)='0' AND A(18)='0' )then
          cVar2S23S111P004N017P002nsss(0) <='1';
          else
          cVar2S23S111P004N017P002nsss(0) <='0';
          end if;
        if(cVar1S24S111N064N016P018N015(0)='1' AND  A(17)='0' AND A(15)='1' )then
          cVar2S24S111N004P008nsss(0) <='1';
          else
          cVar2S24S111N004P008nsss(0) <='0';
          end if;
        if(cVar1S25S111N064N016N018P059(0)='1' AND  D( 6)='0' AND E(12)='0' )then
          cVar2S25S111P042P053nsss(0) <='1';
          else
          cVar2S25S111P042P053nsss(0) <='0';
          end if;
        if(cVar1S26S111N064N016N018N059(0)='1' AND  E(10)='0' AND A(12)='1' AND A(13)='0' )then
          cVar2S26S111P061P014P012nsss(0) <='1';
          else
          cVar2S26S111P061P014P012nsss(0) <='0';
          end if;
        if(cVar1S27S111N064N016N018N059(0)='1' AND  E(10)='1' AND E( 4)='1' )then
          cVar2S27S111P061P052nsss(0) <='1';
          else
          cVar2S27S111P061P052nsss(0) <='0';
          end if;
        if(cVar1S0S112P018P016P027P066(0)='1' AND  A( 5)='0' AND B( 2)='0' AND E( 3)='0' )then
          cVar2S0S112P009P033P056nsss(0) <='1';
          else
          cVar2S0S112P009P033P056nsss(0) <='0';
          end if;
        if(cVar1S1S112P018P016P027P066(0)='1' AND  A( 5)='0' AND B( 2)='1' AND E(10)='1' )then
          cVar2S1S112P009P033P061nsss(0) <='1';
          else
          cVar2S1S112P009P033P061nsss(0) <='0';
          end if;
        if(cVar1S2S112P018P016P027P066(0)='1' AND  A( 5)='1' AND E( 9)='1' AND A( 3)='0' )then
          cVar2S2S112P009P065P013nsss(0) <='1';
          else
          cVar2S2S112P009P065P013nsss(0) <='0';
          end if;
        if(cVar1S3S112P018P016P027P066(0)='1' AND  A( 5)='1' AND E( 9)='0' AND B(11)='1' )then
          cVar2S3S112P009N065P032nsss(0) <='1';
          else
          cVar2S3S112P009N065P032nsss(0) <='0';
          end if;
        if(cVar1S4S112P018P016P027P066(0)='1' AND  A(13)='1' AND A( 5)='1' )then
          cVar2S4S112P012P009nsss(0) <='1';
          else
          cVar2S4S112P012P009nsss(0) <='0';
          end if;
        if(cVar1S5S112P018P016P027P066(0)='1' AND  A(13)='1' AND A( 5)='0' AND A( 1)='0' )then
          cVar2S5S112P012N009P017nsss(0) <='1';
          else
          cVar2S5S112P012N009P017nsss(0) <='0';
          end if;
        if(cVar1S6S112P018P016P027P066(0)='1' AND  A(13)='0' AND E( 8)='0' )then
          cVar2S6S112N012P069nsss(0) <='1';
          else
          cVar2S6S112N012P069nsss(0) <='0';
          end if;
        if(cVar1S7S112P018P016P027P066(0)='1' AND  A(13)='0' AND E( 8)='1' AND B( 1)='1' )then
          cVar2S7S112N012P069P035nsss(0) <='1';
          else
          cVar2S7S112N012P069P035nsss(0) <='0';
          end if;
        if(cVar1S8S112P018P016P027P009(0)='1' AND  D( 0)='0' AND E(13)='1' )then
          cVar2S8S112P066P049nsss(0) <='1';
          else
          cVar2S8S112P066P049nsss(0) <='0';
          end if;
        if(cVar1S9S112P018P016P027P009(0)='1' AND  D( 0)='0' AND E(13)='0' AND E( 4)='0' )then
          cVar2S9S112P066N049P052nsss(0) <='1';
          else
          cVar2S9S112P066N049P052nsss(0) <='0';
          end if;
        if(cVar1S10S112P018P016P027P009(0)='1' AND  D( 0)='1' AND D( 4)='1' )then
          cVar2S10S112P066P050nsss(0) <='1';
          else
          cVar2S10S112P066P050nsss(0) <='0';
          end if;
        if(cVar1S11S112P018P016P027N009(0)='1' AND  D( 9)='1' )then
          cVar2S11S112P063nsss(0) <='1';
          else
          cVar2S11S112P063nsss(0) <='0';
          end if;
        if(cVar1S12S112P018P016P027N009(0)='1' AND  D( 9)='0' AND A( 2)='1' AND A( 1)='0' )then
          cVar2S12S112N063P015P017nsss(0) <='1';
          else
          cVar2S12S112N063P015P017nsss(0) <='0';
          end if;
        if(cVar1S13S112P018P016P027N009(0)='1' AND  D( 9)='0' AND A( 2)='0' AND E( 4)='1' )then
          cVar2S13S112N063N015P052nsss(0) <='1';
          else
          cVar2S13S112N063N015P052nsss(0) <='0';
          end if;
        if(cVar1S14S112P018P016P059P065(0)='1' AND  B(15)='0' AND A(17)='1' )then
          cVar2S14S112P024P004nsss(0) <='1';
          else
          cVar2S14S112P024P004nsss(0) <='0';
          end if;
        if(cVar1S15S112P018P016P059P065(0)='1' AND  B(15)='0' AND A(17)='0' AND A(16)='0' )then
          cVar2S15S112P024N004P006nsss(0) <='1';
          else
          cVar2S15S112P024N004P006nsss(0) <='0';
          end if;
        if(cVar1S16S112P018P016P059P065(0)='1' AND  E( 8)='0' AND E(10)='1' AND A( 0)='0' )then
          cVar2S16S112P069P061P019nsss(0) <='1';
          else
          cVar2S16S112P069P061P019nsss(0) <='0';
          end if;
        if(cVar1S17S112P018P016N059P066(0)='1' AND  E(10)='0' AND D( 9)='1' )then
          cVar2S17S112P061P063nsss(0) <='1';
          else
          cVar2S17S112P061P063nsss(0) <='0';
          end if;
        if(cVar1S18S112P018P016N059P066(0)='1' AND  E(10)='0' AND D( 9)='0' AND E( 3)='1' )then
          cVar2S18S112P061N063P056nsss(0) <='1';
          else
          cVar2S18S112P061N063P056nsss(0) <='0';
          end if;
        if(cVar1S19S112P018P016N059P066(0)='1' AND  E(10)='1' AND A( 0)='1' AND A( 2)='1' )then
          cVar2S19S112P061P019P015nsss(0) <='1';
          else
          cVar2S19S112P061P019P015nsss(0) <='0';
          end if;
        if(cVar1S20S112P018P016N059P066(0)='1' AND  D( 8)='1' AND D(12)='1' )then
          cVar2S20S112P067P051nsss(0) <='1';
          else
          cVar2S20S112P067P051nsss(0) <='0';
          end if;
        if(cVar1S21S112P018P016N059P066(0)='1' AND  D( 8)='1' AND D(12)='0' AND D( 9)='1' )then
          cVar2S21S112P067N051P063nsss(0) <='1';
          else
          cVar2S21S112P067N051P063nsss(0) <='0';
          end if;
        if(cVar1S22S112N018P054P040P065(0)='1' AND  B(15)='1' )then
          cVar2S22S112P024nsss(0) <='1';
          else
          cVar2S22S112P024nsss(0) <='0';
          end if;
        if(cVar1S23S112N018P054P040P065(0)='1' AND  B(15)='0' AND B( 1)='1' AND A( 5)='0' )then
          cVar2S23S112N024P035P009nsss(0) <='1';
          else
          cVar2S23S112N024P035P009nsss(0) <='0';
          end if;
        if(cVar1S24S112N018P054P040P065(0)='1' AND  B(15)='0' AND B( 1)='0' AND E( 3)='1' )then
          cVar2S24S112N024N035P056nsss(0) <='1';
          else
          cVar2S24S112N024N035P056nsss(0) <='0';
          end if;
        if(cVar1S25S112N018P054P040P065(0)='1' AND  B( 0)='1' )then
          cVar2S25S112P037nsss(0) <='1';
          else
          cVar2S25S112P037nsss(0) <='0';
          end if;
        if(cVar1S26S112N018P054P040P065(0)='1' AND  B( 0)='0' AND D( 9)='1' AND A(13)='1' )then
          cVar2S26S112N037P063P012nsss(0) <='1';
          else
          cVar2S26S112N037P063P012nsss(0) <='0';
          end if;
        if(cVar1S27S112N018N054P014P055(0)='1' AND  A( 3)='0' AND E(10)='0' AND E( 2)='0' )then
          cVar2S27S112P013P061P060nsss(0) <='1';
          else
          cVar2S27S112P013P061P060nsss(0) <='0';
          end if;
        if(cVar1S28S112N018N054P014P055(0)='1' AND  A( 3)='1' AND A( 8)='1' )then
          cVar2S28S112P013P003nsss(0) <='1';
          else
          cVar2S28S112P013P003nsss(0) <='0';
          end if;
        if(cVar1S29S112N018N054P014N055(0)='1' AND  E(11)='0' AND A( 4)='0' AND D( 7)='1' )then
          cVar2S29S112P057P011P038nsss(0) <='1';
          else
          cVar2S29S112P057P011P038nsss(0) <='0';
          end if;
        if(cVar1S30S112N018N054P014N055(0)='1' AND  E(11)='0' AND A( 4)='1' AND D( 4)='1' )then
          cVar2S30S112P057P011P050nsss(0) <='1';
          else
          cVar2S30S112P057P011P050nsss(0) <='0';
          end if;
        if(cVar1S31S112N018N054P014N055(0)='1' AND  E(11)='1' AND D(10)='1' AND B( 1)='1' )then
          cVar2S31S112P057P059P035nsss(0) <='1';
          else
          cVar2S31S112P057P059P035nsss(0) <='0';
          end if;
        if(cVar1S32S112N018N054P014N055(0)='1' AND  E(11)='1' AND D(10)='0' AND A( 8)='1' )then
          cVar2S32S112P057N059P003nsss(0) <='1';
          else
          cVar2S32S112P057N059P003nsss(0) <='0';
          end if;
        if(cVar1S33S112N018N054P014P031(0)='1' AND  A( 9)='1' AND D( 0)='0' )then
          cVar2S33S112P001P066nsss(0) <='1';
          else
          cVar2S33S112P001P066nsss(0) <='0';
          end if;
        if(cVar1S34S112N018N054P014P031(0)='1' AND  A( 9)='1' AND D( 0)='1' AND B( 0)='1' )then
          cVar2S34S112P001P066P037nsss(0) <='1';
          else
          cVar2S34S112P001P066P037nsss(0) <='0';
          end if;
        if(cVar1S35S112N018N054P014P031(0)='1' AND  A( 9)='0' AND E( 9)='1' AND E( 2)='0' )then
          cVar2S35S112N001P065P060nsss(0) <='1';
          else
          cVar2S35S112N001P065P060nsss(0) <='0';
          end if;
        if(cVar1S36S112N018N054P014P031(0)='1' AND  A( 9)='0' AND E( 9)='0' AND A( 2)='1' )then
          cVar2S36S112N001N065P015nsss(0) <='1';
          else
          cVar2S36S112N001N065P015nsss(0) <='0';
          end if;
        if(cVar1S37S112N018N054P014P031(0)='1' AND  D(11)='1' AND A( 4)='0' )then
          cVar2S37S112P055P011nsss(0) <='1';
          else
          cVar2S37S112P055P011nsss(0) <='0';
          end if;
        if(cVar1S0S113P014P018P056P011(0)='1' AND  E(11)='0' AND D(11)='0' )then
          cVar2S0S113P057P055nsss(0) <='1';
          else
          cVar2S0S113P057P055nsss(0) <='0';
          end if;
        if(cVar1S1S113P014P018P056P011(0)='1' AND  E(11)='0' AND D(11)='1' AND D( 2)='0' )then
          cVar2S1S113P057P055P058nsss(0) <='1';
          else
          cVar2S1S113P057P055P058nsss(0) <='0';
          end if;
        if(cVar1S2S113P014P018P056P011(0)='1' AND  E(11)='1' AND A(13)='1' )then
          cVar2S2S113P057P012nsss(0) <='1';
          else
          cVar2S2S113P057P012nsss(0) <='0';
          end if;
        if(cVar1S3S113P014P018P056P011(0)='1' AND  E(11)='1' AND A(13)='0' AND A( 8)='1' )then
          cVar2S3S113P057N012P003nsss(0) <='1';
          else
          cVar2S3S113P057N012P003nsss(0) <='0';
          end if;
        if(cVar1S4S113P014P018P056P011(0)='1' AND  D(11)='1' AND B( 4)='1' )then
          cVar2S4S113P055P029nsss(0) <='1';
          else
          cVar2S4S113P055P029nsss(0) <='0';
          end if;
        if(cVar1S5S113P014P018P056P011(0)='1' AND  D(11)='1' AND B( 4)='0' AND A(16)='0' )then
          cVar2S5S113P055N029P006nsss(0) <='1';
          else
          cVar2S5S113P055N029P006nsss(0) <='0';
          end if;
        if(cVar1S6S113P014P018P056P011(0)='1' AND  D(11)='0' AND A(15)='1' AND A( 6)='0' )then
          cVar2S6S113N055P008P007nsss(0) <='1';
          else
          cVar2S6S113N055P008P007nsss(0) <='0';
          end if;
        if(cVar1S7S113P014P018P056P011(0)='1' AND  D(11)='0' AND A(15)='0' AND A(16)='1' )then
          cVar2S7S113N055N008P006nsss(0) <='1';
          else
          cVar2S7S113N055N008P006nsss(0) <='0';
          end if;
        if(cVar1S8S113P014P018P056P017(0)='1' AND  E( 4)='0' AND A(11)='0' )then
          cVar2S8S113P052P016nsss(0) <='1';
          else
          cVar2S8S113P052P016nsss(0) <='0';
          end if;
        if(cVar1S9S113P014P018P056P017(0)='1' AND  E( 4)='0' AND A(11)='1' AND E( 1)='1' )then
          cVar2S9S113P052P016P064nsss(0) <='1';
          else
          cVar2S9S113P052P016P064nsss(0) <='0';
          end if;
        if(cVar1S10S113P014P018P056N017(0)='1' AND  E(11)='0' AND A( 3)='1' )then
          cVar2S10S113P057P013nsss(0) <='1';
          else
          cVar2S10S113P057P013nsss(0) <='0';
          end if;
        if(cVar1S11S113P014P018P056N017(0)='1' AND  E(11)='0' AND A( 3)='0' AND A( 5)='1' )then
          cVar2S11S113P057N013P009nsss(0) <='1';
          else
          cVar2S11S113P057N013P009nsss(0) <='0';
          end if;
        if(cVar1S12S113P014P018P056N017(0)='1' AND  E(11)='1' AND B( 3)='1' AND A( 3)='0' )then
          cVar2S12S113P057P031P013nsss(0) <='1';
          else
          cVar2S12S113P057P031P013nsss(0) <='0';
          end if;
        if(cVar1S13S113P014P018P067P050(0)='1' AND  B(12)='1' AND E( 3)='1' )then
          cVar2S13S113P030P056nsss(0) <='1';
          else
          cVar2S13S113P030P056nsss(0) <='0';
          end if;
        if(cVar1S14S113P014P018P067P050(0)='1' AND  B(12)='1' AND E( 3)='0' AND A(11)='1' )then
          cVar2S14S113P030N056P016nsss(0) <='1';
          else
          cVar2S14S113P030N056P016nsss(0) <='0';
          end if;
        if(cVar1S15S113P014P018P067P050(0)='1' AND  B(12)='0' AND D( 1)='0' AND A(11)='0' )then
          cVar2S15S113N030P062P016nsss(0) <='1';
          else
          cVar2S15S113N030P062P016nsss(0) <='0';
          end if;
        if(cVar1S16S113P014P018P067P050(0)='1' AND  B(12)='0' AND D( 1)='1' AND E( 0)='1' )then
          cVar2S16S113N030P062P068nsss(0) <='1';
          else
          cVar2S16S113N030P062P068nsss(0) <='0';
          end if;
        if(cVar1S17S113P014P018P067P050(0)='1' AND  A(13)='1' )then
          cVar2S17S113P012nsss(0) <='1';
          else
          cVar2S17S113P012nsss(0) <='0';
          end if;
        if(cVar1S18S113P014P018P067P050(0)='1' AND  A(13)='0' AND A(14)='1' )then
          cVar2S18S113N012P010nsss(0) <='1';
          else
          cVar2S18S113N012P010nsss(0) <='0';
          end if;
        if(cVar1S19S113P014P018P067P050(0)='1' AND  A(13)='0' AND A(14)='0' AND E( 0)='1' )then
          cVar2S19S113N012N010P068nsss(0) <='1';
          else
          cVar2S19S113N012N010P068nsss(0) <='0';
          end if;
        if(cVar1S20S113P014P018N067P012(0)='1' AND  E( 1)='1' AND B(11)='1' )then
          cVar2S20S113P064P032nsss(0) <='1';
          else
          cVar2S20S113P064P032nsss(0) <='0';
          end if;
        if(cVar1S21S113P014P018N067P012(0)='1' AND  E( 1)='1' AND B(11)='0' AND A( 3)='0' )then
          cVar2S21S113P064N032P013nsss(0) <='1';
          else
          cVar2S21S113P064N032P013nsss(0) <='0';
          end if;
        if(cVar1S22S113P014P018N067P012(0)='1' AND  E( 1)='0' AND B(10)='1' AND D( 2)='0' )then
          cVar2S22S113N064P034P058nsss(0) <='1';
          else
          cVar2S22S113N064P034P058nsss(0) <='0';
          end if;
        if(cVar1S23S113P014P018N067P012(0)='1' AND  E( 1)='0' AND B(10)='0' AND E( 0)='1' )then
          cVar2S23S113N064N034P068nsss(0) <='1';
          else
          cVar2S23S113N064N034P068nsss(0) <='0';
          end if;
        if(cVar1S24S113P014P018N067N012(0)='1' AND  A(11)='0' AND E( 4)='1' AND A(15)='1' )then
          cVar2S24S113P016P052P008nsss(0) <='1';
          else
          cVar2S24S113P016P052P008nsss(0) <='0';
          end if;
        if(cVar1S25S113P014P018N067N012(0)='1' AND  A(11)='0' AND E( 4)='0' AND B( 6)='1' )then
          cVar2S25S113P016N052P025nsss(0) <='1';
          else
          cVar2S25S113P016N052P025nsss(0) <='0';
          end if;
        if(cVar1S26S113P014P018N067N012(0)='1' AND  A(11)='1' AND B( 1)='1' AND E( 0)='0' )then
          cVar2S26S113P016P035P068nsss(0) <='1';
          else
          cVar2S26S113P016P035P068nsss(0) <='0';
          end if;
        if(cVar1S27S113P014P018N067N012(0)='1' AND  A(11)='1' AND B( 1)='0' AND A( 6)='1' )then
          cVar2S27S113P016N035P007nsss(0) <='1';
          else
          cVar2S27S113P016N035P007nsss(0) <='0';
          end if;
        if(cVar1S28S113P014P018P022P023(0)='1' AND  A(13)='0' )then
          cVar2S28S113P012nsss(0) <='1';
          else
          cVar2S28S113P012nsss(0) <='0';
          end if;
        if(cVar1S29S113P014P018P022N023(0)='1' AND  B( 0)='1' AND B(11)='1' AND A( 0)='0' )then
          cVar2S29S113P037P032P019nsss(0) <='1';
          else
          cVar2S29S113P037P032P019nsss(0) <='0';
          end if;
        if(cVar1S30S113P014P018P022N023(0)='1' AND  B( 0)='1' AND B(11)='0' AND B( 4)='0' )then
          cVar2S30S113P037N032P029nsss(0) <='1';
          else
          cVar2S30S113P037N032P029nsss(0) <='0';
          end if;
        if(cVar1S31S113P014P018P022N023(0)='1' AND  B( 0)='0' AND B( 2)='1' AND A( 0)='0' )then
          cVar2S31S113N037P033P019nsss(0) <='1';
          else
          cVar2S31S113N037P033P019nsss(0) <='0';
          end if;
        if(cVar1S32S113P014P018P022N023(0)='1' AND  B( 0)='0' AND B( 2)='0' AND B(12)='1' )then
          cVar2S32S113N037N033P030nsss(0) <='1';
          else
          cVar2S32S113N037N033P030nsss(0) <='0';
          end if;
        if(cVar1S34S113P014P018P022N037(0)='1' AND  D( 0)='0' AND A( 1)='1' )then
          cVar2S34S113P066P017nsss(0) <='1';
          else
          cVar2S34S113P066P017nsss(0) <='0';
          end if;
        if(cVar1S35S113P014N018P036P035(0)='1' AND  B(10)='0' AND E(10)='0' AND B( 7)='0' )then
          cVar2S35S113P034P061P023nsss(0) <='1';
          else
          cVar2S35S113P034P061P023nsss(0) <='0';
          end if;
        if(cVar1S36S113P014N018P036P035(0)='1' AND  B(10)='0' AND E(10)='1' AND A(11)='1' )then
          cVar2S36S113P034P061P016nsss(0) <='1';
          else
          cVar2S36S113P034P061P016nsss(0) <='0';
          end if;
        if(cVar1S37S113P014N018P036P035(0)='1' AND  B(10)='1' AND A(11)='1' AND D( 9)='1' )then
          cVar2S37S113P034P016P063nsss(0) <='1';
          else
          cVar2S37S113P034P016P063nsss(0) <='0';
          end if;
        if(cVar1S38S113P014N018P036P035(0)='1' AND  B(10)='1' AND A(11)='0' AND D( 9)='0' )then
          cVar2S38S113P034N016P063nsss(0) <='1';
          else
          cVar2S38S113P034N016P063nsss(0) <='0';
          end if;
        if(cVar1S39S113P014N018P036N035(0)='1' AND  E( 1)='0' AND A( 6)='0' AND A(15)='1' )then
          cVar2S39S113P064P007P008nsss(0) <='1';
          else
          cVar2S39S113P064P007P008nsss(0) <='0';
          end if;
        if(cVar1S40S113P014N018P036N035(0)='1' AND  E( 1)='0' AND A( 6)='1' AND D(11)='1' )then
          cVar2S40S113P064P007P055nsss(0) <='1';
          else
          cVar2S40S113P064P007P055nsss(0) <='0';
          end if;
        if(cVar1S41S113P014N018P036N035(0)='1' AND  E( 1)='1' AND E( 0)='1' AND A( 0)='1' )then
          cVar2S41S113P064P068P019nsss(0) <='1';
          else
          cVar2S41S113P064P068P019nsss(0) <='0';
          end if;
        if(cVar1S42S113P014N018P036N035(0)='1' AND  E( 1)='1' AND E( 0)='0' AND B(15)='1' )then
          cVar2S42S113P064N068P024nsss(0) <='1';
          else
          cVar2S42S113P064N068P024nsss(0) <='0';
          end if;
        if(cVar1S43S113P014N018P036P053(0)='1' AND  B(12)='0' AND A(15)='0' AND A(13)='1' )then
          cVar2S43S113P030P008P012nsss(0) <='1';
          else
          cVar2S43S113P030P008P012nsss(0) <='0';
          end if;
        if(cVar1S44S113P014N018P036P053(0)='1' AND  B(12)='1' AND A(13)='1' )then
          cVar2S44S113P030P012nsss(0) <='1';
          else
          cVar2S44S113P030P012nsss(0) <='0';
          end if;
        if(cVar1S0S114P018P064P007P032(0)='1' AND  B( 2)='0' )then
          cVar2S0S114P033nsss(0) <='1';
          else
          cVar2S0S114P033nsss(0) <='0';
          end if;
        if(cVar1S1S114P018P064P007N032(0)='1' AND  E(13)='1' AND A( 5)='1' )then
          cVar2S1S114P049P009nsss(0) <='1';
          else
          cVar2S1S114P049P009nsss(0) <='0';
          end if;
        if(cVar1S2S114P018P064P007N032(0)='1' AND  E(13)='1' AND A( 5)='0' AND B( 1)='1' )then
          cVar2S2S114P049N009P035nsss(0) <='1';
          else
          cVar2S2S114P049N009P035nsss(0) <='0';
          end if;
        if(cVar1S3S114P018P064P007N032(0)='1' AND  E(13)='0' AND E( 2)='0' )then
          cVar2S3S114N049P060nsss(0) <='1';
          else
          cVar2S3S114N049P060nsss(0) <='0';
          end if;
        if(cVar1S4S114P018P064P007N032(0)='1' AND  E(13)='0' AND E( 2)='1' AND B( 2)='1' )then
          cVar2S4S114N049P060P033nsss(0) <='1';
          else
          cVar2S4S114N049P060P033nsss(0) <='0';
          end if;
        if(cVar1S5S114P018P064P007P059(0)='1' AND  A( 3)='0' AND A( 8)='1' )then
          cVar2S5S114P013P003nsss(0) <='1';
          else
          cVar2S5S114P013P003nsss(0) <='0';
          end if;
        if(cVar1S6S114P018P064P007P059(0)='1' AND  A( 3)='0' AND A( 8)='0' AND D( 8)='1' )then
          cVar2S6S114P013N003P067nsss(0) <='1';
          else
          cVar2S6S114P013N003P067nsss(0) <='0';
          end if;
        if(cVar1S7S114P018P064P007P059(0)='1' AND  A( 3)='1' AND B( 9)='1' )then
          cVar2S7S114P013P036nsss(0) <='1';
          else
          cVar2S7S114P013P036nsss(0) <='0';
          end if;
        if(cVar1S8S114P018N064P050P034(0)='1' AND  B( 2)='1' AND D(10)='0' AND A(15)='0' )then
          cVar2S8S114P033P059P008nsss(0) <='1';
          else
          cVar2S8S114P033P059P008nsss(0) <='0';
          end if;
        if(cVar1S9S114P018N064P050P034(0)='1' AND  B( 2)='0' AND B(13)='0' AND B( 1)='0' )then
          cVar2S9S114N033P028P035nsss(0) <='1';
          else
          cVar2S9S114N033P028P035nsss(0) <='0';
          end if;
        if(cVar1S10S114P018N064P050N034(0)='1' AND  A( 6)='1' AND D(10)='1' AND A( 0)='0' )then
          cVar2S10S114P007P059P019nsss(0) <='1';
          else
          cVar2S10S114P007P059P019nsss(0) <='0';
          end if;
        if(cVar1S11S114P018N064P050N034(0)='1' AND  A( 6)='1' AND D(10)='0' AND E( 9)='1' )then
          cVar2S11S114P007N059P065nsss(0) <='1';
          else
          cVar2S11S114P007N059P065nsss(0) <='0';
          end if;
        if(cVar1S12S114P018N064P050N034(0)='1' AND  A( 6)='0' AND B( 1)='1' )then
          cVar2S12S114N007P035nsss(0) <='1';
          else
          cVar2S12S114N007P035nsss(0) <='0';
          end if;
        if(cVar1S13S114P018N064P050N034(0)='1' AND  A( 6)='0' AND B( 1)='0' AND D( 1)='0' )then
          cVar2S13S114N007N035P062nsss(0) <='1';
          else
          cVar2S13S114N007N035P062nsss(0) <='0';
          end if;
        if(cVar1S14S114P018N064P050P008(0)='1' AND  B( 4)='1' )then
          cVar2S14S114P029nsss(0) <='1';
          else
          cVar2S14S114P029nsss(0) <='0';
          end if;
        if(cVar1S15S114P018N064P050P008(0)='1' AND  B( 4)='0' AND B( 9)='0' )then
          cVar2S15S114N029P036nsss(0) <='1';
          else
          cVar2S15S114N029P036nsss(0) <='0';
          end if;
        if(cVar1S16S114P018N064P050N008(0)='1' AND  A( 3)='0' AND B(13)='1' )then
          cVar2S16S114P013P028nsss(0) <='1';
          else
          cVar2S16S114P013P028nsss(0) <='0';
          end if;
        if(cVar1S17S114P018N064P050N008(0)='1' AND  A( 3)='0' AND B(13)='0' AND A(13)='1' )then
          cVar2S17S114P013N028P012nsss(0) <='1';
          else
          cVar2S17S114P013N028P012nsss(0) <='0';
          end if;
        if(cVar1S18S114P018N064P050N008(0)='1' AND  A( 3)='1' AND A(11)='0' AND A(12)='1' )then
          cVar2S18S114P013P016P014nsss(0) <='1';
          else
          cVar2S18S114P013P016P014nsss(0) <='0';
          end if;
        if(cVar1S19S114N018P014P035P015(0)='1' AND  B( 8)='0' AND A( 4)='0' )then
          cVar2S19S114P021P011nsss(0) <='1';
          else
          cVar2S19S114P021P011nsss(0) <='0';
          end if;
        if(cVar1S20S114N018P014P035P015(0)='1' AND  B( 8)='0' AND A( 4)='1' AND A(13)='0' )then
          cVar2S20S114P021P011P012nsss(0) <='1';
          else
          cVar2S20S114P021P011P012nsss(0) <='0';
          end if;
        if(cVar1S21S114N018P014P035P015(0)='1' AND  B( 8)='1' AND A(14)='0' AND B( 0)='1' )then
          cVar2S21S114P021P010P037nsss(0) <='1';
          else
          cVar2S21S114P021P010P037nsss(0) <='0';
          end if;
        if(cVar1S22S114N018P014P035P015(0)='1' AND  B( 2)='0' AND B(11)='1' AND B( 9)='0' )then
          cVar2S22S114P033P032P036nsss(0) <='1';
          else
          cVar2S22S114P033P032P036nsss(0) <='0';
          end if;
        if(cVar1S23S114N018P014P035P015(0)='1' AND  B( 2)='0' AND B(11)='0' AND B(10)='1' )then
          cVar2S23S114P033N032P034nsss(0) <='1';
          else
          cVar2S23S114P033N032P034nsss(0) <='0';
          end if;
        if(cVar1S24S114N018P014P035P015(0)='1' AND  B( 2)='1' AND B(11)='0' AND A( 6)='0' )then
          cVar2S24S114P033P032P007nsss(0) <='1';
          else
          cVar2S24S114P033P032P007nsss(0) <='0';
          end if;
        if(cVar1S25S114N018P014P035P015(0)='1' AND  B( 2)='1' AND B(11)='1' AND D(10)='0' )then
          cVar2S25S114P033P032P059nsss(0) <='1';
          else
          cVar2S25S114P033P032P059nsss(0) <='0';
          end if;
        if(cVar1S26S114N018P014P035P024(0)='1' AND  B(10)='0' AND E( 7)='0' AND A(14)='0' )then
          cVar2S26S114P034P040P010nsss(0) <='1';
          else
          cVar2S26S114P034P040P010nsss(0) <='0';
          end if;
        if(cVar1S27S114N018P014P035P024(0)='1' AND  B(10)='1' AND A( 1)='1' AND A(11)='1' )then
          cVar2S27S114P034P017P016nsss(0) <='1';
          else
          cVar2S27S114P034P017P016nsss(0) <='0';
          end if;
        if(cVar1S28S114N018P014P035P024(0)='1' AND  B(10)='1' AND A( 1)='0' AND B( 2)='1' )then
          cVar2S28S114P034N017P033nsss(0) <='1';
          else
          cVar2S28S114P034N017P033nsss(0) <='0';
          end if;
        if(cVar1S29S114N018N014P010P030(0)='1' AND  E( 3)='0' AND A(13)='1' )then
          cVar2S29S114P056P012nsss(0) <='1';
          else
          cVar2S29S114P056P012nsss(0) <='0';
          end if;
        if(cVar1S30S114N018N014P010P030(0)='1' AND  E( 3)='0' AND A(13)='0' AND B( 0)='0' )then
          cVar2S30S114P056N012P037nsss(0) <='1';
          else
          cVar2S30S114P056N012P037nsss(0) <='0';
          end if;
        if(cVar1S31S114N018N014P010P030(0)='1' AND  E( 3)='1' AND A(13)='0' AND E(11)='0' )then
          cVar2S31S114P056P012P057nsss(0) <='1';
          else
          cVar2S31S114P056P012P057nsss(0) <='0';
          end if;
        if(cVar1S32S114N018N014P010N030(0)='1' AND  A( 3)='1' AND E( 2)='0' AND D(10)='0' )then
          cVar2S32S114P013P060P059nsss(0) <='1';
          else
          cVar2S32S114P013P060P059nsss(0) <='0';
          end if;
        if(cVar1S33S114N018N014P010N030(0)='1' AND  A( 3)='0' AND A(11)='0' AND B( 0)='0' )then
          cVar2S33S114N013P016P037nsss(0) <='1';
          else
          cVar2S33S114N013P016P037nsss(0) <='0';
          end if;
        if(cVar1S34S114N018N014P010N030(0)='1' AND  A( 3)='0' AND A(11)='1' AND E( 0)='1' )then
          cVar2S34S114N013P016P068nsss(0) <='1';
          else
          cVar2S34S114N013P016P068nsss(0) <='0';
          end if;
        if(cVar1S35S114N018N014N010P011(0)='1' AND  A( 6)='0' )then
          cVar2S35S114P007nsss(0) <='1';
          else
          cVar2S35S114P007nsss(0) <='0';
          end if;
        if(cVar1S36S114N018N014N010P011(0)='1' AND  A( 6)='1' AND D( 1)='1' AND A( 2)='0' )then
          cVar2S36S114P007P062P015nsss(0) <='1';
          else
          cVar2S36S114P007P062P015nsss(0) <='0';
          end if;
        if(cVar1S37S114N018N014N010N011(0)='1' AND  A( 1)='0' AND A( 2)='1' AND D( 9)='1' )then
          cVar2S37S114P017P015P063nsss(0) <='1';
          else
          cVar2S37S114P017P015P063nsss(0) <='0';
          end if;
        if(cVar1S38S114N018N014N010N011(0)='1' AND  A( 1)='1' AND E( 6)='1' )then
          cVar2S38S114P017P044nsss(0) <='1';
          else
          cVar2S38S114P017P044nsss(0) <='0';
          end if;
        if(cVar1S0S115P018P014P069P065(0)='1' AND  B(13)='1' AND A( 0)='1' )then
          cVar2S0S115P028P019nsss(0) <='1';
          else
          cVar2S0S115P028P019nsss(0) <='0';
          end if;
        if(cVar1S1S115P018P014P069P065(0)='1' AND  B(13)='1' AND A( 0)='0' AND E( 0)='1' )then
          cVar2S1S115P028N019P068nsss(0) <='1';
          else
          cVar2S1S115P028N019P068nsss(0) <='0';
          end if;
        if(cVar1S2S115P018P014P069P065(0)='1' AND  B(13)='0' AND B( 0)='1' )then
          cVar2S2S115N028P037nsss(0) <='1';
          else
          cVar2S2S115N028P037nsss(0) <='0';
          end if;
        if(cVar1S3S115P018P014P069P065(0)='1' AND  B(13)='0' AND B( 0)='0' AND A(11)='0' )then
          cVar2S3S115N028N037P016nsss(0) <='1';
          else
          cVar2S3S115N028N037P016nsss(0) <='0';
          end if;
        if(cVar1S4S115P018P014P069P065(0)='1' AND  A(11)='1' AND B( 0)='0' AND D(10)='0' )then
          cVar2S4S115P016P037P059nsss(0) <='1';
          else
          cVar2S4S115P016P037P059nsss(0) <='0';
          end if;
        if(cVar1S5S115P018P014P069P065(0)='1' AND  A(11)='1' AND B( 0)='1' AND D( 1)='1' )then
          cVar2S5S115P016P037P062nsss(0) <='1';
          else
          cVar2S5S115P016P037P062nsss(0) <='0';
          end if;
        if(cVar1S6S115P018P014P069P065(0)='1' AND  A(11)='0' AND E( 2)='1' )then
          cVar2S6S115N016P060nsss(0) <='1';
          else
          cVar2S6S115N016P060nsss(0) <='0';
          end if;
        if(cVar1S7S115P018P014N069P067(0)='1' AND  A( 4)='0' AND A( 3)='1' AND B( 9)='0' )then
          cVar2S7S115P011P013P036nsss(0) <='1';
          else
          cVar2S7S115P011P013P036nsss(0) <='0';
          end if;
        if(cVar1S8S115P018P014N069P067(0)='1' AND  A( 4)='0' AND A( 3)='0' AND D( 3)='0' )then
          cVar2S8S115P011N013P054nsss(0) <='1';
          else
          cVar2S8S115P011N013P054nsss(0) <='0';
          end if;
        if(cVar1S9S115P018P014N069P067(0)='1' AND  A( 4)='1' AND D( 0)='0' )then
          cVar2S9S115P011P066nsss(0) <='1';
          else
          cVar2S9S115P011P066nsss(0) <='0';
          end if;
        if(cVar1S10S115P018P014N069P067(0)='1' AND  A( 4)='1' AND D( 0)='1' AND B( 6)='1' )then
          cVar2S10S115P011P066P025nsss(0) <='1';
          else
          cVar2S10S115P011P066P025nsss(0) <='0';
          end if;
        if(cVar1S11S115P018P014N069P067(0)='1' AND  A( 0)='1' AND B( 9)='1' AND A( 2)='0' )then
          cVar2S11S115P019P036P015nsss(0) <='1';
          else
          cVar2S11S115P019P036P015nsss(0) <='0';
          end if;
        if(cVar1S12S115P018P014N069P067(0)='1' AND  A( 0)='1' AND B( 9)='0' AND A(14)='0' )then
          cVar2S12S115P019N036P010nsss(0) <='1';
          else
          cVar2S12S115P019N036P010nsss(0) <='0';
          end if;
        if(cVar1S13S115P018P014N069P067(0)='1' AND  A( 0)='0' AND D( 1)='1' AND D( 0)='0' )then
          cVar2S13S115N019P062P066nsss(0) <='1';
          else
          cVar2S13S115N019P062P066nsss(0) <='0';
          end if;
        if(cVar1S14S115P018P014P007P064(0)='1' AND  B( 9)='0' AND B(12)='1' )then
          cVar2S14S115P036P030nsss(0) <='1';
          else
          cVar2S14S115P036P030nsss(0) <='0';
          end if;
        if(cVar1S15S115P018P014P007P064(0)='1' AND  B( 9)='0' AND B(12)='0' AND A(13)='0' )then
          cVar2S15S115P036N030P012nsss(0) <='1';
          else
          cVar2S15S115P036N030P012nsss(0) <='0';
          end if;
        if(cVar1S16S115P018P014P007P064(0)='1' AND  B( 9)='1' AND E(12)='0' AND A( 0)='1' )then
          cVar2S16S115P036P053P019nsss(0) <='1';
          else
          cVar2S16S115P036P053P019nsss(0) <='0';
          end if;
        if(cVar1S17S115P018P014P007P064(0)='1' AND  B(11)='1' AND E( 8)='1' )then
          cVar2S17S115P032P069nsss(0) <='1';
          else
          cVar2S17S115P032P069nsss(0) <='0';
          end if;
        if(cVar1S18S115P018P014P007P064(0)='1' AND  B(11)='1' AND E( 8)='0' AND B( 1)='1' )then
          cVar2S18S115P032N069P035nsss(0) <='1';
          else
          cVar2S18S115P032N069P035nsss(0) <='0';
          end if;
        if(cVar1S19S115P018P014P007P064(0)='1' AND  B(11)='0' AND A( 9)='1' )then
          cVar2S19S115N032P001nsss(0) <='1';
          else
          cVar2S19S115N032P001nsss(0) <='0';
          end if;
        if(cVar1S20S115P018P014P007P037(0)='1' AND  A(16)='1' )then
          cVar2S20S115P006nsss(0) <='1';
          else
          cVar2S20S115P006nsss(0) <='0';
          end if;
        if(cVar1S21S115P018P014P007P037(0)='1' AND  A(16)='0' AND A(11)='1' AND A(15)='0' )then
          cVar2S21S115N006P016P008nsss(0) <='1';
          else
          cVar2S21S115N006P016P008nsss(0) <='0';
          end if;
        if(cVar1S22S115P018P014P007P037(0)='1' AND  A(16)='0' AND A(11)='0' AND A( 4)='1' )then
          cVar2S22S115N006N016P011nsss(0) <='1';
          else
          cVar2S22S115N006N016P011nsss(0) <='0';
          end if;
        if(cVar1S23S115P018P014P007N037(0)='1' AND  E(14)='1' )then
          cVar2S23S115P045nsss(0) <='1';
          else
          cVar2S23S115P045nsss(0) <='0';
          end if;
        if(cVar1S24S115P018P014P007N037(0)='1' AND  E(14)='0' AND A(18)='1' AND A( 2)='0' )then
          cVar2S24S115N045P002P015nsss(0) <='1';
          else
          cVar2S24S115N045P002P015nsss(0) <='0';
          end if;
        if(cVar1S25S115P018P014P007N037(0)='1' AND  E(14)='0' AND A(18)='0' AND D(12)='1' )then
          cVar2S25S115N045N002P051nsss(0) <='1';
          else
          cVar2S25S115N045N002P051nsss(0) <='0';
          end if;
        if(cVar1S26S115P018P062P066P042(0)='1' AND  A( 6)='0' AND D(13)='1' )then
          cVar2S26S115P007P047nsss(0) <='1';
          else
          cVar2S26S115P007P047nsss(0) <='0';
          end if;
        if(cVar1S27S115P018P062P066P042(0)='1' AND  A( 6)='0' AND D(13)='0' AND B( 8)='0' )then
          cVar2S27S115P007N047P021nsss(0) <='1';
          else
          cVar2S27S115P007N047P021nsss(0) <='0';
          end if;
        if(cVar1S28S115P018P062P066P042(0)='1' AND  A( 6)='1' AND D(10)='0' AND A( 3)='0' )then
          cVar2S28S115P007P059P013nsss(0) <='1';
          else
          cVar2S28S115P007P059P013nsss(0) <='0';
          end if;
        if(cVar1S29S115P018P062P066P068(0)='1' AND  E(10)='1' )then
          cVar2S29S115P061nsss(0) <='1';
          else
          cVar2S29S115P061nsss(0) <='0';
          end if;
        if(cVar1S30S115P018P062P066P068(0)='1' AND  E(10)='0' AND B( 0)='0' AND B( 1)='1' )then
          cVar2S30S115N061P037P035nsss(0) <='1';
          else
          cVar2S30S115N061P037P035nsss(0) <='0';
          end if;
        if(cVar1S31S115P018P062P066N068(0)='1' AND  A( 7)='1' )then
          cVar2S31S115P005nsss(0) <='1';
          else
          cVar2S31S115P005nsss(0) <='0';
          end if;
        if(cVar1S32S115P018P062P066N068(0)='1' AND  A( 7)='0' AND A( 5)='1' )then
          cVar2S32S115N005P009nsss(0) <='1';
          else
          cVar2S32S115N005P009nsss(0) <='0';
          end if;
        if(cVar1S33S115P018N062P007P047(0)='1' AND  D( 0)='1' )then
          cVar2S33S115P066nsss(0) <='1';
          else
          cVar2S33S115P066nsss(0) <='0';
          end if;
        if(cVar1S34S115P018N062P007P047(0)='1' AND  D( 0)='0' AND D( 8)='0' )then
          cVar2S34S115N066P067nsss(0) <='1';
          else
          cVar2S34S115N066P067nsss(0) <='0';
          end if;
        if(cVar1S35S115P018N062P007N047(0)='1' AND  D(10)='1' AND E( 9)='0' )then
          cVar2S35S115P059P065nsss(0) <='1';
          else
          cVar2S35S115P059P065nsss(0) <='0';
          end if;
        if(cVar1S36S115P018N062P007N047(0)='1' AND  D(10)='0' AND B(13)='1' )then
          cVar2S36S115N059P028nsss(0) <='1';
          else
          cVar2S36S115N059P028nsss(0) <='0';
          end if;
        if(cVar1S37S115P018N062P007N047(0)='1' AND  D(10)='0' AND B(13)='0' AND B(11)='0' )then
          cVar2S37S115N059N028P032nsss(0) <='1';
          else
          cVar2S37S115N059N028P032nsss(0) <='0';
          end if;
        if(cVar1S38S115P018N062N007P034(0)='1' AND  B( 2)='1' AND A( 5)='1' )then
          cVar2S38S115P033P009nsss(0) <='1';
          else
          cVar2S38S115P033P009nsss(0) <='0';
          end if;
        if(cVar1S39S115P018N062N007P034(0)='1' AND  B( 2)='1' AND A( 5)='0' AND E( 2)='1' )then
          cVar2S39S115P033N009P060nsss(0) <='1';
          else
          cVar2S39S115P033N009P060nsss(0) <='0';
          end if;
        if(cVar1S40S115P018N062N007P034(0)='1' AND  B( 2)='0' AND B(13)='0' AND D( 8)='0' )then
          cVar2S40S115N033P028P067nsss(0) <='1';
          else
          cVar2S40S115N033P028P067nsss(0) <='0';
          end if;
        if(cVar1S41S115P018N062N007N034(0)='1' AND  D( 2)='1' AND B(11)='1' AND E( 2)='1' )then
          cVar2S41S115P058P032P060nsss(0) <='1';
          else
          cVar2S41S115P058P032P060nsss(0) <='0';
          end if;
        if(cVar1S42S115P018N062N007N034(0)='1' AND  D( 2)='1' AND B(11)='0' AND B( 3)='1' )then
          cVar2S42S115P058N032P031nsss(0) <='1';
          else
          cVar2S42S115P058N032P031nsss(0) <='0';
          end if;
        if(cVar1S0S116P018P063P049P059(0)='1' AND  B(14)='1' )then
          cVar2S0S116P026nsss(0) <='1';
          else
          cVar2S0S116P026nsss(0) <='0';
          end if;
        if(cVar1S1S116P018P063P049P059(0)='1' AND  B(14)='0' AND A(16)='1' )then
          cVar2S1S116N026P006nsss(0) <='1';
          else
          cVar2S1S116N026P006nsss(0) <='0';
          end if;
        if(cVar1S2S116P018P063P049P059(0)='1' AND  B(14)='0' AND A(16)='0' AND D( 2)='1' )then
          cVar2S2S116N026N006P058nsss(0) <='1';
          else
          cVar2S2S116N026N006P058nsss(0) <='0';
          end if;
        if(cVar1S3S116P018P063N049P066(0)='1' AND  D( 5)='1' )then
          cVar2S3S116P046nsss(0) <='1';
          else
          cVar2S3S116P046nsss(0) <='0';
          end if;
        if(cVar1S4S116P018P063N049P066(0)='1' AND  D( 5)='0' AND E( 8)='0' AND A(14)='0' )then
          cVar2S4S116N046P069P010nsss(0) <='1';
          else
          cVar2S4S116N046P069P010nsss(0) <='0';
          end if;
        if(cVar1S5S116P018P063N049P066(0)='1' AND  D( 5)='0' AND E( 8)='1' )then
          cVar2S5S116N046P069psss(0) <='1';
          else
          cVar2S5S116N046P069psss(0) <='0';
          end if;
        if(cVar1S6S116P018P063N049N066(0)='1' AND  E( 5)='0' AND B(13)='1' )then
          cVar2S6S116P048P028nsss(0) <='1';
          else
          cVar2S6S116P048P028nsss(0) <='0';
          end if;
        if(cVar1S7S116P018P063N049N066(0)='1' AND  E( 5)='0' AND B(13)='0' AND E(10)='1' )then
          cVar2S7S116P048N028P061nsss(0) <='1';
          else
          cVar2S7S116P048N028P061nsss(0) <='0';
          end if;
        if(cVar1S8S116P018P063N049N066(0)='1' AND  E( 5)='1' AND A(16)='1' AND A( 1)='0' )then
          cVar2S8S116P048P006P017nsss(0) <='1';
          else
          cVar2S8S116P048P006P017nsss(0) <='0';
          end if;
        if(cVar1S9S116P018P063N049N066(0)='1' AND  E( 5)='1' AND A(16)='0' AND B(14)='1' )then
          cVar2S9S116P048N006P026nsss(0) <='1';
          else
          cVar2S9S116P048N006P026nsss(0) <='0';
          end if;
        if(cVar1S10S116P018P063P031P056(0)='1' AND  A(13)='1' )then
          cVar2S10S116P012nsss(0) <='1';
          else
          cVar2S10S116P012nsss(0) <='0';
          end if;
        if(cVar1S11S116P018P063P031P056(0)='1' AND  A(13)='0' AND A(11)='0' )then
          cVar2S11S116N012P016nsss(0) <='1';
          else
          cVar2S11S116N012P016nsss(0) <='0';
          end if;
        if(cVar1S12S116P018P063P031N056(0)='1' AND  B( 1)='0' AND B( 9)='1' )then
          cVar2S12S116P035P036nsss(0) <='1';
          else
          cVar2S12S116P035P036nsss(0) <='0';
          end if;
        if(cVar1S13S116P018P063N031P033(0)='1' AND  A( 2)='0' AND B( 9)='1' AND E( 8)='0' )then
          cVar2S13S116P015P036P069nsss(0) <='1';
          else
          cVar2S13S116P015P036P069nsss(0) <='0';
          end if;
        if(cVar1S14S116P018P063N031P033(0)='1' AND  A( 2)='0' AND B( 9)='0' AND B( 0)='1' )then
          cVar2S14S116P015N036P037nsss(0) <='1';
          else
          cVar2S14S116P015N036P037nsss(0) <='0';
          end if;
        if(cVar1S15S116P018P063N031P033(0)='1' AND  A( 2)='1' AND E( 9)='1' AND E( 1)='1' )then
          cVar2S15S116P015P065P064nsss(0) <='1';
          else
          cVar2S15S116P015P065P064nsss(0) <='0';
          end if;
        if(cVar1S16S116P018P063N031P033(0)='1' AND  A( 2)='1' AND E( 9)='0' AND A( 1)='0' )then
          cVar2S16S116P015N065P017nsss(0) <='1';
          else
          cVar2S16S116P015N065P017nsss(0) <='0';
          end if;
        if(cVar1S17S116P018P063N031N033(0)='1' AND  A(18)='0' AND D( 8)='1' AND D(10)='0' )then
          cVar2S17S116P002P067P059nsss(0) <='1';
          else
          cVar2S17S116P002P067P059nsss(0) <='0';
          end if;
        if(cVar1S18S116P018P063N031N033(0)='1' AND  A(18)='0' AND D( 8)='0' AND A( 3)='1' )then
          cVar2S18S116P002N067P013nsss(0) <='1';
          else
          cVar2S18S116P002N067P013nsss(0) <='0';
          end if;
        if(cVar1S19S116P018P063N031N033(0)='1' AND  A(18)='1' AND A( 2)='0' AND A( 0)='1' )then
          cVar2S19S116P002N015P019nsss(0) <='1';
          else
          cVar2S19S116P002N015P019nsss(0) <='0';
          end if;
        if(cVar1S20S116N018P069P064P019(0)='1' AND  A( 1)='0' AND B( 0)='0' AND A(11)='1' )then
          cVar2S20S116P017P037P016nsss(0) <='1';
          else
          cVar2S20S116P017P037P016nsss(0) <='0';
          end if;
        if(cVar1S21S116N018P069P064P019(0)='1' AND  A( 1)='0' AND B( 0)='1' AND A( 2)='1' )then
          cVar2S21S116P017P037P015nsss(0) <='1';
          else
          cVar2S21S116P017P037P015nsss(0) <='0';
          end if;
        if(cVar1S22S116N018P069P064P019(0)='1' AND  A( 1)='1' AND A(11)='0' )then
          cVar2S22S116P017P016nsss(0) <='1';
          else
          cVar2S22S116P017P016nsss(0) <='0';
          end if;
        if(cVar1S23S116N018P069P064P019(0)='1' AND  A( 1)='1' AND A(11)='1' AND B( 0)='1' )then
          cVar2S23S116P017P016P037nsss(0) <='1';
          else
          cVar2S23S116P017P016P037nsss(0) <='0';
          end if;
        if(cVar1S24S116N018P069P064P019(0)='1' AND  A(13)='1' AND A( 2)='0' )then
          cVar2S24S116P012P015nsss(0) <='1';
          else
          cVar2S24S116P012P015nsss(0) <='0';
          end if;
        if(cVar1S25S116N018P069P064P019(0)='1' AND  A(13)='0' AND A( 1)='1' AND E( 0)='0' )then
          cVar2S25S116N012P017P068nsss(0) <='1';
          else
          cVar2S25S116N012P017P068nsss(0) <='0';
          end if;
        if(cVar1S26S116N018P069P064P019(0)='1' AND  A(13)='0' AND A( 1)='0' AND A( 2)='1' )then
          cVar2S26S116N012N017P015nsss(0) <='1';
          else
          cVar2S26S116N012N017P015nsss(0) <='0';
          end if;
        if(cVar1S27S116N018P069N064P065(0)='1' AND  E(14)='1' AND D(13)='1' )then
          cVar2S27S116P045P047nsss(0) <='1';
          else
          cVar2S27S116P045P047nsss(0) <='0';
          end if;
        if(cVar1S28S116N018P069N064P065(0)='1' AND  E(14)='1' AND D(13)='0' AND A( 0)='1' )then
          cVar2S28S116P045N047P019nsss(0) <='1';
          else
          cVar2S28S116P045N047P019nsss(0) <='0';
          end if;
        if(cVar1S29S116N018P069N064P065(0)='1' AND  E(14)='0' AND D(14)='0' AND E(15)='1' )then
          cVar2S29S116N045P043P041nsss(0) <='1';
          else
          cVar2S29S116N045P043P041nsss(0) <='0';
          end if;
        if(cVar1S30S116N018P069N064P065(0)='1' AND  E( 2)='1' AND B( 9)='1' )then
          cVar2S30S116P060P036nsss(0) <='1';
          else
          cVar2S30S116P060P036nsss(0) <='0';
          end if;
        if(cVar1S31S116N018P069N064P065(0)='1' AND  E( 2)='0' AND B(10)='1' AND D( 8)='1' )then
          cVar2S31S116N060P034P067nsss(0) <='1';
          else
          cVar2S31S116N060P034P067nsss(0) <='0';
          end if;
        if(cVar1S32S116N018N069P056P012(0)='1' AND  A(14)='0' AND B(10)='1' AND D( 3)='1' )then
          cVar2S32S116P010P034P054nsss(0) <='1';
          else
          cVar2S32S116P010P034P054nsss(0) <='0';
          end if;
        if(cVar1S33S116N018N069P056P012(0)='1' AND  A(14)='0' AND B(10)='0' AND E( 9)='0' )then
          cVar2S33S116P010N034P065nsss(0) <='1';
          else
          cVar2S33S116P010N034P065nsss(0) <='0';
          end if;
        if(cVar1S34S116N018N069P056P012(0)='1' AND  A(14)='1' AND A( 3)='0' AND E( 0)='1' )then
          cVar2S34S116P010P013P068nsss(0) <='1';
          else
          cVar2S34S116P010P013P068nsss(0) <='0';
          end if;
        if(cVar1S35S116N018N069P056N012(0)='1' AND  A( 7)='0' AND D(13)='0' AND B(12)='1' )then
          cVar2S35S116P005P047P030nsss(0) <='1';
          else
          cVar2S35S116P005P047P030nsss(0) <='0';
          end if;
        if(cVar1S36S116N018N069N056P013(0)='1' AND  D( 2)='1' AND A(15)='1' )then
          cVar2S36S116P058P008nsss(0) <='1';
          else
          cVar2S36S116P058P008nsss(0) <='0';
          end if;
        if(cVar1S37S116N018N069N056P013(0)='1' AND  D( 2)='1' AND A(15)='0' AND B(17)='0' )then
          cVar2S37S116P058N008P020nsss(0) <='1';
          else
          cVar2S37S116P058N008P020nsss(0) <='0';
          end if;
        if(cVar1S38S116N018N069N056P013(0)='1' AND  D( 2)='0' AND A(15)='0' AND B( 0)='1' )then
          cVar2S38S116N058P008P037nsss(0) <='1';
          else
          cVar2S38S116N058P008P037nsss(0) <='0';
          end if;
        if(cVar1S39S116N018N069N056P013(0)='1' AND  D( 2)='0' AND A(15)='1' AND B(13)='1' )then
          cVar2S39S116N058P008P028nsss(0) <='1';
          else
          cVar2S39S116N058P008P028nsss(0) <='0';
          end if;
        if(cVar1S40S116N018N069N056N013(0)='1' AND  B( 2)='0' AND B( 9)='1' AND E(15)='0' )then
          cVar2S40S116P033P036P041nsss(0) <='1';
          else
          cVar2S40S116P033P036P041nsss(0) <='0';
          end if;
        if(cVar1S41S116N018N069N056N013(0)='1' AND  B( 2)='0' AND B( 9)='0' AND D(15)='1' )then
          cVar2S41S116P033N036P039nsss(0) <='1';
          else
          cVar2S41S116P033N036P039nsss(0) <='0';
          end if;
        if(cVar1S0S117P066P069P063P067(0)='1' AND  A(11)='1' )then
          cVar2S0S117P016nsss(0) <='1';
          else
          cVar2S0S117P016nsss(0) <='0';
          end if;
        if(cVar1S1S117P066P069P063P067(0)='1' AND  A(11)='0' AND B( 2)='0' )then
          cVar2S1S117N016P033nsss(0) <='1';
          else
          cVar2S1S117N016P033nsss(0) <='0';
          end if;
        if(cVar1S2S117P066P069P063N067(0)='1' AND  B( 1)='1' AND E( 1)='1' )then
          cVar2S2S117P035P064nsss(0) <='1';
          else
          cVar2S2S117P035P064nsss(0) <='0';
          end if;
        if(cVar1S3S117P066P069P063N067(0)='1' AND  B( 1)='0' AND A( 3)='1' AND A( 0)='0' )then
          cVar2S3S117N035P013P019nsss(0) <='1';
          else
          cVar2S3S117N035P013P019nsss(0) <='0';
          end if;
        if(cVar1S4S117P066P069P063P061(0)='1' AND  E( 9)='1' AND B(13)='0' )then
          cVar2S4S117P065P028nsss(0) <='1';
          else
          cVar2S4S117P065P028nsss(0) <='0';
          end if;
        if(cVar1S5S117P066P069P063P061(0)='1' AND  E( 9)='0' AND A( 0)='0' AND A( 1)='1' )then
          cVar2S5S117N065P019P017nsss(0) <='1';
          else
          cVar2S5S117N065P019P017nsss(0) <='0';
          end if;
        if(cVar1S6S117P066P069P063P061(0)='1' AND  D( 2)='1' )then
          cVar2S6S117P058nsss(0) <='1';
          else
          cVar2S6S117P058nsss(0) <='0';
          end if;
        if(cVar1S7S117P066N069P068P047(0)='1' AND  A(10)='1' AND D(12)='0' AND E(13)='1' )then
          cVar2S7S117P018P051P049nsss(0) <='1';
          else
          cVar2S7S117P018P051P049nsss(0) <='0';
          end if;
        if(cVar1S8S117P066N069P068P047(0)='1' AND  A(10)='0' AND E(13)='1' AND E( 5)='0' )then
          cVar2S8S117N018P049P048nsss(0) <='1';
          else
          cVar2S8S117N018P049P048nsss(0) <='0';
          end if;
        if(cVar1S9S117P066N069P068P047(0)='1' AND  A(10)='0' AND E(13)='0' AND E(12)='1' )then
          cVar2S9S117N018N049P053nsss(0) <='1';
          else
          cVar2S9S117N018N049P053nsss(0) <='0';
          end if;
        if(cVar1S10S117P066N069P068N047(0)='1' AND  B( 3)='1' AND A( 6)='0' AND A( 5)='0' )then
          cVar2S10S117P031P007P009nsss(0) <='1';
          else
          cVar2S10S117P031P007P009nsss(0) <='0';
          end if;
        if(cVar1S11S117P066N069P068N047(0)='1' AND  B( 3)='1' AND A( 6)='1' AND A( 0)='1' )then
          cVar2S11S117P031P007P019nsss(0) <='1';
          else
          cVar2S11S117P031P007P019nsss(0) <='0';
          end if;
        if(cVar1S12S117P066N069P068N047(0)='1' AND  B( 3)='0' AND B( 1)='1' )then
          cVar2S12S117N031P035nsss(0) <='1';
          else
          cVar2S12S117N031P035nsss(0) <='0';
          end if;
        if(cVar1S13S117P066N069P068N047(0)='1' AND  B( 3)='0' AND B( 1)='0' AND D(14)='1' )then
          cVar2S13S117N031N035P043nsss(0) <='1';
          else
          cVar2S13S117N031N035P043nsss(0) <='0';
          end if;
        if(cVar1S14S117P066N069P068P064(0)='1' AND  B( 1)='0' AND D( 1)='1' )then
          cVar2S14S117P035P062nsss(0) <='1';
          else
          cVar2S14S117P035P062nsss(0) <='0';
          end if;
        if(cVar1S15S117P066N069P068P064(0)='1' AND  B( 1)='1' AND B( 0)='0' AND A(11)='1' )then
          cVar2S15S117P035P037P016nsss(0) <='1';
          else
          cVar2S15S117P035P037P016nsss(0) <='0';
          end if;
        if(cVar1S16S117P066N069P068N064(0)='1' AND  B( 5)='1' )then
          cVar2S16S117P027nsss(0) <='1';
          else
          cVar2S16S117P027nsss(0) <='0';
          end if;
        if(cVar1S17S117P066P018P006P047(0)='1' AND  A(14)='0' AND A(18)='0' AND A( 3)='0' )then
          cVar2S17S117P010P002P013nsss(0) <='1';
          else
          cVar2S17S117P010P002P013nsss(0) <='0';
          end if;
        if(cVar1S18S117P066P018P006P047(0)='1' AND  A(14)='0' AND A(18)='1' AND B( 0)='1' )then
          cVar2S18S117P010P002P037nsss(0) <='1';
          else
          cVar2S18S117P010P002P037nsss(0) <='0';
          end if;
        if(cVar1S19S117P066P018P006P047(0)='1' AND  A(14)='1' AND D( 3)='1' AND A( 4)='0' )then
          cVar2S19S117P010P054P011nsss(0) <='1';
          else
          cVar2S19S117P010P054P011nsss(0) <='0';
          end if;
        if(cVar1S20S117P066P018P006P047(0)='1' AND  A(14)='1' AND D( 3)='0' AND D( 4)='1' )then
          cVar2S20S117P010N054P050nsss(0) <='1';
          else
          cVar2S20S117P010N054P050nsss(0) <='0';
          end if;
        if(cVar1S21S117P066P018P006P047(0)='1' AND  B(15)='1' AND A( 0)='1' )then
          cVar2S21S117P024P019nsss(0) <='1';
          else
          cVar2S21S117P024P019nsss(0) <='0';
          end if;
        if(cVar1S22S117P066P018P006P047(0)='1' AND  B(15)='0' AND A(14)='1' )then
          cVar2S22S117N024P010nsss(0) <='1';
          else
          cVar2S22S117N024P010nsss(0) <='0';
          end if;
        if(cVar1S23S117P066P018P006P024(0)='1' AND  A( 0)='0' )then
          cVar2S23S117P019nsss(0) <='1';
          else
          cVar2S23S117P019nsss(0) <='0';
          end if;
        if(cVar1S24S117P066P018P006P024(0)='1' AND  A( 0)='1' AND E(13)='0' )then
          cVar2S24S117P019P049nsss(0) <='1';
          else
          cVar2S24S117P019P049nsss(0) <='0';
          end if;
        if(cVar1S25S117P066P018P006N024(0)='1' AND  E( 8)='1' AND A(11)='1' )then
          cVar2S25S117P069P016nsss(0) <='1';
          else
          cVar2S25S117P069P016nsss(0) <='0';
          end if;
        if(cVar1S26S117P066P018P006N024(0)='1' AND  E( 8)='0' AND E( 5)='1' )then
          cVar2S26S117N069P048nsss(0) <='1';
          else
          cVar2S26S117N069P048nsss(0) <='0';
          end if;
        if(cVar1S28S117P066P018P049N051(0)='1' AND  E( 0)='1' AND A( 5)='0' AND A( 1)='0' )then
          cVar2S28S117P068P009P017nsss(0) <='1';
          else
          cVar2S28S117P068P009P017nsss(0) <='0';
          end if;
        if(cVar1S29S117P066P018P049N051(0)='1' AND  E( 0)='1' AND A( 5)='1' AND B( 0)='1' )then
          cVar2S29S117P068P009P037nsss(0) <='1';
          else
          cVar2S29S117P068P009P037nsss(0) <='0';
          end if;
        if(cVar1S30S117P066P018N049P067(0)='1' AND  A(11)='0' AND E( 8)='1' )then
          cVar2S30S117P016P069nsss(0) <='1';
          else
          cVar2S30S117P016P069nsss(0) <='0';
          end if;
        if(cVar1S31S117P066P018N049P067(0)='1' AND  A(11)='0' AND E( 8)='0' AND A( 4)='1' )then
          cVar2S31S117P016N069P011nsss(0) <='1';
          else
          cVar2S31S117P016N069P011nsss(0) <='0';
          end if;
        if(cVar1S32S117P066P018N049P067(0)='1' AND  A(11)='1' AND D(10)='1' AND A( 2)='1' )then
          cVar2S32S117P016P059P015nsss(0) <='1';
          else
          cVar2S32S117P016P059P015nsss(0) <='0';
          end if;
        if(cVar1S33S117P066P018N049P067(0)='1' AND  A(11)='1' AND B(14)='0' AND B( 9)='0' )then
          cVar2S33S117P016P026P036nsss(0) <='1';
          else
          cVar2S33S117P016P026P036nsss(0) <='0';
          end if;
        if(cVar1S34S117P066P018N049P067(0)='1' AND  A(11)='0' AND B(10)='0' AND D( 5)='1' )then
          cVar2S34S117N016P034P046nsss(0) <='1';
          else
          cVar2S34S117N016P034P046nsss(0) <='0';
          end if;
        if(cVar1S35S117P066P018N049P067(0)='1' AND  A(11)='0' AND B(10)='1' AND A( 0)='1' )then
          cVar2S35S117N016P034P019nsss(0) <='1';
          else
          cVar2S35S117N016P034P019nsss(0) <='0';
          end if;
        if(cVar1S0S118P035P033P002P048(0)='1' AND  E( 1)='0' AND D( 9)='0' )then
          cVar2S0S118P064P063nsss(0) <='1';
          else
          cVar2S0S118P064P063nsss(0) <='0';
          end if;
        if(cVar1S1S118P035P033P002N048(0)='1' AND  A(16)='0' AND E(10)='0' AND D( 6)='0' )then
          cVar2S1S118P006P061P042nsss(0) <='1';
          else
          cVar2S1S118P006P061P042nsss(0) <='0';
          end if;
        if(cVar1S2S118P035P033P002N048(0)='1' AND  A(16)='0' AND E(10)='1' AND E( 2)='0' )then
          cVar2S2S118P006P061P060nsss(0) <='1';
          else
          cVar2S2S118P006P061P060nsss(0) <='0';
          end if;
        if(cVar1S3S118P035P033P002N048(0)='1' AND  A(16)='1' AND A( 1)='0' AND A( 2)='1' )then
          cVar2S3S118P006P017P015nsss(0) <='1';
          else
          cVar2S3S118P006P017P015nsss(0) <='0';
          end if;
        if(cVar1S4S118P035P033P002P018(0)='1' AND  A(11)='0' AND A( 1)='0' )then
          cVar2S4S118P016P017nsss(0) <='1';
          else
          cVar2S4S118P016P017nsss(0) <='0';
          end if;
        if(cVar1S5S118P035P033P002N018(0)='1' AND  A( 4)='1' )then
          cVar2S5S118P011nsss(0) <='1';
          else
          cVar2S5S118P011nsss(0) <='0';
          end if;
        if(cVar1S6S118P035P033P002N018(0)='1' AND  A( 4)='0' AND A( 3)='1' )then
          cVar2S6S118N011P013nsss(0) <='1';
          else
          cVar2S6S118N011P013nsss(0) <='0';
          end if;
        if(cVar1S7S118P035N033P019P069(0)='1' AND  E( 0)='0' AND B( 9)='0' )then
          cVar2S7S118P068P036nsss(0) <='1';
          else
          cVar2S7S118P068P036nsss(0) <='0';
          end if;
        if(cVar1S8S118P035N033P019P069(0)='1' AND  E( 0)='0' AND B( 9)='1' AND D( 6)='1' )then
          cVar2S8S118P068P036P042nsss(0) <='1';
          else
          cVar2S8S118P068P036P042nsss(0) <='0';
          end if;
        if(cVar1S9S118P035N033P019P069(0)='1' AND  E( 0)='1' AND A(10)='1' AND A( 1)='1' )then
          cVar2S9S118P068P018P017nsss(0) <='1';
          else
          cVar2S9S118P068P018P017nsss(0) <='0';
          end if;
        if(cVar1S10S118P035N033P019P069(0)='1' AND  E( 0)='1' AND A(10)='0' AND D(11)='1' )then
          cVar2S10S118P068N018P055nsss(0) <='1';
          else
          cVar2S10S118P068N018P055nsss(0) <='0';
          end if;
        if(cVar1S11S118P035N033P019P069(0)='1' AND  D( 0)='1' AND B(10)='0' )then
          cVar2S11S118P066P034nsss(0) <='1';
          else
          cVar2S11S118P066P034nsss(0) <='0';
          end if;
        if(cVar1S12S118P035N033P019P069(0)='1' AND  D( 0)='1' AND B(10)='1' AND A(13)='1' )then
          cVar2S12S118P066P034P012nsss(0) <='1';
          else
          cVar2S12S118P066P034P012nsss(0) <='0';
          end if;
        if(cVar1S13S118P035N033P019P069(0)='1' AND  D( 0)='0' AND B(12)='1' AND A(10)='1' )then
          cVar2S13S118N066P030P018nsss(0) <='1';
          else
          cVar2S13S118N066P030P018nsss(0) <='0';
          end if;
        if(cVar1S14S118P035N033P019P018(0)='1' AND  E( 5)='0' AND B( 4)='1' )then
          cVar2S14S118P048P029nsss(0) <='1';
          else
          cVar2S14S118P048P029nsss(0) <='0';
          end if;
        if(cVar1S15S118P035N033P019P018(0)='1' AND  E( 5)='0' AND B( 4)='0' AND A( 4)='0' )then
          cVar2S15S118P048N029P011nsss(0) <='1';
          else
          cVar2S15S118P048N029P011nsss(0) <='0';
          end if;
        if(cVar1S16S118P035N033P019P018(0)='1' AND  E( 5)='1' AND B( 6)='1' )then
          cVar2S16S118P048P025nsss(0) <='1';
          else
          cVar2S16S118P048P025nsss(0) <='0';
          end if;
        if(cVar1S17S118P035N033P019N018(0)='1' AND  E( 5)='1' AND D( 0)='0' AND B( 0)='0' )then
          cVar2S17S118P048P066P037nsss(0) <='1';
          else
          cVar2S17S118P048P066P037nsss(0) <='0';
          end if;
        if(cVar1S18S118P035N033P019N018(0)='1' AND  E( 5)='1' AND D( 0)='1' AND B(14)='1' )then
          cVar2S18S118P048P066P026nsss(0) <='1';
          else
          cVar2S18S118P048P066P026nsss(0) <='0';
          end if;
        if(cVar1S19S118P035N033P019N018(0)='1' AND  E( 5)='0' AND E(14)='1' )then
          cVar2S19S118N048P045nsss(0) <='1';
          else
          cVar2S19S118N048P045nsss(0) <='0';
          end if;
        if(cVar1S20S118P035N033P019N018(0)='1' AND  E( 5)='0' AND E(14)='0' AND D( 1)='1' )then
          cVar2S20S118N048N045P062nsss(0) <='1';
          else
          cVar2S20S118N048N045P062nsss(0) <='0';
          end if;
        if(cVar1S21S118P035P046P058P033(0)='1' AND  D( 9)='1' )then
          cVar2S21S118P063nsss(0) <='1';
          else
          cVar2S21S118P063nsss(0) <='0';
          end if;
        if(cVar1S22S118P035P046P058P033(0)='1' AND  D( 9)='0' AND A( 0)='0' )then
          cVar2S22S118N063P019nsss(0) <='1';
          else
          cVar2S22S118N063P019nsss(0) <='0';
          end if;
        if(cVar1S23S118P035N046P022P034(0)='1' AND  A(16)='0' AND E( 9)='1' )then
          cVar2S23S118P006P065nsss(0) <='1';
          else
          cVar2S23S118P006P065nsss(0) <='0';
          end if;
        if(cVar1S24S118P035N046P022P034(0)='1' AND  A(16)='1' AND B(13)='1' )then
          cVar2S24S118P006P028nsss(0) <='1';
          else
          cVar2S24S118P006P028nsss(0) <='0';
          end if;
        if(cVar1S25S118P035N046P022P034(0)='1' AND  A(16)='1' AND B(13)='0' AND E( 3)='1' )then
          cVar2S25S118P006N028P056nsss(0) <='1';
          else
          cVar2S25S118P006N028P056nsss(0) <='0';
          end if;
        if(cVar1S26S118P035N046P022P034(0)='1' AND  A(15)='0' AND B( 2)='1' AND B( 9)='0' )then
          cVar2S26S118P008P033P036nsss(0) <='1';
          else
          cVar2S26S118P008P033P036nsss(0) <='0';
          end if;
        if(cVar1S27S118P035N046P022P034(0)='1' AND  A(15)='0' AND B( 2)='0' AND A( 7)='1' )then
          cVar2S27S118P008N033P005nsss(0) <='1';
          else
          cVar2S27S118P008N033P005nsss(0) <='0';
          end if;
        if(cVar1S28S118P035N046P022P034(0)='1' AND  A(15)='1' AND E( 2)='0' AND B( 9)='1' )then
          cVar2S28S118P008P060P036nsss(0) <='1';
          else
          cVar2S28S118P008P060P036nsss(0) <='0';
          end if;
        if(cVar1S30S118P035N046P022N065(0)='1' AND  A( 3)='1' )then
          cVar2S30S118P013nsss(0) <='1';
          else
          cVar2S30S118P013nsss(0) <='0';
          end if;
        if(cVar1S31S118P035N046P022N065(0)='1' AND  A( 3)='0' AND A(16)='1' )then
          cVar2S31S118N013P006nsss(0) <='1';
          else
          cVar2S31S118N013P006nsss(0) <='0';
          end if;
        if(cVar1S0S119P065P027P010P032(0)='1' AND  A( 9)='0' AND B(14)='0' )then
          cVar2S0S119P001P026nsss(0) <='1';
          else
          cVar2S0S119P001P026nsss(0) <='0';
          end if;
        if(cVar1S1S119P065P027P010P032(0)='1' AND  A( 9)='0' AND B(14)='1' AND D( 8)='0' )then
          cVar2S1S119P001P026P067nsss(0) <='1';
          else
          cVar2S1S119P001P026P067nsss(0) <='0';
          end if;
        if(cVar1S2S119P065P027P010P032(0)='1' AND  E( 4)='0' AND E(10)='1' )then
          cVar2S2S119P052P061nsss(0) <='1';
          else
          cVar2S2S119P052P061nsss(0) <='0';
          end if;
        if(cVar1S3S119P065P027P010P031(0)='1' AND  B( 9)='1' AND A(10)='0' )then
          cVar2S3S119P036P018nsss(0) <='1';
          else
          cVar2S3S119P036P018nsss(0) <='0';
          end if;
        if(cVar1S4S119P065P027P010P031(0)='1' AND  B( 9)='0' AND D( 4)='1' AND A( 0)='1' )then
          cVar2S4S119N036P050P019nsss(0) <='1';
          else
          cVar2S4S119N036P050P019nsss(0) <='0';
          end if;
        if(cVar1S5S119P065P027P010P031(0)='1' AND  B( 9)='0' AND D( 4)='0' AND A( 4)='1' )then
          cVar2S5S119N036N050P011nsss(0) <='1';
          else
          cVar2S5S119N036N050P011nsss(0) <='0';
          end if;
        if(cVar1S6S119P065N027P037P016(0)='1' AND  B(10)='1' AND A( 0)='0' AND B(12)='0' )then
          cVar2S6S119P034P019P030nsss(0) <='1';
          else
          cVar2S6S119P034P019P030nsss(0) <='0';
          end if;
        if(cVar1S7S119P065N027P037P016(0)='1' AND  B(10)='0' AND E( 8)='1' AND D( 0)='0' )then
          cVar2S7S119N034P069P066nsss(0) <='1';
          else
          cVar2S7S119N034P069P066nsss(0) <='0';
          end if;
        if(cVar1S8S119P065N027P037P016(0)='1' AND  B(10)='0' AND E( 8)='0' AND D( 4)='0' )then
          cVar2S8S119N034N069P050nsss(0) <='1';
          else
          cVar2S8S119N034N069P050nsss(0) <='0';
          end if;
        if(cVar1S9S119P065N027P037N016(0)='1' AND  B( 9)='0' AND E( 0)='1' AND A(15)='0' )then
          cVar2S9S119P036P068P008nsss(0) <='1';
          else
          cVar2S9S119P036P068P008nsss(0) <='0';
          end if;
        if(cVar1S10S119P065N027P037N016(0)='1' AND  B( 9)='0' AND E( 0)='0' AND D( 0)='0' )then
          cVar2S10S119P036N068P066nsss(0) <='1';
          else
          cVar2S10S119P036N068P066nsss(0) <='0';
          end if;
        if(cVar1S11S119P065N027P037N016(0)='1' AND  B( 9)='1' AND E(12)='0' AND B(16)='1' )then
          cVar2S11S119P036P053P022nsss(0) <='1';
          else
          cVar2S11S119P036P053P022nsss(0) <='0';
          end if;
        if(cVar1S12S119P065N027P037P008(0)='1' AND  B(15)='1' AND D(13)='1' )then
          cVar2S12S119P024P047nsss(0) <='1';
          else
          cVar2S12S119P024P047nsss(0) <='0';
          end if;
        if(cVar1S13S119P065N027P037P008(0)='1' AND  B(15)='1' AND D(13)='0' AND A( 1)='1' )then
          cVar2S13S119P024N047P017nsss(0) <='1';
          else
          cVar2S13S119P024N047P017nsss(0) <='0';
          end if;
        if(cVar1S14S119P065N027P037P008(0)='1' AND  B(15)='0' AND E( 4)='1' )then
          cVar2S14S119N024P052nsss(0) <='1';
          else
          cVar2S14S119N024P052nsss(0) <='0';
          end if;
        if(cVar1S15S119P065N027P037P008(0)='1' AND  B(15)='0' AND E( 4)='0' AND A( 3)='0' )then
          cVar2S15S119N024N052P013nsss(0) <='1';
          else
          cVar2S15S119N024N052P013nsss(0) <='0';
          end if;
        if(cVar1S16S119P065N027P037N008(0)='1' AND  E(11)='1' AND E(12)='0' )then
          cVar2S16S119P057P053nsss(0) <='1';
          else
          cVar2S16S119P057P053nsss(0) <='0';
          end if;
        if(cVar1S17S119P065N027P037N008(0)='1' AND  E(11)='0' AND A( 5)='1' AND E( 8)='1' )then
          cVar2S17S119N057P009P069nsss(0) <='1';
          else
          cVar2S17S119N057P009P069nsss(0) <='0';
          end if;
        if(cVar1S18S119P065P008P064P069(0)='1' AND  E( 2)='0' AND D( 0)='0' )then
          cVar2S18S119P060P066nsss(0) <='1';
          else
          cVar2S18S119P060P066nsss(0) <='0';
          end if;
        if(cVar1S19S119P065P008P064P069(0)='1' AND  E( 2)='0' AND D( 0)='1' AND E(12)='0' )then
          cVar2S19S119P060P066P053nsss(0) <='1';
          else
          cVar2S19S119P060P066P053nsss(0) <='0';
          end if;
        if(cVar1S20S119P065P008P064P069(0)='1' AND  E( 2)='1' AND E(11)='0' AND A( 1)='1' )then
          cVar2S20S119P060P057P017nsss(0) <='1';
          else
          cVar2S20S119P060P057P017nsss(0) <='0';
          end if;
        if(cVar1S21S119P065P008P064P069(0)='1' AND  D(10)='0' AND A(10)='1' AND A( 0)='1' )then
          cVar2S21S119P059P018P019nsss(0) <='1';
          else
          cVar2S21S119P059P018P019nsss(0) <='0';
          end if;
        if(cVar1S22S119P065P008P064P069(0)='1' AND  D(10)='1' AND B( 0)='1' )then
          cVar2S22S119P059P037nsss(0) <='1';
          else
          cVar2S22S119P059P037nsss(0) <='0';
          end if;
        if(cVar1S23S119P065P008P064P014(0)='1' AND  B( 1)='0' AND B(10)='0' AND A( 3)='0' )then
          cVar2S23S119P035P034P013nsss(0) <='1';
          else
          cVar2S23S119P035P034P013nsss(0) <='0';
          end if;
        if(cVar1S24S119P065P008P064P014(0)='1' AND  B( 1)='0' AND B(10)='1' AND A( 1)='0' )then
          cVar2S24S119P035P034P017nsss(0) <='1';
          else
          cVar2S24S119P035P034P017nsss(0) <='0';
          end if;
        if(cVar1S25S119P065P008P064P014(0)='1' AND  B( 1)='1' AND A( 5)='0' AND D( 0)='1' )then
          cVar2S25S119P035P009P066nsss(0) <='1';
          else
          cVar2S25S119P035P009P066nsss(0) <='0';
          end if;
        if(cVar1S26S119P065P008P064N014(0)='1' AND  D( 9)='0' AND D( 8)='0' AND B( 1)='1' )then
          cVar2S26S119P063P067P035nsss(0) <='1';
          else
          cVar2S26S119P063P067P035nsss(0) <='0';
          end if;
        if(cVar1S27S119P065P008P064N014(0)='1' AND  D( 9)='0' AND D( 8)='1' AND A(10)='0' )then
          cVar2S27S119P063P067P018nsss(0) <='1';
          else
          cVar2S27S119P063P067P018nsss(0) <='0';
          end if;
        if(cVar1S28S119P065P008P064N014(0)='1' AND  D( 9)='1' AND E( 8)='1' AND A( 0)='0' )then
          cVar2S28S119P063P069P019nsss(0) <='1';
          else
          cVar2S28S119P063P069P019nsss(0) <='0';
          end if;
        if(cVar1S29S119P065P008P064N014(0)='1' AND  D( 9)='1' AND E( 8)='0' AND A(17)='1' )then
          cVar2S29S119P063N069P004nsss(0) <='1';
          else
          cVar2S29S119P063N069P004nsss(0) <='0';
          end if;
        if(cVar1S30S119P065P008P011P014(0)='1' AND  D( 9)='1' AND B( 9)='1' )then
          cVar2S30S119P063P036nsss(0) <='1';
          else
          cVar2S30S119P063P036nsss(0) <='0';
          end if;
        if(cVar1S31S119P065P008P011P014(0)='1' AND  D( 9)='1' AND B( 9)='0' AND B(10)='1' )then
          cVar2S31S119P063N036P034nsss(0) <='1';
          else
          cVar2S31S119P063N036P034nsss(0) <='0';
          end if;
        if(cVar1S32S119P065P008P011P014(0)='1' AND  D( 0)='0' AND A( 0)='0' )then
          cVar2S32S119P066P019nsss(0) <='1';
          else
          cVar2S32S119P066P019nsss(0) <='0';
          end if;
        if(cVar1S34S119P065P008N011N056(0)='1' AND  A( 0)='1' AND A( 2)='0' AND D( 8)='0' )then
          cVar2S34S119P019P015P067nsss(0) <='1';
          else
          cVar2S34S119P019P015P067nsss(0) <='0';
          end if;
        if(cVar1S35S119P065P008N011N056(0)='1' AND  A( 0)='0' AND D( 2)='1' )then
          cVar2S35S119N019P058nsss(0) <='1';
          else
          cVar2S35S119N019P058nsss(0) <='0';
          end if;
        if(cVar1S0S120P037P001P032P018(0)='1' AND  A( 1)='0' AND A( 0)='0' )then
          cVar2S0S120P017P019nsss(0) <='1';
          else
          cVar2S0S120P017P019nsss(0) <='0';
          end if;
        if(cVar1S1S120P037P001P032P018(0)='1' AND  A( 1)='0' AND A( 0)='1' AND A( 3)='1' )then
          cVar2S1S120P017P019P013nsss(0) <='1';
          else
          cVar2S1S120P017P019P013nsss(0) <='0';
          end if;
        if(cVar1S2S120P037P001P032P018(0)='1' AND  A( 1)='1' AND E( 2)='1' )then
          cVar2S2S120P017P060nsss(0) <='1';
          else
          cVar2S2S120P017P060nsss(0) <='0';
          end if;
        if(cVar1S3S120P037P001P032P018(0)='1' AND  A( 1)='1' AND E( 2)='0' AND B(10)='1' )then
          cVar2S3S120P017N060P034nsss(0) <='1';
          else
          cVar2S3S120P017N060P034nsss(0) <='0';
          end if;
        if(cVar1S4S120P037P001P032N018(0)='1' AND  E( 0)='0' AND E( 3)='0' )then
          cVar2S4S120P068P056nsss(0) <='1';
          else
          cVar2S4S120P068P056nsss(0) <='0';
          end if;
        if(cVar1S5S120P037P001P032N018(0)='1' AND  E( 0)='1' AND B( 9)='0' AND E(10)='0' )then
          cVar2S5S120P068P036P061nsss(0) <='1';
          else
          cVar2S5S120P068P036P061nsss(0) <='0';
          end if;
        if(cVar1S6S120P037P001N032P056(0)='1' AND  A(10)='0' AND E( 8)='1' AND B( 9)='0' )then
          cVar2S6S120P018P069P036nsss(0) <='1';
          else
          cVar2S6S120P018P069P036nsss(0) <='0';
          end if;
        if(cVar1S7S120P037P001N032P056(0)='1' AND  A(10)='0' AND E( 8)='0' )then
          cVar2S7S120P018N069psss(0) <='1';
          else
          cVar2S7S120P018N069psss(0) <='0';
          end if;
        if(cVar1S8S120P037P001N032P056(0)='1' AND  A(10)='1' AND A( 1)='0' )then
          cVar2S8S120P018P017nsss(0) <='1';
          else
          cVar2S8S120P018P017nsss(0) <='0';
          end if;
        if(cVar1S9S120P037P001N032P056(0)='1' AND  A(10)='1' AND A( 1)='1' AND B( 1)='1' )then
          cVar2S9S120P018P017P035nsss(0) <='1';
          else
          cVar2S9S120P018P017P035nsss(0) <='0';
          end if;
        if(cVar1S10S120P037P001N032N056(0)='1' AND  E( 4)='1' )then
          cVar2S10S120P052nsss(0) <='1';
          else
          cVar2S10S120P052nsss(0) <='0';
          end if;
        if(cVar1S11S120P037P001N032N056(0)='1' AND  E( 4)='0' AND B( 3)='0' )then
          cVar2S11S120N052P031nsss(0) <='1';
          else
          cVar2S11S120N052P031nsss(0) <='0';
          end if;
        if(cVar1S12S120P037P001N032N056(0)='1' AND  E( 4)='0' AND B( 3)='1' AND A( 3)='1' )then
          cVar2S12S120N052P031P013nsss(0) <='1';
          else
          cVar2S12S120N052P031P013nsss(0) <='0';
          end if;
        if(cVar1S13S120P037P001P036P019(0)='1' AND  A(11)='0' AND E( 0)='1' )then
          cVar2S13S120P016P068nsss(0) <='1';
          else
          cVar2S13S120P016P068nsss(0) <='0';
          end if;
        if(cVar1S14S120P037P001P036P019(0)='1' AND  A(11)='0' AND E( 0)='0' AND A(10)='0' )then
          cVar2S14S120P016N068P018nsss(0) <='1';
          else
          cVar2S14S120P016N068P018nsss(0) <='0';
          end if;
        if(cVar1S15S120P037P001P036P019(0)='1' AND  A(11)='1' AND A(12)='1' )then
          cVar2S15S120P016P014nsss(0) <='1';
          else
          cVar2S15S120P016P014nsss(0) <='0';
          end if;
        if(cVar1S16S120P037P001P036N019(0)='1' AND  A(12)='1' AND A( 1)='1' )then
          cVar2S16S120P014P017nsss(0) <='1';
          else
          cVar2S16S120P014P017nsss(0) <='0';
          end if;
        if(cVar1S17S120P037P001P036P008(0)='1' AND  A(10)='1' AND A(11)='0' )then
          cVar2S17S120P018P016nsss(0) <='1';
          else
          cVar2S17S120P018P016nsss(0) <='0';
          end if;
        if(cVar1S18S120N037P036P065P017(0)='1' AND  B( 5)='1' )then
          cVar2S18S120P027nsss(0) <='1';
          else
          cVar2S18S120P027nsss(0) <='0';
          end if;
        if(cVar1S19S120N037P036P065P017(0)='1' AND  B( 5)='0' AND A(14)='0' AND B(11)='0' )then
          cVar2S19S120N027P010P032nsss(0) <='1';
          else
          cVar2S19S120N027P010P032nsss(0) <='0';
          end if;
        if(cVar1S20S120N037P036P065P017(0)='1' AND  B( 5)='0' AND A(14)='1' AND E( 3)='1' )then
          cVar2S20S120N027P010P056nsss(0) <='1';
          else
          cVar2S20S120N027P010P056nsss(0) <='0';
          end if;
        if(cVar1S21S120N037P036P065N017(0)='1' AND  E( 3)='1' AND A( 8)='0' AND B( 4)='0' )then
          cVar2S21S120P056P003P029nsss(0) <='1';
          else
          cVar2S21S120P056P003P029nsss(0) <='0';
          end if;
        if(cVar1S22S120N037P036P065N017(0)='1' AND  E( 3)='0' AND A(13)='0' )then
          cVar2S22S120N056P012nsss(0) <='1';
          else
          cVar2S22S120N056P012nsss(0) <='0';
          end if;
        if(cVar1S23S120N037P036P065N017(0)='1' AND  E( 3)='0' AND A(13)='1' AND E( 2)='1' )then
          cVar2S23S120N056P012P060nsss(0) <='1';
          else
          cVar2S23S120N056P012P060nsss(0) <='0';
          end if;
        if(cVar1S24S120N037P036P065P016(0)='1' AND  E( 5)='1' )then
          cVar2S24S120P048nsss(0) <='1';
          else
          cVar2S24S120P048nsss(0) <='0';
          end if;
        if(cVar1S25S120N037P036P065P016(0)='1' AND  E( 5)='0' AND E( 0)='0' AND A(10)='1' )then
          cVar2S25S120N048P068P018nsss(0) <='1';
          else
          cVar2S25S120N048P068P018nsss(0) <='0';
          end if;
        if(cVar1S26S120N037P036P065P016(0)='1' AND  B(15)='0' AND B(11)='1' )then
          cVar2S26S120P024P032nsss(0) <='1';
          else
          cVar2S26S120P024P032nsss(0) <='0';
          end if;
        if(cVar1S27S120N037N036P034P050(0)='1' AND  E(10)='1' AND A( 0)='1' )then
          cVar2S27S120P061P019nsss(0) <='1';
          else
          cVar2S27S120P061P019nsss(0) <='0';
          end if;
        if(cVar1S28S120N037N036P034P050(0)='1' AND  E(10)='1' AND A( 0)='0' AND D( 8)='0' )then
          cVar2S28S120P061N019P067nsss(0) <='1';
          else
          cVar2S28S120P061N019P067nsss(0) <='0';
          end if;
        if(cVar1S29S120N037N036P034P050(0)='1' AND  E(10)='0' AND D(10)='0' AND B( 6)='0' )then
          cVar2S29S120N061P059P025nsss(0) <='1';
          else
          cVar2S29S120N061P059P025nsss(0) <='0';
          end if;
        if(cVar1S30S120N037N036P034P050(0)='1' AND  E(10)='0' AND D(10)='1' AND E( 1)='1' )then
          cVar2S30S120N061P059P064nsss(0) <='1';
          else
          cVar2S30S120N061P059P064nsss(0) <='0';
          end if;
        if(cVar1S31S120N037N036P034P050(0)='1' AND  A( 1)='1' AND A( 0)='0' )then
          cVar2S31S120P017P019nsss(0) <='1';
          else
          cVar2S31S120P017P019nsss(0) <='0';
          end if;
        if(cVar1S32S120N037N036P034P050(0)='1' AND  A( 1)='0' AND B( 5)='1' )then
          cVar2S32S120N017P027nsss(0) <='1';
          else
          cVar2S32S120N017P027nsss(0) <='0';
          end if;
        if(cVar1S33S120N037N036N034P065(0)='1' AND  A( 1)='0' AND D( 9)='1' AND E(11)='1' )then
          cVar2S33S120P017P063P057nsss(0) <='1';
          else
          cVar2S33S120P017P063P057nsss(0) <='0';
          end if;
        if(cVar1S34S120N037N036N034P065(0)='1' AND  A( 1)='1' AND E(10)='1' AND D(11)='0' )then
          cVar2S34S120P017P061P055nsss(0) <='1';
          else
          cVar2S34S120P017P061P055nsss(0) <='0';
          end if;
        if(cVar1S35S120N037N036N034P065(0)='1' AND  A( 1)='1' AND E(10)='0' AND B( 4)='1' )then
          cVar2S35S120P017N061P029nsss(0) <='1';
          else
          cVar2S35S120P017N061P029nsss(0) <='0';
          end if;
        if(cVar1S36S120N037N036N034P065(0)='1' AND  B( 1)='1' AND A( 6)='0' )then
          cVar2S36S120P035P007nsss(0) <='1';
          else
          cVar2S36S120P035P007nsss(0) <='0';
          end if;
        if(cVar1S37S120N037N036N034P065(0)='1' AND  B( 1)='0' AND D( 9)='0' AND A( 4)='1' )then
          cVar2S37S120N035P063P011nsss(0) <='1';
          else
          cVar2S37S120N035P063P011nsss(0) <='0';
          end if;
        if(cVar1S0S121P065P052P034P009(0)='1' AND  E( 3)='1' )then
          cVar2S0S121P056nsss(0) <='1';
          else
          cVar2S0S121P056nsss(0) <='0';
          end if;
        if(cVar1S1S121P065P052P034P009(0)='1' AND  E( 3)='0' AND A(15)='1' )then
          cVar2S1S121N056P008nsss(0) <='1';
          else
          cVar2S1S121N056P008nsss(0) <='0';
          end if;
        if(cVar1S2S121P065P052P034P009(0)='1' AND  E( 3)='0' AND A(15)='0' AND A( 0)='1' )then
          cVar2S2S121N056N008P019nsss(0) <='1';
          else
          cVar2S2S121N056N008P019nsss(0) <='0';
          end if;
        if(cVar1S3S121P065P052P034N009(0)='1' AND  E( 3)='0' AND E( 5)='0' AND D( 5)='0' )then
          cVar2S3S121P056P048P046nsss(0) <='1';
          else
          cVar2S3S121P056P048P046nsss(0) <='0';
          end if;
        if(cVar1S4S121P065P052P034N009(0)='1' AND  E( 3)='1' AND A( 2)='1' )then
          cVar2S4S121P056P015nsss(0) <='1';
          else
          cVar2S4S121P056P015nsss(0) <='0';
          end if;
        if(cVar1S5S121P065P052P034P011(0)='1' AND  A(12)='1' )then
          cVar2S5S121P014nsss(0) <='1';
          else
          cVar2S5S121P014nsss(0) <='0';
          end if;
        if(cVar1S6S121P065P052P034N011(0)='1' AND  A( 2)='0' AND D( 1)='0' AND D( 4)='0' )then
          cVar2S6S121P015P062P050nsss(0) <='1';
          else
          cVar2S6S121P015P062P050nsss(0) <='0';
          end if;
        if(cVar1S7S121P065N052P050P046(0)='1' AND  A(17)='1' AND B( 6)='1' )then
          cVar2S7S121P004P025nsss(0) <='1';
          else
          cVar2S7S121P004P025nsss(0) <='0';
          end if;
        if(cVar1S8S121P065N052P050P046(0)='1' AND  A(17)='1' AND B( 6)='0' AND A( 2)='1' )then
          cVar2S8S121P004N025P015nsss(0) <='1';
          else
          cVar2S8S121P004N025P015nsss(0) <='0';
          end if;
        if(cVar1S9S121P065N052P050P046(0)='1' AND  A(17)='0' AND B( 5)='1' )then
          cVar2S9S121N004P027nsss(0) <='1';
          else
          cVar2S9S121N004P027nsss(0) <='0';
          end if;
        if(cVar1S10S121P065N052P050N046(0)='1' AND  D(12)='1' AND A( 5)='1' AND D(11)='0' )then
          cVar2S10S121P051P009P055nsss(0) <='1';
          else
          cVar2S10S121P051P009P055nsss(0) <='0';
          end if;
        if(cVar1S11S121P065N052P050N046(0)='1' AND  D(12)='1' AND A( 5)='0' AND A( 7)='0' )then
          cVar2S11S121P051N009P005nsss(0) <='1';
          else
          cVar2S11S121P051N009P005nsss(0) <='0';
          end if;
        if(cVar1S12S121P065N052P050N046(0)='1' AND  D(12)='0' AND B( 5)='0' AND A(15)='0' )then
          cVar2S12S121N051P027P008nsss(0) <='1';
          else
          cVar2S12S121N051P027P008nsss(0) <='0';
          end if;
        if(cVar1S13S121P065N052P050P060(0)='1' AND  D( 8)='1' )then
          cVar2S13S121P067nsss(0) <='1';
          else
          cVar2S13S121P067nsss(0) <='0';
          end if;
        if(cVar1S14S121P065N052P050P060(0)='1' AND  D( 8)='0' AND A(11)='1' )then
          cVar2S14S121N067P016nsss(0) <='1';
          else
          cVar2S14S121N067P016nsss(0) <='0';
          end if;
        if(cVar1S15S121P065N052P050P060(0)='1' AND  D( 8)='0' AND A(11)='0' AND E( 5)='1' )then
          cVar2S15S121N067N016P048nsss(0) <='1';
          else
          cVar2S15S121N067N016P048nsss(0) <='0';
          end if;
        if(cVar1S16S121P065N052P050N060(0)='1' AND  E( 5)='1' AND D( 5)='0' AND A(10)='0' )then
          cVar2S16S121P048P046P018nsss(0) <='1';
          else
          cVar2S16S121P048P046P018nsss(0) <='0';
          end if;
        if(cVar1S17S121P065N052P050N060(0)='1' AND  E( 5)='0' AND D( 8)='1' AND B( 0)='1' )then
          cVar2S17S121N048P067P037nsss(0) <='1';
          else
          cVar2S17S121N048P067P037nsss(0) <='0';
          end if;
        if(cVar1S18S121P065N052P050N060(0)='1' AND  E( 5)='0' AND D( 8)='0' AND D(10)='1' )then
          cVar2S18S121N048N067P059nsss(0) <='1';
          else
          cVar2S18S121N048N067P059nsss(0) <='0';
          end if;
        if(cVar1S19S121P065P036P024P030(0)='1' AND  A( 2)='0' )then
          cVar2S19S121P015nsss(0) <='1';
          else
          cVar2S19S121P015nsss(0) <='0';
          end if;
        if(cVar1S20S121P065P036P024N030(0)='1' AND  D( 0)='0' AND A(11)='0' )then
          cVar2S20S121P066P016nsss(0) <='1';
          else
          cVar2S20S121P066P016nsss(0) <='0';
          end if;
        if(cVar1S21S121P065P036P024N030(0)='1' AND  D( 0)='0' AND A(11)='1' AND B(11)='1' )then
          cVar2S21S121P066P016P032nsss(0) <='1';
          else
          cVar2S21S121P066P016P032nsss(0) <='0';
          end if;
        if(cVar1S22S121P065P036P024N030(0)='1' AND  D( 0)='1' AND A( 3)='1' AND A(13)='0' )then
          cVar2S22S121P066P013P012nsss(0) <='1';
          else
          cVar2S22S121P066P013P012nsss(0) <='0';
          end if;
        if(cVar1S23S121P065P036P024N030(0)='1' AND  D( 0)='1' AND A( 3)='0' AND A(12)='1' )then
          cVar2S23S121P066N013P014nsss(0) <='1';
          else
          cVar2S23S121P066N013P014nsss(0) <='0';
          end if;
        if(cVar1S24S121P065P036P024P034(0)='1' AND  D( 8)='0' AND A( 0)='1' )then
          cVar2S24S121P067P019nsss(0) <='1';
          else
          cVar2S24S121P067P019nsss(0) <='0';
          end if;
        if(cVar1S25S121P065N036P008P041(0)='1' AND  E( 2)='1' AND B(11)='1' )then
          cVar2S25S121P060P032nsss(0) <='1';
          else
          cVar2S25S121P060P032nsss(0) <='0';
          end if;
        if(cVar1S26S121P065N036P008P041(0)='1' AND  E( 2)='1' AND B(11)='0' AND A( 6)='1' )then
          cVar2S26S121P060N032P007nsss(0) <='1';
          else
          cVar2S26S121P060N032P007nsss(0) <='0';
          end if;
        if(cVar1S27S121P065N036P008P041(0)='1' AND  E( 2)='0' AND B(11)='0' AND E(14)='1' )then
          cVar2S27S121N060P032P045nsss(0) <='1';
          else
          cVar2S27S121N060P032P045nsss(0) <='0';
          end if;
        if(cVar1S28S121P065N036P008P041(0)='1' AND  D(15)='1' )then
          cVar2S28S121P039nsss(0) <='1';
          else
          cVar2S28S121P039nsss(0) <='0';
          end if;
        if(cVar1S29S121P065N036P008P037(0)='1' AND  D( 1)='1' )then
          cVar2S29S121P062nsss(0) <='1';
          else
          cVar2S29S121P062nsss(0) <='0';
          end if;
        if(cVar1S30S121P065N036P008P037(0)='1' AND  D( 1)='0' AND A(10)='0' AND B(10)='0' )then
          cVar2S30S121N062P018P034nsss(0) <='1';
          else
          cVar2S30S121N062P018P034nsss(0) <='0';
          end if;
        if(cVar1S31S121P065N036P008N037(0)='1' AND  D( 9)='1' AND A( 4)='1' )then
          cVar2S31S121P063P011nsss(0) <='1';
          else
          cVar2S31S121P063P011nsss(0) <='0';
          end if;
        if(cVar1S32S121P065N036P008N037(0)='1' AND  D( 9)='1' AND A( 4)='0' AND E(12)='1' )then
          cVar2S32S121P063N011P053nsss(0) <='1';
          else
          cVar2S32S121P063N011P053nsss(0) <='0';
          end if;
        if(cVar1S1S122P052P009N056P010(0)='1' AND  B( 0)='0' )then
          cVar2S1S122P037nsss(0) <='1';
          else
          cVar2S1S122P037nsss(0) <='0';
          end if;
        if(cVar1S2S122P052P009N056N010(0)='1' AND  D( 4)='1' )then
          cVar2S2S122P050nsss(0) <='1';
          else
          cVar2S2S122P050nsss(0) <='0';
          end if;
        if(cVar1S3S122P052P009N056N010(0)='1' AND  D( 4)='0' AND A( 0)='1' )then
          cVar2S3S122N050P019nsss(0) <='1';
          else
          cVar2S3S122N050P019nsss(0) <='0';
          end if;
        if(cVar1S4S122P052N009P056P046(0)='1' AND  E(10)='0' AND E( 5)='0' AND B( 8)='0' )then
          cVar2S4S122P061P048P021nsss(0) <='1';
          else
          cVar2S4S122P061P048P021nsss(0) <='0';
          end if;
        if(cVar1S5S122P052N009P056P046(0)='1' AND  E(10)='0' AND E( 5)='1' AND A( 1)='1' )then
          cVar2S5S122P061P048P017nsss(0) <='1';
          else
          cVar2S5S122P061P048P017nsss(0) <='0';
          end if;
        if(cVar1S6S122P052N009P056P046(0)='1' AND  E(10)='1' AND D(10)='0' )then
          cVar2S6S122P061P059nsss(0) <='1';
          else
          cVar2S6S122P061P059nsss(0) <='0';
          end if;
        if(cVar1S7S122P052N009P056P046(0)='1' AND  E( 5)='1' )then
          cVar2S7S122P048nsss(0) <='1';
          else
          cVar2S7S122P048nsss(0) <='0';
          end if;
        if(cVar1S9S122P052N009P056N015(0)='1' AND  A(13)='1' )then
          cVar2S9S122P012nsss(0) <='1';
          else
          cVar2S9S122P012nsss(0) <='0';
          end if;
        if(cVar1S10S122N052P046P050P042(0)='1' AND  A(17)='1' AND B( 6)='1' )then
          cVar2S10S122P004P025nsss(0) <='1';
          else
          cVar2S10S122P004P025nsss(0) <='0';
          end if;
        if(cVar1S11S122N052P046P050P042(0)='1' AND  A(17)='1' AND B( 6)='0' AND A(11)='0' )then
          cVar2S11S122P004N025P016nsss(0) <='1';
          else
          cVar2S11S122P004N025P016nsss(0) <='0';
          end if;
        if(cVar1S12S122N052P046P050P042(0)='1' AND  A(17)='0' AND B( 5)='1' AND B( 6)='0' )then
          cVar2S12S122N004P027P025nsss(0) <='1';
          else
          cVar2S12S122N004P027P025nsss(0) <='0';
          end if;
        if(cVar1S13S122N052P046P050P042(0)='1' AND  A(17)='0' AND B( 5)='0' AND B( 1)='1' )then
          cVar2S13S122N004N027P035nsss(0) <='1';
          else
          cVar2S13S122N004N027P035nsss(0) <='0';
          end if;
        if(cVar1S14S122N052P046P050P042(0)='1' AND  A(11)='1' )then
          cVar2S14S122P016nsss(0) <='1';
          else
          cVar2S14S122P016nsss(0) <='0';
          end if;
        if(cVar1S16S122N052N046P065P008(0)='1' AND  E(15)='0' AND B( 9)='1' AND A( 0)='0' )then
          cVar2S16S122P041P036P019nsss(0) <='1';
          else
          cVar2S16S122P041P036P019nsss(0) <='0';
          end if;
        if(cVar1S17S122N052N046P065P008(0)='1' AND  E(15)='0' AND B( 9)='0' AND B( 1)='1' )then
          cVar2S17S122P041N036P035nsss(0) <='1';
          else
          cVar2S17S122P041N036P035nsss(0) <='0';
          end if;
        if(cVar1S18S122N052N046P065P008(0)='1' AND  E(15)='1' AND A( 7)='1' )then
          cVar2S18S122P041P005nsss(0) <='1';
          else
          cVar2S18S122P041P005nsss(0) <='0';
          end if;
        if(cVar1S19S122N052N046P065P008(0)='1' AND  A( 4)='1' AND B( 9)='1' AND D( 1)='0' )then
          cVar2S19S122P011P036P062nsss(0) <='1';
          else
          cVar2S19S122P011P036P062nsss(0) <='0';
          end if;
        if(cVar1S20S122N052N046P065P008(0)='1' AND  A( 4)='0' AND E( 3)='1' )then
          cVar2S20S122N011P056nsss(0) <='1';
          else
          cVar2S20S122N011P056nsss(0) <='0';
          end if;
        if(cVar1S21S122N052N046N065P049(0)='1' AND  A( 9)='0' AND A(10)='1' AND D(10)='0' )then
          cVar2S21S122P001P018P059nsss(0) <='1';
          else
          cVar2S21S122P001P018P059nsss(0) <='0';
          end if;
        if(cVar1S22S122N052N046N065P049(0)='1' AND  A( 9)='0' AND A(10)='0' AND A( 8)='1' )then
          cVar2S22S122P001N018P003nsss(0) <='1';
          else
          cVar2S22S122P001N018P003nsss(0) <='0';
          end if;
        if(cVar1S23S122N052N046N065N049(0)='1' AND  A( 6)='1' AND B( 4)='0' AND B(16)='1' )then
          cVar2S23S122P007P029P022nsss(0) <='1';
          else
          cVar2S23S122P007P029P022nsss(0) <='0';
          end if;
        if(cVar1S0S123P017P036P016P021(0)='1' AND  E( 6)='1' AND A( 2)='0' AND D( 0)='0' )then
          cVar2S0S123P044P015P066nsss(0) <='1';
          else
          cVar2S0S123P044P015P066nsss(0) <='0';
          end if;
        if(cVar1S1S123P017P036P016P021(0)='1' AND  E( 6)='1' AND A( 2)='1' AND A(10)='0' )then
          cVar2S1S123P044P015P018nsss(0) <='1';
          else
          cVar2S1S123P044P015P018nsss(0) <='0';
          end if;
        if(cVar1S2S123P017P036P016P021(0)='1' AND  E( 6)='0' AND D( 2)='1' AND A( 6)='0' )then
          cVar2S2S123N044P058P007nsss(0) <='1';
          else
          cVar2S2S123N044P058P007nsss(0) <='0';
          end if;
        if(cVar1S3S123P017P036P016P021(0)='1' AND  E( 6)='0' AND D( 2)='0' )then
          cVar2S3S123N044N058psss(0) <='1';
          else
          cVar2S3S123N044N058psss(0) <='0';
          end if;
        if(cVar1S4S123P017P036P016P021(0)='1' AND  A(17)='1' )then
          cVar2S4S123P004nsss(0) <='1';
          else
          cVar2S4S123P004nsss(0) <='0';
          end if;
        if(cVar1S5S123P017P036P016P021(0)='1' AND  A(17)='0' AND A( 8)='1' )then
          cVar2S5S123N004P003nsss(0) <='1';
          else
          cVar2S5S123N004P003nsss(0) <='0';
          end if;
        if(cVar1S6S123P017P036N016P034(0)='1' AND  E( 9)='0' AND D( 9)='0' )then
          cVar2S6S123P065P063nsss(0) <='1';
          else
          cVar2S6S123P065P063nsss(0) <='0';
          end if;
        if(cVar1S7S123P017P036N016P034(0)='1' AND  E( 9)='1' AND E( 8)='0' AND B( 1)='1' )then
          cVar2S7S123P065P069P035nsss(0) <='1';
          else
          cVar2S7S123P065P069P035nsss(0) <='0';
          end if;
        if(cVar1S8S123P017P036N016P034(0)='1' AND  E( 9)='1' AND E( 8)='1' AND E(11)='1' )then
          cVar2S8S123P065P069P057nsss(0) <='1';
          else
          cVar2S8S123P065P069P057nsss(0) <='0';
          end if;
        if(cVar1S9S123P017P036N016P034(0)='1' AND  B(12)='1' )then
          cVar2S9S123P030nsss(0) <='1';
          else
          cVar2S9S123P030nsss(0) <='0';
          end if;
        if(cVar1S10S123P017P036N016P034(0)='1' AND  B(12)='0' AND A( 2)='1' AND E( 8)='0' )then
          cVar2S10S123N030P015P069nsss(0) <='1';
          else
          cVar2S10S123N030P015P069nsss(0) <='0';
          end if;
        if(cVar1S11S123P017P036N016P034(0)='1' AND  B(12)='0' AND A( 2)='0' AND B( 2)='1' )then
          cVar2S11S123N030N015P033nsss(0) <='1';
          else
          cVar2S11S123N030N015P033nsss(0) <='0';
          end if;
        if(cVar1S12S123P017P036P056P052(0)='1' AND  A( 3)='0' AND B(11)='0' )then
          cVar2S12S123P013P032nsss(0) <='1';
          else
          cVar2S12S123P013P032nsss(0) <='0';
          end if;
        if(cVar1S13S123P017P036P056P052(0)='1' AND  A( 3)='1' AND A( 4)='1' AND B( 3)='1' )then
          cVar2S13S123P013P011P031nsss(0) <='1';
          else
          cVar2S13S123P013P011P031nsss(0) <='0';
          end if;
        if(cVar1S14S123P017P036P056P052(0)='1' AND  A( 3)='1' AND A( 4)='0' AND D( 3)='0' )then
          cVar2S14S123P013N011P054nsss(0) <='1';
          else
          cVar2S14S123P013N011P054nsss(0) <='0';
          end if;
        if(cVar1S15S123P017P036N056P065(0)='1' AND  A( 7)='0' )then
          cVar2S15S123P005nsss(0) <='1';
          else
          cVar2S15S123P005nsss(0) <='0';
          end if;
        if(cVar1S16S123P017P036N056P065(0)='1' AND  A( 7)='1' AND A(13)='1' )then
          cVar2S16S123P005P012nsss(0) <='1';
          else
          cVar2S16S123P005P012nsss(0) <='0';
          end if;
        if(cVar1S17S123P017P036N056N065(0)='1' AND  D(14)='1' )then
          cVar2S17S123P043nsss(0) <='1';
          else
          cVar2S17S123P043nsss(0) <='0';
          end if;
        if(cVar1S18S123P017P036P065P019(0)='1' AND  E( 1)='0' AND A(17)='1' AND A(12)='0' )then
          cVar2S18S123P064P004P014nsss(0) <='1';
          else
          cVar2S18S123P064P004P014nsss(0) <='0';
          end if;
        if(cVar1S19S123P017P036P065P019(0)='1' AND  E( 1)='0' AND A(17)='0' AND A( 6)='0' )then
          cVar2S19S123P064N004P007nsss(0) <='1';
          else
          cVar2S19S123P064N004P007nsss(0) <='0';
          end if;
        if(cVar1S20S123P017P036P065P019(0)='1' AND  E( 1)='1' AND D( 8)='0' )then
          cVar2S20S123P064P067nsss(0) <='1';
          else
          cVar2S20S123P064P067nsss(0) <='0';
          end if;
        if(cVar1S21S123P017P036P065P019(0)='1' AND  E( 1)='1' AND D( 8)='1' AND A(11)='0' )then
          cVar2S21S123P064P067P016nsss(0) <='1';
          else
          cVar2S21S123P064P067P016nsss(0) <='0';
          end if;
        if(cVar1S22S123P017P036P065P019(0)='1' AND  A(10)='0' AND D( 2)='0' AND D( 8)='1' )then
          cVar2S22S123P018P058P067nsss(0) <='1';
          else
          cVar2S22S123P018P058P067nsss(0) <='0';
          end if;
        if(cVar1S23S123P017P036P065P019(0)='1' AND  A(10)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar2S23S123P018P058P033nsss(0) <='1';
          else
          cVar2S23S123P018P058P033nsss(0) <='0';
          end if;
        if(cVar1S24S123P017P036P065P019(0)='1' AND  A(10)='1' AND D( 2)='1' AND A( 2)='0' )then
          cVar2S24S123P018P058P015nsss(0) <='1';
          else
          cVar2S24S123P018P058P015nsss(0) <='0';
          end if;
        if(cVar1S25S123P017P036P065P019(0)='1' AND  A(10)='1' AND D( 2)='0' AND A(13)='1' )then
          cVar2S25S123P018N058P012nsss(0) <='1';
          else
          cVar2S25S123P018N058P012nsss(0) <='0';
          end if;
        if(cVar1S26S123P017P036P065P063(0)='1' AND  A( 4)='1' AND E( 8)='1' )then
          cVar2S26S123P011P069nsss(0) <='1';
          else
          cVar2S26S123P011P069nsss(0) <='0';
          end if;
        if(cVar1S27S123P017P036P065P063(0)='1' AND  A( 4)='1' AND E( 8)='0' AND D( 0)='1' )then
          cVar2S27S123P011N069P066nsss(0) <='1';
          else
          cVar2S27S123P011N069P066nsss(0) <='0';
          end if;
        if(cVar1S28S123P017P036P065P063(0)='1' AND  A( 4)='0' AND E( 3)='1' )then
          cVar2S28S123N011P056nsss(0) <='1';
          else
          cVar2S28S123N011P056nsss(0) <='0';
          end if;
        if(cVar1S29S123P017P036P065P063(0)='1' AND  A( 4)='0' AND E( 3)='0' AND B( 5)='1' )then
          cVar2S29S123N011N056P027nsss(0) <='1';
          else
          cVar2S29S123N011N056P027nsss(0) <='0';
          end if;
        if(cVar1S30S123P017P036P065N063(0)='1' AND  D( 1)='0' AND A(10)='0' )then
          cVar2S30S123P062P018nsss(0) <='1';
          else
          cVar2S30S123P062P018nsss(0) <='0';
          end if;
        if(cVar1S31S123P017N036P060P069(0)='1' AND  A( 2)='0' AND B(10)='1' )then
          cVar2S31S123P015P034nsss(0) <='1';
          else
          cVar2S31S123P015P034nsss(0) <='0';
          end if;
        if(cVar1S32S123P017N036P060P069(0)='1' AND  A( 2)='0' AND B(10)='0' AND D( 0)='0' )then
          cVar2S32S123P015N034P066nsss(0) <='1';
          else
          cVar2S32S123P015N034P066nsss(0) <='0';
          end if;
        if(cVar1S33S123P017N036P060P069(0)='1' AND  A( 2)='1' AND A(12)='1' )then
          cVar2S33S123P015P014nsss(0) <='1';
          else
          cVar2S33S123P015P014nsss(0) <='0';
          end if;
        if(cVar1S34S123P017N036P060N069(0)='1' AND  A(19)='1' )then
          cVar2S34S123P000nsss(0) <='1';
          else
          cVar2S34S123P000nsss(0) <='0';
          end if;
        if(cVar1S35S123P017N036P060N069(0)='1' AND  A(19)='0' AND E(10)='0' )then
          cVar2S35S123N000P061nsss(0) <='1';
          else
          cVar2S35S123N000P061nsss(0) <='0';
          end if;
        if(cVar1S36S123P017N036P060N069(0)='1' AND  A(19)='0' AND E(10)='1' AND A( 4)='1' )then
          cVar2S36S123N000P061P011nsss(0) <='1';
          else
          cVar2S36S123N000P061P011nsss(0) <='0';
          end if;
        if(cVar1S37S123P017N036N060P037(0)='1' AND  A(14)='1' AND B(13)='1' )then
          cVar2S37S123P010P028nsss(0) <='1';
          else
          cVar2S37S123P010P028nsss(0) <='0';
          end if;
        if(cVar1S38S123P017N036N060P037(0)='1' AND  A(14)='1' AND B(13)='0' AND D(11)='0' )then
          cVar2S38S123P010N028P055nsss(0) <='1';
          else
          cVar2S38S123P010N028P055nsss(0) <='0';
          end if;
        if(cVar1S39S123P017N036N060P037(0)='1' AND  A(14)='0' AND D( 6)='0' AND A(11)='0' )then
          cVar2S39S123N010P042P016nsss(0) <='1';
          else
          cVar2S39S123N010P042P016nsss(0) <='0';
          end if;
        if(cVar1S40S123P017N036N060P037(0)='1' AND  A(14)='0' AND D( 6)='1' AND A( 0)='0' )then
          cVar2S40S123N010P042P019nsss(0) <='1';
          else
          cVar2S40S123N010P042P019nsss(0) <='0';
          end if;
        if(cVar1S41S123P017N036N060N037(0)='1' AND  A(12)='1' AND B(10)='1' AND B( 1)='0' )then
          cVar2S41S123P014P034P035nsss(0) <='1';
          else
          cVar2S41S123P014P034P035nsss(0) <='0';
          end if;
        if(cVar1S42S123P017N036N060N037(0)='1' AND  A(12)='1' AND B(10)='0' AND B( 6)='1' )then
          cVar2S42S123P014N034P025nsss(0) <='1';
          else
          cVar2S42S123P014N034P025nsss(0) <='0';
          end if;
        if(cVar1S43S123P017N036N060N037(0)='1' AND  A(12)='0' AND B(13)='1' )then
          cVar2S43S123N014P028nsss(0) <='1';
          else
          cVar2S43S123N014P028nsss(0) <='0';
          end if;
        if(cVar1S0S124P036P065P032P019(0)='1' AND  E( 7)='0' AND A(13)='0' AND B( 7)='0' )then
          cVar2S0S124P040P012P023nsss(0) <='1';
          else
          cVar2S0S124P040P012P023nsss(0) <='0';
          end if;
        if(cVar1S1S124P036P065P032P019(0)='1' AND  E( 7)='0' AND A(13)='1' AND E(11)='1' )then
          cVar2S1S124P040P012P057nsss(0) <='1';
          else
          cVar2S1S124P040P012P057nsss(0) <='0';
          end if;
        if(cVar1S2S124P036P065P032P019(0)='1' AND  E( 7)='1' AND A( 1)='1' )then
          cVar2S2S124P040P017nsss(0) <='1';
          else
          cVar2S2S124P040P017nsss(0) <='0';
          end if;
        if(cVar1S3S124P036P065P032P019(0)='1' AND  D( 6)='1' AND E( 8)='1' AND A(11)='0' )then
          cVar2S3S124P042P069P016nsss(0) <='1';
          else
          cVar2S3S124P042P069P016nsss(0) <='0';
          end if;
        if(cVar1S4S124P036P065P032P019(0)='1' AND  D( 6)='0' AND B( 7)='0' )then
          cVar2S4S124N042P023nsss(0) <='1';
          else
          cVar2S4S124N042P023nsss(0) <='0';
          end if;
        if(cVar1S5S124P036P065P032P055(0)='1' AND  A( 8)='0' AND D( 0)='1' AND A( 2)='1' )then
          cVar2S5S124P003P066P015nsss(0) <='1';
          else
          cVar2S5S124P003P066P015nsss(0) <='0';
          end if;
        if(cVar1S6S124P036P065P032P055(0)='1' AND  A( 8)='0' AND D( 0)='0' AND A( 0)='1' )then
          cVar2S6S124P003N066P019nsss(0) <='1';
          else
          cVar2S6S124P003N066P019nsss(0) <='0';
          end if;
        if(cVar1S7S124P036P065P024P063(0)='1' AND  A( 1)='1' AND B( 0)='0' )then
          cVar2S7S124P017P037nsss(0) <='1';
          else
          cVar2S7S124P017P037nsss(0) <='0';
          end if;
        if(cVar1S8S124P036P065P024P063(0)='1' AND  A( 1)='1' AND B( 0)='1' AND B(10)='1' )then
          cVar2S8S124P017P037P034nsss(0) <='1';
          else
          cVar2S8S124P017P037P034nsss(0) <='0';
          end if;
        if(cVar1S9S124P036P065P024P063(0)='1' AND  A( 1)='0' AND B( 2)='1' AND E( 2)='0' )then
          cVar2S9S124N017P033P060nsss(0) <='1';
          else
          cVar2S9S124N017P033P060nsss(0) <='0';
          end if;
        if(cVar1S10S124P036P065P024P063(0)='1' AND  A( 1)='0' AND B( 2)='0' AND E( 2)='1' )then
          cVar2S10S124N017N033P060nsss(0) <='1';
          else
          cVar2S10S124N017N033P060nsss(0) <='0';
          end if;
        if(cVar1S11S124P036P065P024N063(0)='1' AND  A( 2)='1' AND A( 0)='1' )then
          cVar2S11S124P015P019nsss(0) <='1';
          else
          cVar2S11S124P015P019nsss(0) <='0';
          end if;
        if(cVar1S12S124P036P065P024N063(0)='1' AND  A( 2)='0' AND A(10)='0' AND E( 0)='0' )then
          cVar2S12S124N015P018P068nsss(0) <='1';
          else
          cVar2S12S124N015P018P068nsss(0) <='0';
          end if;
        if(cVar1S13S124P036P065P024N063(0)='1' AND  A( 2)='0' AND A(10)='1' AND A(12)='1' )then
          cVar2S13S124N015P018P014nsss(0) <='1';
          else
          cVar2S13S124N015P018P014nsss(0) <='0';
          end if;
        if(cVar1S14S124P036P065P024P034(0)='1' AND  D( 8)='0' AND A( 1)='1' )then
          cVar2S14S124P067P017nsss(0) <='1';
          else
          cVar2S14S124P067P017nsss(0) <='0';
          end if;
        if(cVar1S16S124N036P017P034N043(0)='1' AND  A( 5)='1' AND D( 2)='1' )then
          cVar2S16S124P009P058nsss(0) <='1';
          else
          cVar2S16S124P009P058nsss(0) <='0';
          end if;
        if(cVar1S17S124N036P017P034N043(0)='1' AND  A( 5)='1' AND D( 2)='0' AND D( 0)='1' )then
          cVar2S17S124P009N058P066nsss(0) <='1';
          else
          cVar2S17S124P009N058P066nsss(0) <='0';
          end if;
        if(cVar1S18S124N036P017P034N043(0)='1' AND  A( 5)='0' AND B(17)='1' AND A(10)='1' )then
          cVar2S18S124N009P020P018nsss(0) <='1';
          else
          cVar2S18S124N009P020P018nsss(0) <='0';
          end if;
        if(cVar1S19S124N036P017P034N043(0)='1' AND  A( 5)='0' AND B(17)='0' AND B( 4)='0' )then
          cVar2S19S124N009N020P029nsss(0) <='1';
          else
          cVar2S19S124N009N020P029nsss(0) <='0';
          end if;
        if(cVar1S20S124N036P017N034P002(0)='1' AND  A(14)='1' AND D(15)='0' )then
          cVar2S20S124P010P039nsss(0) <='1';
          else
          cVar2S20S124P010P039nsss(0) <='0';
          end if;
        if(cVar1S21S124N036P017N034P002(0)='1' AND  A(14)='0' AND D( 5)='1' AND D( 2)='0' )then
          cVar2S21S124N010P046P058nsss(0) <='1';
          else
          cVar2S21S124N010P046P058nsss(0) <='0';
          end if;
        if(cVar1S22S124N036P017N034P002(0)='1' AND  E( 7)='1' )then
          cVar2S22S124P040nsss(0) <='1';
          else
          cVar2S22S124P040nsss(0) <='0';
          end if;
        if(cVar1S23S124N036P017N034P002(0)='1' AND  E( 7)='0' AND B( 0)='1' AND A(11)='1' )then
          cVar2S23S124N040P037P016nsss(0) <='1';
          else
          cVar2S23S124N040P037P016nsss(0) <='0';
          end if;
        if(cVar1S24S124N036N017P032P031(0)='1' AND  E( 4)='0' AND A( 7)='0' AND E(15)='0' )then
          cVar2S24S124P052P005P041nsss(0) <='1';
          else
          cVar2S24S124P052P005P041nsss(0) <='0';
          end if;
        if(cVar1S25S124N036N017P032P031(0)='1' AND  E( 4)='1' AND D(10)='0' AND A(12)='1' )then
          cVar2S25S124P052P059P014nsss(0) <='1';
          else
          cVar2S25S124P052P059P014nsss(0) <='0';
          end if;
        if(cVar1S26S124N036N017P032P031(0)='1' AND  A(13)='0' AND A(12)='0' )then
          cVar2S26S124P012P014nsss(0) <='1';
          else
          cVar2S26S124P012P014nsss(0) <='0';
          end if;
        if(cVar1S27S124N036N017P032P031(0)='1' AND  A(13)='0' AND A(12)='1' AND D( 3)='1' )then
          cVar2S27S124P012P014P054nsss(0) <='1';
          else
          cVar2S27S124P012P014P054nsss(0) <='0';
          end if;
        if(cVar1S28S124N036N017N032P046(0)='1' AND  E( 7)='0' AND B( 6)='1' )then
          cVar2S28S124P040P025nsss(0) <='1';
          else
          cVar2S28S124P040P025nsss(0) <='0';
          end if;
        if(cVar1S29S124N036N017N032P046(0)='1' AND  E( 7)='0' AND B( 6)='0' AND A(15)='1' )then
          cVar2S29S124P040N025P008nsss(0) <='1';
          else
          cVar2S29S124P040N025P008nsss(0) <='0';
          end if;
        if(cVar1S30S124N036N017N032N046(0)='1' AND  B( 6)='0' AND B( 7)='1' AND B(10)='0' )then
          cVar2S30S124P025P023P034nsss(0) <='1';
          else
          cVar2S30S124P025P023P034nsss(0) <='0';
          end if;
        if(cVar1S31S124N036N017N032N046(0)='1' AND  B( 6)='1' AND D(13)='1' AND A( 6)='1' )then
          cVar2S31S124P025P047P007nsss(0) <='1';
          else
          cVar2S31S124P025P047P007nsss(0) <='0';
          end if;
        if(cVar1S0S125P032P064P050P022(0)='1' AND  D( 8)='0' AND E( 8)='1' AND E( 0)='0' )then
          cVar2S0S125P067P069P068nsss(0) <='1';
          else
          cVar2S0S125P067P069P068nsss(0) <='0';
          end if;
        if(cVar1S1S125P032P064P050P022(0)='1' AND  D( 8)='0' AND E( 8)='0' )then
          cVar2S1S125P067N069psss(0) <='1';
          else
          cVar2S1S125P067N069psss(0) <='0';
          end if;
        if(cVar1S2S125P032P064P050P022(0)='1' AND  D( 8)='1' AND B( 0)='0' )then
          cVar2S2S125P067P037nsss(0) <='1';
          else
          cVar2S2S125P067P037nsss(0) <='0';
          end if;
        if(cVar1S3S125P032P064P050P022(0)='1' AND  B( 9)='0' AND A(12)='1' )then
          cVar2S3S125P036P014nsss(0) <='1';
          else
          cVar2S3S125P036P014nsss(0) <='0';
          end if;
        if(cVar1S4S125P032P064P050P022(0)='1' AND  B( 9)='0' AND A(12)='0' AND A(10)='1' )then
          cVar2S4S125P036N014P018nsss(0) <='1';
          else
          cVar2S4S125P036N014P018nsss(0) <='0';
          end if;
        if(cVar1S5S125P032P064P050P027(0)='1' AND  D( 9)='0' )then
          cVar2S5S125P063nsss(0) <='1';
          else
          cVar2S5S125P063nsss(0) <='0';
          end if;
        if(cVar1S6S125P032P064P050N027(0)='1' AND  B( 1)='1' AND B( 0)='1' )then
          cVar2S6S125P035P037nsss(0) <='1';
          else
          cVar2S6S125P035P037nsss(0) <='0';
          end if;
        if(cVar1S7S125P032P064P050N027(0)='1' AND  B( 1)='1' AND B( 0)='0' AND E( 4)='1' )then
          cVar2S7S125P035N037P052nsss(0) <='1';
          else
          cVar2S7S125P035N037P052nsss(0) <='0';
          end if;
        if(cVar1S8S125P032P064P050N027(0)='1' AND  B( 1)='0' AND E( 8)='1' )then
          cVar2S8S125N035P069nsss(0) <='1';
          else
          cVar2S8S125N035P069nsss(0) <='0';
          end if;
        if(cVar1S9S125P032N064P037P068(0)='1' AND  E( 4)='0' AND A( 3)='1' AND B(13)='0' )then
          cVar2S9S125P052P013P028nsss(0) <='1';
          else
          cVar2S9S125P052P013P028nsss(0) <='0';
          end if;
        if(cVar1S10S125P032N064P037P068(0)='1' AND  E( 4)='0' AND A( 3)='0' )then
          cVar2S10S125P052N013psss(0) <='1';
          else
          cVar2S10S125P052N013psss(0) <='0';
          end if;
        if(cVar1S11S125P032N064P037P068(0)='1' AND  E( 4)='1' AND D( 4)='1' AND A(12)='0' )then
          cVar2S11S125P052P050P014nsss(0) <='1';
          else
          cVar2S11S125P052P050P014nsss(0) <='0';
          end if;
        if(cVar1S12S125P032N064P037N068(0)='1' AND  B(12)='1' AND B( 3)='0' AND A(13)='1' )then
          cVar2S12S125P030P031P012nsss(0) <='1';
          else
          cVar2S12S125P030P031P012nsss(0) <='0';
          end if;
        if(cVar1S13S125P032N064P037N068(0)='1' AND  B(12)='0' AND A(17)='1' )then
          cVar2S13S125N030P004nsss(0) <='1';
          else
          cVar2S13S125N030P004nsss(0) <='0';
          end if;
        if(cVar1S14S125P032N064P037N068(0)='1' AND  B(12)='0' AND A(17)='0' AND B( 2)='1' )then
          cVar2S14S125N030N004P033nsss(0) <='1';
          else
          cVar2S14S125N030N004P033nsss(0) <='0';
          end if;
        if(cVar1S15S125P032N064P037P056(0)='1' AND  D( 8)='1' AND D( 0)='0' )then
          cVar2S15S125P067P066nsss(0) <='1';
          else
          cVar2S15S125P067P066nsss(0) <='0';
          end if;
        if(cVar1S16S125P032N064P037P056(0)='1' AND  D( 8)='1' AND D( 0)='1' AND A(11)='0' )then
          cVar2S16S125P067P066P016nsss(0) <='1';
          else
          cVar2S16S125P067P066P016nsss(0) <='0';
          end if;
        if(cVar1S17S125P032N064P037P056(0)='1' AND  D( 8)='0' AND E( 9)='1' AND A(11)='0' )then
          cVar2S17S125N067P065P016nsss(0) <='1';
          else
          cVar2S17S125N067P065P016nsss(0) <='0';
          end if;
        if(cVar1S18S125P032N064P037P056(0)='1' AND  D( 8)='0' AND E( 9)='0' AND B( 3)='1' )then
          cVar2S18S125N067N065P031nsss(0) <='1';
          else
          cVar2S18S125N067N065P031nsss(0) <='0';
          end if;
        if(cVar1S19S125P032N064P037N056(0)='1' AND  A(11)='1' AND B(15)='0' AND E( 0)='1' )then
          cVar2S19S125P016P024P068nsss(0) <='1';
          else
          cVar2S19S125P016P024P068nsss(0) <='0';
          end if;
        if(cVar1S20S125P032N064P037N056(0)='1' AND  A(11)='1' AND B(15)='1' AND E( 0)='0' )then
          cVar2S20S125P016P024P068nsss(0) <='1';
          else
          cVar2S20S125P016P024P068nsss(0) <='0';
          end if;
        if(cVar1S21S125P032N064P037N056(0)='1' AND  A(11)='0' AND A( 6)='0' AND B( 2)='1' )then
          cVar2S21S125N016P007P033nsss(0) <='1';
          else
          cVar2S21S125N016P007P033nsss(0) <='0';
          end if;
        if(cVar1S22S125P032P037P063P016(0)='1' AND  A( 0)='1' )then
          cVar2S22S125P019nsss(0) <='1';
          else
          cVar2S22S125P019nsss(0) <='0';
          end if;
        if(cVar1S23S125P032P037P063P016(0)='1' AND  A( 0)='0' AND A(12)='1' )then
          cVar2S23S125N019P014nsss(0) <='1';
          else
          cVar2S23S125N019P014nsss(0) <='0';
          end if;
        if(cVar1S24S125P032P037P063P016(0)='1' AND  A(12)='0' )then
          cVar2S24S125P014nsss(0) <='1';
          else
          cVar2S24S125P014nsss(0) <='0';
          end if;
        if(cVar1S25S125P032P037N063P012(0)='1' AND  A( 4)='0' AND A( 5)='0' AND B(12)='0' )then
          cVar2S25S125P011P009P030nsss(0) <='1';
          else
          cVar2S25S125P011P009P030nsss(0) <='0';
          end if;
        if(cVar1S26S125P032P037N063P012(0)='1' AND  A( 4)='1' AND A( 0)='1' )then
          cVar2S26S125P011P019nsss(0) <='1';
          else
          cVar2S26S125P011P019nsss(0) <='0';
          end if;
        if(cVar1S27S125P032P037N063N012(0)='1' AND  E( 3)='0' AND A( 2)='1' )then
          cVar2S27S125P056P015nsss(0) <='1';
          else
          cVar2S27S125P056P015nsss(0) <='0';
          end if;
        if(cVar1S28S125P032P037N063N012(0)='1' AND  E( 3)='1' AND A(12)='1' )then
          cVar2S28S125P056P014nsss(0) <='1';
          else
          cVar2S28S125P056P014nsss(0) <='0';
          end if;
        if(cVar1S29S125P032N037P031P068(0)='1' AND  A( 1)='1' AND D(10)='1' )then
          cVar2S29S125P017P059nsss(0) <='1';
          else
          cVar2S29S125P017P059nsss(0) <='0';
          end if;
        if(cVar1S30S125P032N037P031P068(0)='1' AND  A( 1)='1' AND D(10)='0' AND A(10)='0' )then
          cVar2S30S125P017N059P018nsss(0) <='1';
          else
          cVar2S30S125P017N059P018nsss(0) <='0';
          end if;
        if(cVar1S31S125P032N037P031P068(0)='1' AND  A( 1)='0' AND A( 8)='0' AND D( 9)='1' )then
          cVar2S31S125N017P003P063nsss(0) <='1';
          else
          cVar2S31S125N017P003P063nsss(0) <='0';
          end if;
        if(cVar1S32S125P032N037P031N068(0)='1' AND  A(15)='1' AND B( 2)='1' AND A(12)='1' )then
          cVar2S32S125P008P033P014nsss(0) <='1';
          else
          cVar2S32S125P008P033P014nsss(0) <='0';
          end if;
        if(cVar1S33S125P032N037P031N068(0)='1' AND  A(15)='1' AND B( 2)='0' AND A( 4)='1' )then
          cVar2S33S125P008N033P011nsss(0) <='1';
          else
          cVar2S33S125P008N033P011nsss(0) <='0';
          end if;
        if(cVar1S34S125P032N037P031P012(0)='1' AND  D( 3)='1' AND A( 3)='0' )then
          cVar2S34S125P054P013nsss(0) <='1';
          else
          cVar2S34S125P054P013nsss(0) <='0';
          end if;
        if(cVar1S35S125P032N037P031P012(0)='1' AND  D( 3)='0' AND E(11)='1' )then
          cVar2S35S125N054P057nsss(0) <='1';
          else
          cVar2S35S125N054P057nsss(0) <='0';
          end if;
        if(cVar1S36S125P032N037P031P012(0)='1' AND  E( 3)='1' AND A( 2)='0' )then
          cVar2S36S125P056P015nsss(0) <='1';
          else
          cVar2S36S125P056P015nsss(0) <='0';
          end if;
        if(cVar1S1S126P069P018P026N064(0)='1' AND  A( 0)='1' )then
          cVar2S1S126P019nsss(0) <='1';
          else
          cVar2S1S126P019nsss(0) <='0';
          end if;
        if(cVar1S2S126P069P018P026N064(0)='1' AND  A( 0)='0' AND A(13)='0' AND A( 1)='1' )then
          cVar2S2S126N019P012P017nsss(0) <='1';
          else
          cVar2S2S126N019P012P017nsss(0) <='0';
          end if;
        if(cVar1S3S126P069P018N026P031(0)='1' AND  A(15)='0' )then
          cVar2S3S126P008nsss(0) <='1';
          else
          cVar2S3S126P008nsss(0) <='0';
          end if;
        if(cVar1S4S126P069P018N026N031(0)='1' AND  D( 8)='0' AND E( 1)='1' )then
          cVar2S4S126P067P064nsss(0) <='1';
          else
          cVar2S4S126P067P064nsss(0) <='0';
          end if;
        if(cVar1S5S126P069P018N026N031(0)='1' AND  D( 8)='0' AND E( 1)='0' AND E( 2)='1' )then
          cVar2S5S126P067N064P060nsss(0) <='1';
          else
          cVar2S5S126P067N064P060nsss(0) <='0';
          end if;
        if(cVar1S6S126P069P018N026N031(0)='1' AND  D( 8)='1' AND E(14)='1' )then
          cVar2S6S126P067P045nsss(0) <='1';
          else
          cVar2S6S126P067P045nsss(0) <='0';
          end if;
        if(cVar1S7S126P069P018N026N031(0)='1' AND  D( 8)='1' AND E(14)='0' AND A(12)='0' )then
          cVar2S7S126P067N045P014nsss(0) <='1';
          else
          cVar2S7S126P067N045P014nsss(0) <='0';
          end if;
        if(cVar1S8S126P069P018P068P067(0)='1' AND  D( 1)='0' AND A( 0)='0' )then
          cVar2S8S126P062P019nsss(0) <='1';
          else
          cVar2S8S126P062P019nsss(0) <='0';
          end if;
        if(cVar1S9S126P069P018P068P067(0)='1' AND  D( 1)='0' AND A( 0)='1' AND A( 1)='0' )then
          cVar2S9S126P062P019P017nsss(0) <='1';
          else
          cVar2S9S126P062P019P017nsss(0) <='0';
          end if;
        if(cVar1S10S126P069P018P068P067(0)='1' AND  D( 1)='1' AND D( 9)='0' AND A(12)='1' )then
          cVar2S10S126P062P063P014nsss(0) <='1';
          else
          cVar2S10S126P062P063P014nsss(0) <='0';
          end if;
        if(cVar1S11S126P069P018P068N067(0)='1' AND  E( 1)='1' AND D( 9)='1' )then
          cVar2S11S126P064P063nsss(0) <='1';
          else
          cVar2S11S126P064P063nsss(0) <='0';
          end if;
        if(cVar1S12S126P069P018P068N067(0)='1' AND  E( 1)='0' AND A( 0)='0' AND A( 3)='1' )then
          cVar2S12S126N064P019P013nsss(0) <='1';
          else
          cVar2S12S126N064P019P013nsss(0) <='0';
          end if;
        if(cVar1S14S126P069P018P068N040(0)='1' AND  D( 9)='1' AND A( 0)='1' )then
          cVar2S14S126P063P019nsss(0) <='1';
          else
          cVar2S14S126P063P019nsss(0) <='0';
          end if;
        if(cVar1S15S126P069P018P068N040(0)='1' AND  D( 9)='1' AND A( 0)='0' AND E( 9)='1' )then
          cVar2S15S126P063N019P065nsss(0) <='1';
          else
          cVar2S15S126P063N019P065nsss(0) <='0';
          end if;
        if(cVar1S16S126P069P018P068N040(0)='1' AND  D( 9)='0' AND B( 2)='0' AND A(13)='1' )then
          cVar2S16S126N063P033P012nsss(0) <='1';
          else
          cVar2S16S126N063P033P012nsss(0) <='0';
          end if;
        if(cVar1S17S126N069P018P049P032(0)='1' AND  A(12)='0' AND A( 2)='0' )then
          cVar2S17S126P014P015nsss(0) <='1';
          else
          cVar2S17S126P014P015nsss(0) <='0';
          end if;
        if(cVar1S18S126N069P018P049P032(0)='1' AND  A(12)='0' AND A( 2)='1' AND A(13)='1' )then
          cVar2S18S126P014P015P012nsss(0) <='1';
          else
          cVar2S18S126P014P015P012nsss(0) <='0';
          end if;
        if(cVar1S19S126N069P018P049P032(0)='1' AND  A(12)='1' AND A( 3)='0' AND D(13)='0' )then
          cVar2S19S126P014P013P047nsss(0) <='1';
          else
          cVar2S19S126P014P013P047nsss(0) <='0';
          end if;
        if(cVar1S20S126N069P018N049P032(0)='1' AND  E(14)='0' AND A(18)='0' )then
          cVar2S20S126P045P002nsss(0) <='1';
          else
          cVar2S20S126P045P002nsss(0) <='0';
          end if;
        if(cVar1S21S126N069P018N049N032(0)='1' AND  D(14)='1' AND B(16)='1' )then
          cVar2S21S126P043P022nsss(0) <='1';
          else
          cVar2S21S126P043P022nsss(0) <='0';
          end if;
        if(cVar1S22S126N069P018N049N032(0)='1' AND  D(14)='1' AND B(16)='0' AND B( 7)='1' )then
          cVar2S22S126P043N022P023nsss(0) <='1';
          else
          cVar2S22S126P043N022P023nsss(0) <='0';
          end if;
        if(cVar1S23S126N069P018N049N032(0)='1' AND  D(14)='0' AND B(16)='0' AND B( 3)='1' )then
          cVar2S23S126N043P022P031nsss(0) <='1';
          else
          cVar2S23S126N043P022P031nsss(0) <='0';
          end if;
        if(cVar1S24S126N069N018P066P064(0)='1' AND  E( 0)='0' AND E( 9)='1' AND E( 2)='0' )then
          cVar2S24S126P068P065P060nsss(0) <='1';
          else
          cVar2S24S126P068P065P060nsss(0) <='0';
          end if;
        if(cVar1S25S126N069N018P066P064(0)='1' AND  E( 0)='1' AND D( 2)='1' AND D( 1)='0' )then
          cVar2S25S126P068P058P062nsss(0) <='1';
          else
          cVar2S25S126P068P058P062nsss(0) <='0';
          end if;
        if(cVar1S26S126N069N018P066P064(0)='1' AND  E( 0)='1' AND D( 2)='0' AND B(11)='1' )then
          cVar2S26S126P068N058P032nsss(0) <='1';
          else
          cVar2S26S126P068N058P032nsss(0) <='0';
          end if;
        if(cVar1S27S126N069N018P066P064(0)='1' AND  D( 1)='1' AND E( 0)='1' AND A(11)='1' )then
          cVar2S27S126P062P068P016nsss(0) <='1';
          else
          cVar2S27S126P062P068P016nsss(0) <='0';
          end if;
        if(cVar1S28S126N069N018P066P064(0)='1' AND  D( 1)='1' AND E( 0)='0' AND E( 9)='0' )then
          cVar2S28S126P062N068P065nsss(0) <='1';
          else
          cVar2S28S126P062N068P065nsss(0) <='0';
          end if;
        if(cVar1S29S126N069N018P066P064(0)='1' AND  D( 1)='0' AND A( 2)='1' AND A(11)='0' )then
          cVar2S29S126N062P015P016nsss(0) <='1';
          else
          cVar2S29S126N062P015P016nsss(0) <='0';
          end if;
        if(cVar1S30S126N069N018P066P064(0)='1' AND  D( 1)='0' AND A( 2)='0' AND A(16)='1' )then
          cVar2S30S126N062N015P006nsss(0) <='1';
          else
          cVar2S30S126N062N015P006nsss(0) <='0';
          end if;
        if(cVar1S31S126N069N018P066P006(0)='1' AND  D(13)='0' AND A( 6)='1' AND E(12)='1' )then
          cVar2S31S126P047P007P053nsss(0) <='1';
          else
          cVar2S31S126P047P007P053nsss(0) <='0';
          end if;
        if(cVar1S32S126N069N018P066P006(0)='1' AND  D(13)='1' AND A( 0)='1' AND B(15)='1' )then
          cVar2S32S126P047P019P024nsss(0) <='1';
          else
          cVar2S32S126P047P019P024nsss(0) <='0';
          end if;
        if(cVar1S33S126N069N018P066P006(0)='1' AND  B(15)='1' AND A( 0)='0' )then
          cVar2S33S126P024P019nsss(0) <='1';
          else
          cVar2S33S126P024P019nsss(0) <='0';
          end if;
        if(cVar1S34S126N069N018P066P006(0)='1' AND  B(15)='1' AND A( 0)='1' AND E(13)='0' )then
          cVar2S34S126P024P019P049nsss(0) <='1';
          else
          cVar2S34S126P024P019P049nsss(0) <='0';
          end if;
        if(cVar1S35S126N069N018P066P006(0)='1' AND  B(15)='0' AND B( 1)='1' AND A( 2)='1' )then
          cVar2S35S126N024P035P015nsss(0) <='1';
          else
          cVar2S35S126N024P035P015nsss(0) <='0';
          end if;
        if(cVar1S36S126N069N018P066P006(0)='1' AND  B(15)='0' AND B( 1)='0' AND E( 5)='1' )then
          cVar2S36S126N024N035P048nsss(0) <='1';
          else
          cVar2S36S126N024N035P048nsss(0) <='0';
          end if;
        if(cVar1S0S127P064P069P034P016(0)='1' AND  A(19)='0' )then
          cVar2S0S127P000nsss(0) <='1';
          else
          cVar2S0S127P000nsss(0) <='0';
          end if;
        if(cVar1S1S127P064P069P034P016(0)='1' AND  A(19)='1' AND E( 6)='0' AND E( 4)='1' )then
          cVar2S1S127P000P044P052nsss(0) <='1';
          else
          cVar2S1S127P000P044P052nsss(0) <='0';
          end if;
        if(cVar1S2S127P064P069P034P016(0)='1' AND  D( 8)='0' AND B( 6)='0' )then
          cVar2S2S127P067P025nsss(0) <='1';
          else
          cVar2S2S127P067P025nsss(0) <='0';
          end if;
        if(cVar1S3S127P064P069P034P016(0)='1' AND  D( 8)='0' AND B( 6)='1' AND A(14)='1' )then
          cVar2S3S127P067P025P010nsss(0) <='1';
          else
          cVar2S3S127P067P025P010nsss(0) <='0';
          end if;
        if(cVar1S4S127P064P069P034P016(0)='1' AND  D( 8)='1' AND D( 0)='1' AND A( 0)='1' )then
          cVar2S4S127P067P066P019nsss(0) <='1';
          else
          cVar2S4S127P067P066P019nsss(0) <='0';
          end if;
        if(cVar1S5S127P064P069P034P016(0)='1' AND  D( 8)='1' AND D( 0)='0' AND B(14)='1' )then
          cVar2S5S127P067N066P026nsss(0) <='1';
          else
          cVar2S5S127P067N066P026nsss(0) <='0';
          end if;
        if(cVar1S6S127P064P069P034P008(0)='1' AND  B( 9)='0' AND D(12)='1' AND B(13)='1' )then
          cVar2S6S127P036P051P028nsss(0) <='1';
          else
          cVar2S6S127P036P051P028nsss(0) <='0';
          end if;
        if(cVar1S7S127P064P069P034P008(0)='1' AND  B( 9)='0' AND D(12)='0' AND A(14)='0' )then
          cVar2S7S127P036N051P010nsss(0) <='1';
          else
          cVar2S7S127P036N051P010nsss(0) <='0';
          end if;
        if(cVar1S8S127P064P069P034P008(0)='1' AND  B( 9)='1' AND B(12)='0' AND A(12)='0' )then
          cVar2S8S127P036P030P014nsss(0) <='1';
          else
          cVar2S8S127P036P030P014nsss(0) <='0';
          end if;
        if(cVar1S9S127P064P069P034P008(0)='1' AND  B(14)='1' )then
          cVar2S9S127P026nsss(0) <='1';
          else
          cVar2S9S127P026nsss(0) <='0';
          end if;
        if(cVar1S10S127P064P069P034P008(0)='1' AND  B(14)='0' AND D( 8)='0' AND D( 0)='1' )then
          cVar2S10S127N026P067P066nsss(0) <='1';
          else
          cVar2S10S127N026P067P066nsss(0) <='0';
          end if;
        if(cVar1S11S127P064P069P037P016(0)='1' AND  A( 6)='0' AND A(19)='1' AND E( 0)='1' )then
          cVar2S11S127P007P000P068nsss(0) <='1';
          else
          cVar2S11S127P007P000P068nsss(0) <='0';
          end if;
        if(cVar1S12S127P064P069P037P016(0)='1' AND  A( 6)='0' AND A(19)='0' )then
          cVar2S12S127P007N000psss(0) <='1';
          else
          cVar2S12S127P007N000psss(0) <='0';
          end if;
        if(cVar1S13S127P064P069P037P016(0)='1' AND  A( 6)='1' AND A( 4)='1' )then
          cVar2S13S127P007P011nsss(0) <='1';
          else
          cVar2S13S127P007P011nsss(0) <='0';
          end if;
        if(cVar1S14S127P064P069P037P016(0)='1' AND  A( 7)='0' AND D(12)='1' )then
          cVar2S14S127P005P051nsss(0) <='1';
          else
          cVar2S14S127P005P051nsss(0) <='0';
          end if;
        if(cVar1S15S127P064P069N037P016(0)='1' AND  A(15)='1' AND E( 2)='1' )then
          cVar2S15S127P008P060nsss(0) <='1';
          else
          cVar2S15S127P008P060nsss(0) <='0';
          end if;
        if(cVar1S16S127P064P069N037P016(0)='1' AND  A(15)='1' AND E( 2)='0' AND A(12)='0' )then
          cVar2S16S127P008N060P014nsss(0) <='1';
          else
          cVar2S16S127P008N060P014nsss(0) <='0';
          end if;
        if(cVar1S17S127P064P069N037P016(0)='1' AND  A(15)='0' AND E( 4)='1' )then
          cVar2S17S127N008P052nsss(0) <='1';
          else
          cVar2S17S127N008P052nsss(0) <='0';
          end if;
        if(cVar1S18S127P064P069N037P016(0)='1' AND  A(15)='0' AND E( 4)='0' AND A(14)='0' )then
          cVar2S18S127N008N052P010nsss(0) <='1';
          else
          cVar2S18S127N008N052P010nsss(0) <='0';
          end if;
        if(cVar1S19S127P064P069N037N016(0)='1' AND  E(12)='0' AND A( 1)='1' AND D( 0)='1' )then
          cVar2S19S127P053P017P066nsss(0) <='1';
          else
          cVar2S19S127P053P017P066nsss(0) <='0';
          end if;
        if(cVar1S20S127P064P069N037N016(0)='1' AND  E(12)='0' AND A( 1)='0' AND A( 6)='1' )then
          cVar2S20S127P053N017P007nsss(0) <='1';
          else
          cVar2S20S127P053N017P007nsss(0) <='0';
          end if;
        if(cVar1S21S127P064P069N037N016(0)='1' AND  E(12)='1' AND A(14)='1' )then
          cVar2S21S127P053P010nsss(0) <='1';
          else
          cVar2S21S127P053P010nsss(0) <='0';
          end if;
        if(cVar1S22S127P064P018P054P035(0)='1' AND  A( 2)='0' AND A( 3)='0' )then
          cVar2S22S127P015P013nsss(0) <='1';
          else
          cVar2S22S127P015P013nsss(0) <='0';
          end if;
        if(cVar1S23S127P064P018P054P035(0)='1' AND  A( 2)='1' AND D( 9)='1' AND A( 4)='0' )then
          cVar2S23S127P015P063P011nsss(0) <='1';
          else
          cVar2S23S127P015P063P011nsss(0) <='0';
          end if;
        if(cVar1S24S127P064P018P054P035(0)='1' AND  A( 2)='1' AND D( 9)='0' AND A( 3)='1' )then
          cVar2S24S127P015N063P013nsss(0) <='1';
          else
          cVar2S24S127P015N063P013nsss(0) <='0';
          end if;
        if(cVar1S25S127P064P018P054P035(0)='1' AND  D( 9)='0' AND D( 8)='0' AND B(10)='0' )then
          cVar2S25S127P063P067P034nsss(0) <='1';
          else
          cVar2S25S127P063P067P034nsss(0) <='0';
          end if;
        if(cVar1S26S127P064P018P054P035(0)='1' AND  D( 9)='0' AND D( 8)='1' AND A( 1)='0' )then
          cVar2S26S127P063P067P017nsss(0) <='1';
          else
          cVar2S26S127P063P067P017nsss(0) <='0';
          end if;
        if(cVar1S27S127P064P018P054P035(0)='1' AND  D( 9)='1' AND A( 0)='1' AND A( 1)='1' )then
          cVar2S27S127P063P019P017nsss(0) <='1';
          else
          cVar2S27S127P063P019P017nsss(0) <='0';
          end if;
        if(cVar1S28S127P064P018P054P035(0)='1' AND  D( 9)='1' AND A( 0)='0' AND A( 1)='0' )then
          cVar2S28S127P063N019P017nsss(0) <='1';
          else
          cVar2S28S127P063N019P017nsss(0) <='0';
          end if;
        if(cVar1S30S127P064P018P054N065(0)='1' AND  E( 4)='1' )then
          cVar2S30S127P052nsss(0) <='1';
          else
          cVar2S30S127P052nsss(0) <='0';
          end if;
        if(cVar1S31S127P064P018P054N065(0)='1' AND  E( 4)='0' AND A( 0)='1' AND A(11)='1' )then
          cVar2S31S127N052P019P016nsss(0) <='1';
          else
          cVar2S31S127N052P019P016nsss(0) <='0';
          end if;
        if(cVar1S32S127P064N018P050P048(0)='1' AND  A( 8)='1' AND A( 2)='1' AND B( 0)='0' )then
          cVar2S32S127P003P015P037nsss(0) <='1';
          else
          cVar2S32S127P003P015P037nsss(0) <='0';
          end if;
        if(cVar1S33S127P064N018P050P048(0)='1' AND  A( 8)='1' AND A( 2)='0' AND A(12)='1' )then
          cVar2S33S127P003N015P014nsss(0) <='1';
          else
          cVar2S33S127P003N015P014nsss(0) <='0';
          end if;
        if(cVar1S34S127P064N018P050P048(0)='1' AND  A( 8)='0' AND D(14)='0' AND A(17)='1' )then
          cVar2S34S127N003P043P004nsss(0) <='1';
          else
          cVar2S34S127N003P043P004nsss(0) <='0';
          end if;
        if(cVar1S35S127P064N018P050P048(0)='1' AND  E(13)='1' )then
          cVar2S35S127P049nsss(0) <='1';
          else
          cVar2S35S127P049nsss(0) <='0';
          end if;
        if(cVar1S37S127P064N018P050N027(0)='1' AND  B( 1)='1' AND B( 0)='1' )then
          cVar2S37S127P035P037nsss(0) <='1';
          else
          cVar2S37S127P035P037nsss(0) <='0';
          end if;
        if(cVar1S38S127P064N018P050N027(0)='1' AND  B( 1)='0' AND E( 8)='1' )then
          cVar2S38S127N035P069nsss(0) <='1';
          else
          cVar2S38S127N035P069nsss(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV3 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar2S0S0P062P011nsss(0)='1'  OR cVar2S1S0P062P011P014nsss(0)='1'  OR cVar2S2S0N062P066nsss(0)='1'  OR cVar2S3S0P058P033nsss(0)='1'  )then
          oVar1S0(0) <='1';
          else
          oVar1S0(0) <='0';
          end if;
        if(cVar2S4S0P058N033P013nsss(0)='1'  OR cVar2S5S0N058P068P066nsss(0)='1'  OR cVar2S6S0N058N068P054nsss(0)='1'  OR cVar2S7S0P036P017nsss(0)='1'  )then
          oVar1S1(0) <='1';
          else
          oVar1S1(0) <='0';
          end if;
        if(cVar2S8S0N036P065P068nsss(0)='1'  OR cVar2S9S0P062nsss(0)='1'  OR cVar2S10S0N062P068P067nsss(0)='1'  OR cVar2S11S0N062N068P060nsss(0)='1'  )then
          oVar1S2(0) <='1';
          else
          oVar1S2(0) <='0';
          end if;
        if(cVar2S12S0P018P062nsss(0)='1'  OR cVar2S13S0P018N062P068nsss(0)='1'  OR cVar2S14S0N018P016P058nsss(0)='1'  OR cVar2S15S0P068P066P012nsss(0)='1'  )then
          oVar1S3(0) <='1';
          else
          oVar1S3(0) <='0';
          end if;
        if(cVar2S16S0N068P067P062nsss(0)='1'  OR cVar2S17S0P060P033nsss(0)='1'  OR cVar2S18S0P068P066nsss(0)='1'  OR cVar2S19S0P068N066P019nsss(0)='1'  )then
          oVar1S4(0) <='1';
          else
          oVar1S4(0) <='0';
          end if;
        if(cVar2S20S0N068P064nsss(0)='1'  OR cVar2S21S0N068N064P060nsss(0)='1'  OR cVar2S22S0P064P016nsss(0)='1'  OR cVar2S23S0P064N016P037nsss(0)='1'  )then
          oVar1S5(0) <='1';
          else
          oVar1S5(0) <='0';
          end if;
        if(cVar2S24S0N064P068P018nsss(0)='1'  OR cVar2S25S0N064N068P060nsss(0)='1'  OR cVar2S26S0P034P062nsss(0)='1'  OR cVar2S27S0P034N062P068nsss(0)='1'  )then
          oVar1S6(0) <='1';
          else
          oVar1S6(0) <='0';
          end if;
        if(cVar2S28S0P015P032nsss(0)='1'  OR cVar2S29S0P015N032P064nsss(0)='1'  OR cVar2S30S0N015P066nsss(0)='1'  OR cVar2S31S0N015N066P062nsss(0)='1'  )then
          oVar1S7(0) <='1';
          else
          oVar1S7(0) <='0';
          end if;
        if(cVar2S32S0P013P030nsss(0)='1'  OR cVar2S33S0P013N030P066nsss(0)='1'  OR cVar2S34S0N013P068P018nsss(0)='1'  OR cVar2S35S0N013N068P064nsss(0)='1'  )then
          oVar1S8(0) <='1';
          else
          oVar1S8(0) <='0';
          end if;
        if(cVar2S36S0P051P028P066nsss(0)='1'  OR cVar2S37S0N051P047P068nsss(0)='1'  )then
          oVar1S9(0) <='1';
          else
          oVar1S9(0) <='0';
          end if;
        if(cVar2S0S1P062nsss(0)='1'  OR cVar2S1S1P062P029nsss(0)='1'  OR cVar2S2S1P029nsss(0)='1'  OR cVar2S3S1N029P028nsss(0)='1'  )then
          oVar1S10(0) <='1';
          else
          oVar1S10(0) <='0';
          end if;
        if(cVar2S4S1P066nsss(0)='1'  OR cVar2S5S1P066P036P019nsss(0)='1'  OR cVar2S6S1P008P064nsss(0)='1'  OR cVar2S7S1N008psss(0)='1'  )then
          oVar1S11(0) <='1';
          else
          oVar1S11(0) <='0';
          end if;
        if(cVar1S8S1P052N050P029nsss(0)='1'  OR cVar2S9S1P054nsss(0)='1'  OR cVar2S10S1P049nsss(0)='1'  OR cVar2S11S1P062nsss(0)='1'  )then
          oVar1S12(0) <='1';
          else
          oVar1S12(0) <='0';
          end if;
        if(cVar2S12S1P062P016nsss(0)='1'  OR cVar1S13S1N052P056P031N063psss(0)='1'  OR cVar2S14S1P003nsss(0)='1'  OR cVar2S15S1P030P012P064nsss(0)='1'  )then
          oVar1S13(0) <='1';
          else
          oVar1S13(0) <='0';
          end if;
        if(cVar2S16S1P030N012P054nsss(0)='1'  OR cVar2S17S1N030P028nsss(0)='1'  OR cVar2S18S1N030N028P027nsss(0)='1'  OR cVar2S19S1P033P069nsss(0)='1'  )then
          oVar1S14(0) <='1';
          else
          oVar1S14(0) <='0';
          end if;
        if(cVar2S20S1P033P069P018nsss(0)='1'  OR cVar2S21S1N033P035nsss(0)='1'  OR cVar2S22S1N033N035P032nsss(0)='1'  OR cVar2S23S1P035P058P064nsss(0)='1'  )then
          oVar1S15(0) <='1';
          else
          oVar1S15(0) <='0';
          end if;
        if(cVar2S24S1P035N058P019nsss(0)='1'  OR cVar2S25S1N035P014P032nsss(0)='1'  OR cVar2S26S1P006nsss(0)='1'  OR cVar2S27S1N006P008nsss(0)='1'  )then
          oVar1S16(0) <='1';
          else
          oVar1S16(0) <='0';
          end if;
        if(cVar2S28S1N006N008P027nsss(0)='1'  OR cVar2S29S1P064P051nsss(0)='1'  OR cVar2S30S1P064N051P035nsss(0)='1'  OR cVar2S31S1N064N068P069nsss(0)='1'  )then
          oVar1S17(0) <='1';
          else
          oVar1S17(0) <='0';
          end if;
        if(cVar2S0S2P043P022nsss(0)='1'  OR cVar2S1S2P043N022P045nsss(0)='1'  OR cVar2S2S2N043P047nsss(0)='1'  OR cVar2S3S2N043P047P049nsss(0)='1'  )then
          oVar1S19(0) <='1';
          else
          oVar1S19(0) <='0';
          end if;
        if(cVar2S4S2P064P015nsss(0)='1'  OR cVar2S5S2P064N015P017nsss(0)='1'  OR cVar2S6S2P064P059P062nsss(0)='1'  OR cVar2S7S2P064P019nsss(0)='1'  )then
          oVar1S20(0) <='1';
          else
          oVar1S20(0) <='0';
          end if;
        if(cVar2S8S2P064N019P012nsss(0)='1'  OR cVar2S9S2P028P018nsss(0)='1'  OR cVar2S10S2N028P039nsss(0)='1'  OR cVar2S11S2P018P019P058nsss(0)='1'  )then
          oVar1S21(0) <='1';
          else
          oVar1S21(0) <='0';
          end if;
        if(cVar2S12S2P018P019psss(0)='1'  OR cVar2S13S2P018P066nsss(0)='1'  OR cVar2S14S2P018P069P065nsss(0)='1'  OR cVar2S15S2P018P069psss(0)='1'  )then
          oVar1S22(0) <='1';
          else
          oVar1S22(0) <='0';
          end if;
        if(cVar2S16S2N018P044nsss(0)='1'  OR cVar1S17S2P068P067P035P031nsss(0)='1'  OR cVar2S18S2P006P014P062nsss(0)='1'  OR cVar2S19S2P060P069P064nsss(0)='1'  )then
          oVar1S23(0) <='1';
          else
          oVar1S23(0) <='0';
          end if;
        if(cVar2S20S2P060P069psss(0)='1'  OR cVar2S21S2P060P058P033nsss(0)='1'  OR cVar2S22S2P064P018nsss(0)='1'  OR cVar2S23S2N064P060P061nsss(0)='1'  )then
          oVar1S24(0) <='1';
          else
          oVar1S24(0) <='0';
          end if;
        if(cVar2S24S2P066P010nsss(0)='1'  OR cVar2S25S2P064P014nsss(0)='1'  OR cVar2S26S2P064N014P060nsss(0)='1'  OR cVar2S27S2P064P017P014nsss(0)='1'  )then
          oVar1S25(0) <='1';
          else
          oVar1S25(0) <='0';
          end if;
        if(cVar2S28S2P064P017P030nsss(0)='1'  OR cVar1S29S2N068N063P051P028nsss(0)='1'  OR cVar2S30S2P026nsss(0)='1'  OR cVar2S31S2N026P029nsss(0)='1'  )then
          oVar1S26(0) <='1';
          else
          oVar1S26(0) <='0';
          end if;
        if(cVar2S32S2N026N029P027nsss(0)='1'  OR cVar2S33S2P050P052nsss(0)='1'  OR cVar2S34S2P050N052P027nsss(0)='1'  OR cVar2S35S2N050P046nsss(0)='1'  )then
          oVar1S27(0) <='1';
          else
          oVar1S27(0) <='0';
          end if;
        if(cVar2S36S2N050N046P060nsss(0)='1'  OR cVar2S37S2P064P037P035nsss(0)='1'  OR cVar2S38S2P064N037P049nsss(0)='1'  OR cVar2S39S2N064P059nsss(0)='1'  )then
          oVar1S28(0) <='1';
          else
          oVar1S28(0) <='0';
          end if;
        if(cVar2S40S2N064N059P055nsss(0)='1'  )then
          oVar1S29(0) <='1';
          else
          oVar1S29(0) <='0';
          end if;
        if(cVar1S0S3P043P022nsss(0)='1'  OR cVar2S1S3P024nsss(0)='1'  OR cVar2S2S3N024P069nsss(0)='1'  OR cVar1S3S3P043N022P007P015psss(0)='1'  )then
          oVar1S30(0) <='1';
          else
          oVar1S30(0) <='0';
          end if;
        if(cVar2S4S3P024P045nsss(0)='1'  OR cVar2S5S3N024P023nsss(0)='1'  OR cVar2S6S3N024N023P016nsss(0)='1'  OR cVar2S7S3P065nsss(0)='1'  )then
          oVar1S31(0) <='1';
          else
          oVar1S31(0) <='0';
          end if;
        if(cVar2S8S3P065P016P069nsss(0)='1'  OR cVar2S9S3P065N016P028nsss(0)='1'  OR cVar2S10S3P014P017P010nsss(0)='1'  OR cVar2S11S3P062P019nsss(0)='1'  )then
          oVar1S32(0) <='1';
          else
          oVar1S32(0) <='0';
          end if;
        if(cVar2S12S3P062P019P018nsss(0)='1'  OR cVar2S13S3P018P069P054nsss(0)='1'  OR cVar2S14S3P018P069P066nsss(0)='1'  OR cVar2S15S3P018P069P034nsss(0)='1'  )then
          oVar1S33(0) <='1';
          else
          oVar1S33(0) <='0';
          end if;
        if(cVar2S16S3P065P069nsss(0)='1'  OR cVar2S17S3P065P069P017nsss(0)='1'  OR cVar2S18S3N065P061P032nsss(0)='1'  OR cVar2S19S3N065N061P049nsss(0)='1'  )then
          oVar1S34(0) <='1';
          else
          oVar1S34(0) <='0';
          end if;
        if(cVar2S20S3P065P064P016nsss(0)='1'  OR cVar2S21S3P065P016P068nsss(0)='1'  OR cVar2S22S3P009nsss(0)='1'  OR cVar2S23S3N009P011nsss(0)='1'  )then
          oVar1S35(0) <='1';
          else
          oVar1S35(0) <='0';
          end if;
        if(cVar2S24S3N009N011P056nsss(0)='1'  OR cVar2S25S3P039P041nsss(0)='1'  OR cVar2S26S3P039N041P020nsss(0)='1'  OR cVar2S27S3N039P047P068nsss(0)='1'  )then
          oVar1S36(0) <='1';
          else
          oVar1S36(0) <='0';
          end if;
        if(cVar1S0S4P044P023P006nsss(0)='1'  OR cVar1S1S4P044P023N006P004nsss(0)='1'  OR cVar2S2S4P046nsss(0)='1'  OR cVar2S3S4P017nsss(0)='1'  )then
          oVar1S38(0) <='1';
          else
          oVar1S38(0) <='0';
          end if;
        if(cVar2S4S4N017P048nsss(0)='1'  OR cVar1S5S4P044N023P025P018psss(0)='1'  OR cVar2S6S4P042nsss(0)='1'  OR cVar2S7S4P011P024nsss(0)='1'  )then
          oVar1S39(0) <='1';
          else
          oVar1S39(0) <='0';
          end if;
        if(cVar2S8S4P011N024P021nsss(0)='1'  OR cVar2S9S4P034P014nsss(0)='1'  OR cVar2S10S4P034P014P033nsss(0)='1'  OR cVar2S11S4P034P015nsss(0)='1'  )then
          oVar1S40(0) <='1';
          else
          oVar1S40(0) <='0';
          end if;
        if(cVar2S12S4P016P010P003nsss(0)='1'  OR cVar2S13S4N016P017nsss(0)='1'  OR cVar2S14S4P036P015nsss(0)='1'  OR cVar2S15S4P011P033P069nsss(0)='1'  )then
          oVar1S41(0) <='1';
          else
          oVar1S41(0) <='0';
          end if;
        if(cVar2S16S4P011P007P026nsss(0)='1'  OR cVar2S17S4P012P030nsss(0)='1'  OR cVar2S18S4P012P030P013nsss(0)='1'  OR cVar2S19S4N012P064P062nsss(0)='1'  )then
          oVar1S42(0) <='1';
          else
          oVar1S42(0) <='0';
          end if;
        if(cVar2S20S4N012N064psss(0)='1'  OR cVar2S21S4P014P035P056nsss(0)='1'  OR cVar2S22S4P069P063nsss(0)='1'  OR cVar2S23S4P069N063P064nsss(0)='1'  )then
          oVar1S43(0) <='1';
          else
          oVar1S43(0) <='0';
          end if;
        if(cVar2S24S4P069P029nsss(0)='1'  OR cVar2S25S4P069N029P059nsss(0)='1'  OR cVar2S26S4P033P069nsss(0)='1'  OR cVar2S27S4N033P035P067nsss(0)='1'  )then
          oVar1S44(0) <='1';
          else
          oVar1S44(0) <='0';
          end if;
        if(cVar2S28S4N033N035P030nsss(0)='1'  )then
          oVar1S45(0) <='1';
          else
          oVar1S45(0) <='0';
          end if;
        if(cVar1S0S5P027P048P052P050nsss(0)='1'  OR cVar2S1S5P008nsss(0)='1'  OR cVar2S2S5N008P019nsss(0)='1'  OR cVar2S3S5N008N019P046nsss(0)='1'  )then
          oVar1S46(0) <='1';
          else
          oVar1S46(0) <='0';
          end if;
        if(cVar1S4S5P027P048P052P009nsss(0)='1'  OR cVar1S5S5P027N048P050P008nsss(0)='1'  OR cVar2S6S5P053P016nsss(0)='1'  OR cVar2S7S5P053P016P034nsss(0)='1'  )then
          oVar1S47(0) <='1';
          else
          oVar1S47(0) <='0';
          end if;
        if(cVar2S8S5P053P018nsss(0)='1'  OR cVar2S9S5P036nsss(0)='1'  OR cVar2S10S5P038nsss(0)='1'  OR cVar2S11S5N038P012P003nsss(0)='1'  )then
          oVar1S48(0) <='1';
          else
          oVar1S48(0) <='0';
          end if;
        if(cVar2S12S5N038N012P051nsss(0)='1'  OR cVar1S13S5N027P043P022nsss(0)='1'  OR cVar2S14S5P063nsss(0)='1'  OR cVar2S15S5P036P066nsss(0)='1'  )then
          oVar1S49(0) <='1';
          else
          oVar1S49(0) <='0';
          end if;
        if(cVar2S16S5P036N066P069nsss(0)='1'  OR cVar2S17S5N036P018P017nsss(0)='1'  OR cVar2S18S5N036N018P039nsss(0)='1'  OR cVar2S19S5P056P019P068nsss(0)='1'  )then
          oVar1S50(0) <='1';
          else
          oVar1S50(0) <='0';
          end if;
        if(cVar2S20S5P056P019P065nsss(0)='1'  OR cVar2S21S5N056P019nsss(0)='1'  OR cVar2S22S5N056N019P016nsss(0)='1'  OR cVar2S23S5P016P013P011nsss(0)='1'  )then
          oVar1S51(0) <='1';
          else
          oVar1S51(0) <='0';
          end if;
        if(cVar2S24S5P016P030P037nsss(0)='1'  OR cVar2S25S5P016N030P051nsss(0)='1'  OR cVar2S26S5P065P018nsss(0)='1'  OR cVar2S27S5P065N018P057nsss(0)='1'  )then
          oVar1S52(0) <='1';
          else
          oVar1S52(0) <='0';
          end if;
        if(cVar2S28S5P065P011P064nsss(0)='1'  OR cVar2S29S5P029P010nsss(0)='1'  OR cVar2S30S5P029N010P051nsss(0)='1'  OR cVar2S31S5N029P064P016nsss(0)='1'  )then
          oVar1S53(0) <='1';
          else
          oVar1S53(0) <='0';
          end if;
        if(cVar2S32S5N029N064P042nsss(0)='1'  )then
          oVar1S54(0) <='1';
          else
          oVar1S54(0) <='0';
          end if;
        if(cVar1S0S6P040P021nsss(0)='1'  OR cVar1S1S6P040N021P023P018nsss(0)='1'  OR cVar2S2S6P005nsss(0)='1'  OR cVar2S3S6P018nsss(0)='1'  )then
          oVar1S55(0) <='1';
          else
          oVar1S55(0) <='0';
          end if;
        if(cVar2S4S6N018P038nsss(0)='1'  OR cVar2S5S6P033P019nsss(0)='1'  OR cVar2S6S6N033P053nsss(0)='1'  OR cVar2S7S6P042nsss(0)='1'  )then
          oVar1S56(0) <='1';
          else
          oVar1S56(0) <='0';
          end if;
        if(cVar2S8S6P048nsss(0)='1'  OR cVar1S9S6N040P025N046P044nsss(0)='1'  OR cVar2S10S6P058P034nsss(0)='1'  OR cVar2S11S6N058P045nsss(0)='1'  )then
          oVar1S57(0) <='1';
          else
          oVar1S57(0) <='0';
          end if;
        if(cVar2S12S6N058N045P047nsss(0)='1'  OR cVar2S13S6P019nsss(0)='1'  OR cVar2S14S6P019P069nsss(0)='1'  OR cVar2S15S6P019P069P066nsss(0)='1'  )then
          oVar1S58(0) <='1';
          else
          oVar1S58(0) <='0';
          end if;
        if(cVar2S16S6P012P011nsss(0)='1'  OR cVar2S17S6P012N011P031nsss(0)='1'  OR cVar2S18S6N012P028P010nsss(0)='1'  OR cVar2S19S6N012N028P035nsss(0)='1'  )then
          oVar1S59(0) <='1';
          else
          oVar1S59(0) <='0';
          end if;
        if(cVar2S20S6P066P058nsss(0)='1'  OR cVar2S21S6P066N058P061nsss(0)='1'  OR cVar2S22S6P066P019P018nsss(0)='1'  OR cVar2S23S6P061P059nsss(0)='1'  )then
          oVar1S60(0) <='1';
          else
          oVar1S60(0) <='0';
          end if;
        if(cVar2S24S6P061N059P051nsss(0)='1'  OR cVar2S25S6N061P050nsss(0)='1'  OR cVar2S26S6N061N050P066nsss(0)='1'  )then
          oVar1S61(0) <='1';
          else
          oVar1S61(0) <='0';
          end if;
        if(cVar1S0S7P066P028P055nsss(0)='1'  OR cVar1S1S7P066P028N055P053nsss(0)='1'  OR cVar2S2S7P010P052nsss(0)='1'  OR cVar2S3S7P010N052P054nsss(0)='1'  )then
          oVar1S62(0) <='1';
          else
          oVar1S62(0) <='0';
          end if;
        if(cVar2S4S7N010P025nsss(0)='1'  OR cVar2S5S7N010N025P034nsss(0)='1'  OR cVar1S6S7P066N028P044P023nsss(0)='1'  OR cVar2S7S7P025P017nsss(0)='1'  )then
          oVar1S63(0) <='1';
          else
          oVar1S63(0) <='0';
          end if;
        if(cVar2S8S7P025N017P018nsss(0)='1'  OR cVar2S9S7N025P006nsss(0)='1'  OR cVar2S10S7N025N006P010nsss(0)='1'  OR cVar2S11S7P021nsss(0)='1'  )then
          oVar1S64(0) <='1';
          else
          oVar1S64(0) <='0';
          end if;
        if(cVar2S12S7N021P023nsss(0)='1'  OR cVar2S13S7N021N023P013nsss(0)='1'  OR cVar2S14S7P069P000nsss(0)='1'  OR cVar2S15S7N069P031nsss(0)='1'  )then
          oVar1S65(0) <='1';
          else
          oVar1S65(0) <='0';
          end if;
        if(cVar2S16S7N069N031P048nsss(0)='1'  OR cVar2S17S7P041nsss(0)='1'  OR cVar2S18S7N041P020P063nsss(0)='1'  OR cVar2S19S7P051P008nsss(0)='1'  )then
          oVar1S66(0) <='1';
          else
          oVar1S66(0) <='0';
          end if;
        if(cVar2S20S7P051N008P037nsss(0)='1'  OR cVar1S21S7P066P065P003P041nsss(0)='1'  OR cVar2S22S7P022nsss(0)='1'  OR cVar2S23S7P064P035nsss(0)='1'  )then
          oVar1S67(0) <='1';
          else
          oVar1S67(0) <='0';
          end if;
        if(cVar2S24S7P017P019nsss(0)='1'  OR cVar2S25S7N017P037P019nsss(0)='1'  OR cVar2S26S7P017P064P063nsss(0)='1'  OR cVar2S27S7P017P069P016nsss(0)='1'  )then
          oVar1S68(0) <='1';
          else
          oVar1S68(0) <='0';
          end if;
        if(cVar2S28S7P016N017P035nsss(0)='1'  OR cVar2S29S7P016P067P034nsss(0)='1'  )then
          oVar1S69(0) <='1';
          else
          oVar1S69(0) <='0';
          end if;
        if(cVar1S0S8P043P045P064nsss(0)='1'  OR cVar2S1S8P044P047nsss(0)='1'  OR cVar2S2S8P044P005nsss(0)='1'  OR cVar2S3S8P044N005P046nsss(0)='1'  )then
          oVar1S70(0) <='1';
          else
          oVar1S70(0) <='0';
          end if;
        if(cVar1S4S8P043N045P005P022nsss(0)='1'  OR cVar2S5S8P018nsss(0)='1'  OR cVar2S6S8P041nsss(0)='1'  OR cVar2S7S8P068P066P011nsss(0)='1'  )then
          oVar1S71(0) <='1';
          else
          oVar1S71(0) <='0';
          end if;
        if(cVar2S8S8N068P014P018nsss(0)='1'  OR cVar1S9S8N043P003P040P021nsss(0)='1'  OR cVar2S10S8P004nsss(0)='1'  OR cVar2S11S8N004P017P037nsss(0)='1'  )then
          oVar1S72(0) <='1';
          else
          oVar1S72(0) <='0';
          end if;
        if(cVar2S12S8N004N017P061nsss(0)='1'  OR cVar2S13S8P049nsss(0)='1'  OR cVar2S14S8N049P051P053nsss(0)='1'  OR cVar2S15S8N049N051P056nsss(0)='1'  )then
          oVar1S73(0) <='1';
          else
          oVar1S73(0) <='0';
          end if;
        if(cVar2S16S8P057P049P055nsss(0)='1'  OR cVar2S17S8N057P025nsss(0)='1'  OR cVar2S18S8N057N025P064nsss(0)='1'  OR cVar1S19S8N043P003P039P020nsss(0)='1'  )then
          oVar1S74(0) <='1';
          else
          oVar1S74(0) <='0';
          end if;
        if(cVar2S20S8P016nsss(0)='1'  OR cVar2S21S8N016P021nsss(0)='1'  OR cVar2S22S8P001P010P058nsss(0)='1'  OR cVar2S23S8P044P018nsss(0)='1'  )then
          oVar1S75(0) <='1';
          else
          oVar1S75(0) <='0';
          end if;
        if(cVar2S24S8N044P021P040nsss(0)='1'  )then
          oVar1S76(0) <='1';
          else
          oVar1S76(0) <='0';
          end if;
        if(cVar2S0S9P066P069nsss(0)='1'  OR cVar2S1S9P066P069P060nsss(0)='1'  OR cVar2S2S9P066P018nsss(0)='1'  OR cVar2S3S9P066N018P069nsss(0)='1'  )then
          oVar1S77(0) <='1';
          else
          oVar1S77(0) <='0';
          end if;
        if(cVar2S4S9P058P067nsss(0)='1'  OR cVar2S5S9P058P067P036nsss(0)='1'  OR cVar2S6S9N058P057nsss(0)='1'  OR cVar2S7S9N058N057P050nsss(0)='1'  )then
          oVar1S78(0) <='1';
          else
          oVar1S78(0) <='0';
          end if;
        if(cVar2S8S9P006P065nsss(0)='1'  OR cVar2S9S9P006N065P060nsss(0)='1'  OR cVar1S10S9P032P015P063P059nsss(0)='1'  OR cVar2S11S9P068P016nsss(0)='1'  )then
          oVar1S79(0) <='1';
          else
          oVar1S79(0) <='0';
          end if;
        if(cVar2S12S9P059P064nsss(0)='1'  OR cVar2S13S9N059P058nsss(0)='1'  OR cVar2S14S9P064P017nsss(0)='1'  OR cVar2S15S9P064P017P013nsss(0)='1'  )then
          oVar1S80(0) <='1';
          else
          oVar1S80(0) <='0';
          end if;
        if(cVar2S16S9N064P061P019nsss(0)='1'  OR cVar2S17S9N064P061P069nsss(0)='1'  OR cVar1S18S9N032P043P045P062nsss(0)='1'  OR cVar2S19S9P022nsss(0)='1'  )then
          oVar1S81(0) <='1';
          else
          oVar1S81(0) <='0';
          end if;
        if(cVar2S20S9N022P049nsss(0)='1'  OR cVar1S21S9N032P043N045P005nsss(0)='1'  OR cVar2S22S9P068P012nsss(0)='1'  OR cVar2S23S9N068P041P013nsss(0)='1'  )then
          oVar1S82(0) <='1';
          else
          oVar1S82(0) <='0';
          end if;
        if(cVar2S24S9N068N041P034nsss(0)='1'  OR cVar1S25S9N032N043P044P023nsss(0)='1'  OR cVar2S26S9P025nsss(0)='1'  OR cVar2S27S9N025P022nsss(0)='1'  )then
          oVar1S83(0) <='1';
          else
          oVar1S83(0) <='0';
          end if;
        if(cVar2S28S9N025N022P009nsss(0)='1'  OR cVar2S29S9P021nsss(0)='1'  OR cVar2S30S9N021P023nsss(0)='1'  OR cVar2S31S9N021N023P041nsss(0)='1'  )then
          oVar1S84(0) <='1';
          else
          oVar1S84(0) <='0';
          end if;
        if(cVar2S32S9P003P033P034nsss(0)='1'  OR cVar2S33S9P003N033psss(0)='1'  OR cVar2S34S9P003P039P020nsss(0)='1'  OR cVar2S35S9P003N039P036nsss(0)='1'  )then
          oVar1S85(0) <='1';
          else
          oVar1S85(0) <='0';
          end if;
        if(cVar2S0S10P066P069nsss(0)='1'  OR cVar2S1S10P066P069P058nsss(0)='1'  OR cVar2S2S10P066P069nsss(0)='1'  OR cVar2S3S10P066N069P014nsss(0)='1'  )then
          oVar1S87(0) <='1';
          else
          oVar1S87(0) <='0';
          end if;
        if(cVar2S4S10P033P047nsss(0)='1'  OR cVar2S5S10P033N047P014nsss(0)='1'  OR cVar2S6S10P006P065nsss(0)='1'  OR cVar2S7S10P006N065P061nsss(0)='1'  )then
          oVar1S88(0) <='1';
          else
          oVar1S88(0) <='0';
          end if;
        if(cVar2S8S10P059nsss(0)='1'  OR cVar2S9S10N059P016nsss(0)='1'  OR cVar2S10S10N059N016P017nsss(0)='1'  OR cVar2S11S10P059P011nsss(0)='1'  )then
          oVar1S89(0) <='1';
          else
          oVar1S89(0) <='0';
          end if;
        if(cVar2S12S10N059P060P017nsss(0)='1'  OR cVar2S13S10P061P066nsss(0)='1'  OR cVar2S14S10P061P068nsss(0)='1'  OR cVar2S15S10P061N068P064nsss(0)='1'  )then
          oVar1S90(0) <='1';
          else
          oVar1S90(0) <='0';
          end if;
        if(cVar1S16S10N032P040P021nsss(0)='1'  OR cVar2S17S10P036P017nsss(0)='1'  OR cVar2S18S10P036N017P068nsss(0)='1'  OR cVar2S19S10N036P044P003nsss(0)='1'  )then
          oVar1S91(0) <='1';
          else
          oVar1S91(0) <='0';
          end if;
        if(cVar2S20S10N036P044P042nsss(0)='1'  OR cVar2S21S10P036P042nsss(0)='1'  OR cVar2S22S10P036N042P018nsss(0)='1'  OR cVar2S23S10P045nsss(0)='1'  )then
          oVar1S92(0) <='1';
          else
          oVar1S92(0) <='0';
          end if;
        if(cVar2S24S10N045P019nsss(0)='1'  OR cVar2S25S10P022P007nsss(0)='1'  OR cVar2S26S10P022N007P005nsss(0)='1'  OR cVar2S27S10N022P024P047nsss(0)='1'  )then
          oVar1S93(0) <='1';
          else
          oVar1S93(0) <='0';
          end if;
        if(cVar2S28S10N022N024P023nsss(0)='1'  OR cVar2S29S10P058P014nsss(0)='1'  OR cVar2S30S10P058N014P012nsss(0)='1'  OR cVar2S31S10N058P059P015nsss(0)='1'  )then
          oVar1S94(0) <='1';
          else
          oVar1S94(0) <='0';
          end if;
        if(cVar2S32S10P044P023nsss(0)='1'  OR cVar2S33S10P044N023P016nsss(0)='1'  OR cVar2S34S10N044P047P068nsss(0)='1'  OR cVar2S35S10N044N047P028nsss(0)='1'  )then
          oVar1S95(0) <='1';
          else
          oVar1S95(0) <='0';
          end if;
        if(cVar1S0S11P027P008P046nsss(0)='1'  OR cVar1S1S11P027P008N046P050nsss(0)='1'  OR cVar2S2S11P069P037nsss(0)='1'  OR cVar2S3S11P046nsss(0)='1'  )then
          oVar1S97(0) <='1';
          else
          oVar1S97(0) <='0';
          end if;
        if(cVar2S4S11P010nsss(0)='1'  OR cVar2S5S11N010P048P006nsss(0)='1'  OR cVar2S6S11P049nsss(0)='1'  OR cVar2S7S11N049P062nsss(0)='1'  )then
          oVar1S98(0) <='1';
          else
          oVar1S98(0) <='0';
          end if;
        if(cVar2S8S11P024P001P049nsss(0)='1'  OR cVar1S9S11N027P039P020P005nsss(0)='1'  OR cVar2S10S11P041P038nsss(0)='1'  OR cVar2S11S11P022nsss(0)='1'  )then
          oVar1S99(0) <='1';
          else
          oVar1S99(0) <='0';
          end if;
        if(cVar2S12S11N022P023nsss(0)='1'  OR cVar2S13S11N022N023P019nsss(0)='1'  OR cVar2S14S11P066P019P015nsss(0)='1'  OR cVar2S15S11P035P066nsss(0)='1'  )then
          oVar1S100(0) <='1';
          else
          oVar1S100(0) <='0';
          end if;
        if(cVar2S16S11P035P066P015nsss(0)='1'  OR cVar2S17S11P068P065nsss(0)='1'  OR cVar2S18S11N068P054P057nsss(0)='1'  OR cVar2S19S11N068N054P035nsss(0)='1'  )then
          oVar1S101(0) <='1';
          else
          oVar1S101(0) <='0';
          end if;
        if(cVar2S20S11P038nsss(0)='1'  OR cVar2S21S11N038P042nsss(0)='1'  OR cVar2S22S11P013P065P017nsss(0)='1'  OR cVar2S23S11P013P031nsss(0)='1'  )then
          oVar1S102(0) <='1';
          else
          oVar1S102(0) <='0';
          end if;
        if(cVar2S0S12P062nsss(0)='1'  OR cVar2S1S12P062P018P013nsss(0)='1'  OR cVar2S2S12P062N018P037nsss(0)='1'  OR cVar2S3S12P063P069nsss(0)='1'  )then
          oVar1S104(0) <='1';
          else
          oVar1S104(0) <='0';
          end if;
        if(cVar2S4S12N063P055nsss(0)='1'  OR cVar2S5S12N063N055P046nsss(0)='1'  OR cVar2S6S12P014P034nsss(0)='1'  OR cVar2S7S12P014P034P048nsss(0)='1'  )then
          oVar1S105(0) <='1';
          else
          oVar1S105(0) <='0';
          end if;
        if(cVar2S8S12P014P056P017nsss(0)='1'  OR cVar2S9S12P014N056P064nsss(0)='1'  OR cVar2S10S12P034P017P060nsss(0)='1'  OR cVar2S11S12P034N017psss(0)='1'  )then
          oVar1S106(0) <='1';
          else
          oVar1S106(0) <='0';
          end if;
        if(cVar2S12S12N034P037nsss(0)='1'  OR cVar2S13S12N034N037P033nsss(0)='1'  OR cVar2S14S12P013P012nsss(0)='1'  OR cVar2S15S12P013P012P018nsss(0)='1'  )then
          oVar1S107(0) <='1';
          else
          oVar1S107(0) <='0';
          end if;
        if(cVar2S16S12P013P059P015nsss(0)='1'  OR cVar2S17S12P013N059P036nsss(0)='1'  OR cVar2S18S12P064P033P012nsss(0)='1'  OR cVar2S19S12P064P017P019nsss(0)='1'  )then
          oVar1S108(0) <='1';
          else
          oVar1S108(0) <='0';
          end if;
        if(cVar2S20S12P055nsss(0)='1'  OR cVar2S21S12N055P069P037nsss(0)='1'  OR cVar2S22S12P036P051nsss(0)='1'  OR cVar2S23S12N036P053P037nsss(0)='1'  )then
          oVar1S109(0) <='1';
          else
          oVar1S109(0) <='0';
          end if;
        if(cVar2S24S12P054nsss(0)='1'  OR cVar2S25S12N054P012P062nsss(0)='1'  OR cVar2S26S12N054P012P058nsss(0)='1'  OR cVar2S27S12P064P003P017nsss(0)='1'  )then
          oVar1S110(0) <='1';
          else
          oVar1S110(0) <='0';
          end if;
        if(cVar2S28S12P064P032P019nsss(0)='1'  OR cVar2S29S12P064N032P059nsss(0)='1'  OR cVar2S30S12P055P012P001nsss(0)='1'  OR cVar2S31S12P055P012P064nsss(0)='1'  )then
          oVar1S111(0) <='1';
          else
          oVar1S111(0) <='0';
          end if;
        if(cVar2S32S12P064P034P010nsss(0)='1'  OR cVar2S33S12P005P009nsss(0)='1'  OR cVar2S34S12P016P018nsss(0)='1'  OR cVar2S35S12P016P018nsss(0)='1'  )then
          oVar1S112(0) <='1';
          else
          oVar1S112(0) <='0';
          end if;
        if(cVar2S36S12P010P036P017nsss(0)='1'  OR cVar2S37S12P010P036P017nsss(0)='1'  OR cVar2S38S12P065P064nsss(0)='1'  )then
          oVar1S113(0) <='1';
          else
          oVar1S113(0) <='0';
          end if;
        if(cVar2S0S13P012nsss(0)='1'  OR cVar2S1S13P012P052nsss(0)='1'  OR cVar2S2S13P031P028nsss(0)='1'  OR cVar2S3S13P031P028P011nsss(0)='1'  )then
          oVar1S114(0) <='1';
          else
          oVar1S114(0) <='0';
          end if;
        if(cVar2S4S13P031P012nsss(0)='1'  OR cVar2S5S13P048P040nsss(0)='1'  OR cVar2S6S13N048P025nsss(0)='1'  OR cVar2S7S13N048N025P023nsss(0)='1'  )then
          oVar1S115(0) <='1';
          else
          oVar1S115(0) <='0';
          end if;
        if(cVar2S8S13P030P012P066nsss(0)='1'  OR cVar2S9S13P030N012P036nsss(0)='1'  OR cVar2S10S13N030psss(0)='1'  OR cVar2S11S13P001P065P024nsss(0)='1'  )then
          oVar1S116(0) <='1';
          else
          oVar1S116(0) <='0';
          end if;
        if(cVar2S12S13P001P065P034nsss(0)='1'  OR cVar2S13S13P055nsss(0)='1'  OR cVar2S14S13N055P019P058nsss(0)='1'  OR cVar2S15S13N055N019P056nsss(0)='1'  )then
          oVar1S117(0) <='1';
          else
          oVar1S117(0) <='0';
          end if;
        if(cVar2S16S13P049P003nsss(0)='1'  OR cVar2S17S13P049P003P068nsss(0)='1'  OR cVar2S18S13P009P065P066nsss(0)='1'  OR cVar2S19S13P009P026P018nsss(0)='1'  )then
          oVar1S118(0) <='1';
          else
          oVar1S118(0) <='0';
          end if;
        if(cVar2S20S13P009N026P027nsss(0)='1'  OR cVar2S21S13P069P062nsss(0)='1'  OR cVar2S22S13P069N062P036nsss(0)='1'  OR cVar2S23S13P069P058P057nsss(0)='1'  )then
          oVar1S119(0) <='1';
          else
          oVar1S119(0) <='0';
          end if;
        if(cVar2S24S13P032P066nsss(0)='1'  OR cVar2S25S13N032P014P037nsss(0)='1'  OR cVar2S26S13P065P015P011nsss(0)='1'  OR cVar2S27S13P065N015P012nsss(0)='1'  )then
          oVar1S120(0) <='1';
          else
          oVar1S120(0) <='0';
          end if;
        if(cVar2S28S13N065P067P036nsss(0)='1'  OR cVar2S29S13P065P037P036nsss(0)='1'  OR cVar2S30S13P065N037P015nsss(0)='1'  OR cVar2S31S13P065P014P016nsss(0)='1'  )then
          oVar1S121(0) <='1';
          else
          oVar1S121(0) <='0';
          end if;
        if(cVar2S32S13P065N014P060nsss(0)='1'  OR cVar1S33S13P064P010P032P061nsss(0)='1'  OR cVar2S34S13P030P015nsss(0)='1'  OR cVar2S35S13P030N015P035nsss(0)='1'  )then
          oVar1S122(0) <='1';
          else
          oVar1S122(0) <='0';
          end if;
        if(cVar2S36S13N030P055P029nsss(0)='1'  )then
          oVar1S123(0) <='1';
          else
          oVar1S123(0) <='0';
          end if;
        if(cVar1S0S14P030P057P063nsss(0)='1'  OR cVar2S1S14P011P018nsss(0)='1'  OR cVar2S2S14P011P018P068nsss(0)='1'  OR cVar2S3S14N011P064nsss(0)='1'  )then
          oVar1S124(0) <='1';
          else
          oVar1S124(0) <='0';
          end if;
        if(cVar2S4S14N011P064P037nsss(0)='1'  OR cVar2S5S14P018nsss(0)='1'  OR cVar2S6S14N018P037nsss(0)='1'  OR cVar2S7S14N018N037P059nsss(0)='1'  )then
          oVar1S125(0) <='1';
          else
          oVar1S125(0) <='0';
          end if;
        if(cVar2S8S14P008P019nsss(0)='1'  OR cVar2S9S14P008P019P018nsss(0)='1'  OR cVar2S10S14P069P012nsss(0)='1'  OR cVar2S11S14P013P062nsss(0)='1'  )then
          oVar1S126(0) <='1';
          else
          oVar1S126(0) <='0';
          end if;
        if(cVar2S12S14N013P034P011nsss(0)='1'  OR cVar2S13S14P029N062P051nsss(0)='1'  OR cVar2S14S14P064nsss(0)='1'  OR cVar2S15S14P064P017nsss(0)='1'  )then
          oVar1S127(0) <='1';
          else
          oVar1S127(0) <='0';
          end if;
        if(cVar2S16S14P062P052nsss(0)='1'  OR cVar2S17S14P062N052P054nsss(0)='1'  OR cVar2S18S14P050nsss(0)='1'  OR cVar2S19S14P050P014nsss(0)='1'  )then
          oVar1S128(0) <='1';
          else
          oVar1S128(0) <='0';
          end if;
        if(cVar2S20S14P050N014P018nsss(0)='1'  OR cVar2S21S14P052P008nsss(0)='1'  OR cVar2S22S14P052N008P012nsss(0)='1'  OR cVar2S23S14P000P034P040nsss(0)='1'  )then
          oVar1S129(0) <='1';
          else
          oVar1S129(0) <='0';
          end if;
        if(cVar2S24S14P000P034P017nsss(0)='1'  OR cVar2S25S14P025P048nsss(0)='1'  OR cVar2S26S14N025P027nsss(0)='1'  OR cVar2S27S14N025N027P062nsss(0)='1'  )then
          oVar1S130(0) <='1';
          else
          oVar1S130(0) <='0';
          end if;
        if(cVar2S28S14P012P052P009nsss(0)='1'  OR cVar2S29S14P012P052P027nsss(0)='1'  OR cVar2S30S14P012P031P062nsss(0)='1'  OR cVar2S31S14P040P021nsss(0)='1'  )then
          oVar1S131(0) <='1';
          else
          oVar1S131(0) <='0';
          end if;
        if(cVar2S32S14P040N021P013nsss(0)='1'  OR cVar2S33S14N040P032P013nsss(0)='1'  )then
          oVar1S132(0) <='1';
          else
          oVar1S132(0) <='0';
          end if;
        if(cVar1S0S15P037P039P020nsss(0)='1'  OR cVar1S1S15P037P039N020P022nsss(0)='1'  OR cVar2S2S15P021P038nsss(0)='1'  OR cVar2S3S15N021P035P062nsss(0)='1'  )then
          oVar1S133(0) <='1';
          else
          oVar1S133(0) <='0';
          end if;
        if(cVar2S4S15N021N035P026nsss(0)='1'  OR cVar2S5S15P046nsss(0)='1'  OR cVar2S6S15P046P009nsss(0)='1'  OR cVar2S7S15P008P046nsss(0)='1'  )then
          oVar1S134(0) <='1';
          else
          oVar1S134(0) <='0';
          end if;
        if(cVar2S8S15N008P049P018nsss(0)='1'  OR cVar2S9S15P009P013P007nsss(0)='1'  OR cVar2S10S15P009P013P011nsss(0)='1'  OR cVar2S11S15N009P068P006nsss(0)='1'  )then
          oVar1S135(0) <='1';
          else
          oVar1S135(0) <='0';
          end if;
        if(cVar2S12S15P008P067P058nsss(0)='1'  OR cVar2S13S15P008N067P058nsss(0)='1'  OR cVar2S14S15P008P052P029nsss(0)='1'  OR cVar1S15S15P037P030P057P016nsss(0)='1'  )then
          oVar1S136(0) <='1';
          else
          oVar1S136(0) <='0';
          end if;
        if(cVar2S16S15P069nsss(0)='1'  OR cVar2S17S15N069P019P056nsss(0)='1'  OR cVar2S18S15N069N019P013nsss(0)='1'  OR cVar2S19S15P018nsss(0)='1'  )then
          oVar1S137(0) <='1';
          else
          oVar1S137(0) <='0';
          end if;
        if(cVar2S20S15N018P017nsss(0)='1'  OR cVar2S21S15P047P026nsss(0)='1'  OR cVar2S22S15P047N026P018nsss(0)='1'  OR cVar2S23S15N047P058P017nsss(0)='1'  )then
          oVar1S138(0) <='1';
          else
          oVar1S138(0) <='0';
          end if;
        if(cVar2S24S15P047P031P061nsss(0)='1'  OR cVar2S25S15P047N031P029nsss(0)='1'  OR cVar2S26S15P047P007P024nsss(0)='1'  OR cVar2S27S15P018nsss(0)='1'  )then
          oVar1S139(0) <='1';
          else
          oVar1S139(0) <='0';
          end if;
        if(cVar2S28S15N018P068nsss(0)='1'  OR cVar2S29S15P028P018P053nsss(0)='1'  OR cVar2S30S15N028P069P018nsss(0)='1'  )then
          oVar1S140(0) <='1';
          else
          oVar1S140(0) <='0';
          end if;
        if(cVar1S0S16P043P022P007nsss(0)='1'  OR cVar2S1S16P068nsss(0)='1'  OR cVar2S2S16P068P004nsss(0)='1'  OR cVar2S3S16P069P005nsss(0)='1'  )then
          oVar1S141(0) <='1';
          else
          oVar1S141(0) <='0';
          end if;
        if(cVar2S4S16P069N005P062nsss(0)='1'  OR cVar1S5S16P043N022P062P016nsss(0)='1'  OR cVar2S6S16P019nsss(0)='1'  OR cVar2S7S16P068P024nsss(0)='1'  )then
          oVar1S142(0) <='1';
          else
          oVar1S142(0) <='0';
          end if;
        if(cVar2S8S16P068psss(0)='1'  OR cVar2S9S16P049P044P048nsss(0)='1'  OR cVar2S10S16P055nsss(0)='1'  OR cVar2S11S16P011P013nsss(0)='1'  )then
          oVar1S143(0) <='1';
          else
          oVar1S143(0) <='0';
          end if;
        if(cVar2S12S16P011P013P066nsss(0)='1'  OR cVar2S13S16N011P018nsss(0)='1'  OR cVar2S14S16N011N018P013nsss(0)='1'  OR cVar2S15S16P014P061nsss(0)='1'  )then
          oVar1S144(0) <='1';
          else
          oVar1S144(0) <='0';
          end if;
        if(cVar2S16S16P014N061P054nsss(0)='1'  OR cVar2S17S16P014P058P066nsss(0)='1'  OR cVar2S18S16P014N058P053nsss(0)='1'  OR cVar2S19S16P013P012nsss(0)='1'  )then
          oVar1S145(0) <='1';
          else
          oVar1S145(0) <='0';
          end if;
        if(cVar2S20S16P005nsss(0)='1'  OR cVar2S21S16N005P041nsss(0)='1'  OR cVar2S22S16P013P022nsss(0)='1'  OR cVar2S23S16P013N022P053nsss(0)='1'  )then
          oVar1S146(0) <='1';
          else
          oVar1S146(0) <='0';
          end if;
        if(cVar2S24S16P033P054nsss(0)='1'  OR cVar2S25S16P033P054P063nsss(0)='1'  OR cVar2S26S16P033P069P015nsss(0)='1'  OR cVar2S27S16P033N069P027nsss(0)='1'  )then
          oVar1S147(0) <='1';
          else
          oVar1S147(0) <='0';
          end if;
        if(cVar2S28S16P044P023nsss(0)='1'  OR cVar2S29S16P044N023P022nsss(0)='1'  OR cVar2S30S16N044P029nsss(0)='1'  OR cVar2S31S16N044N029P027nsss(0)='1'  )then
          oVar1S148(0) <='1';
          else
          oVar1S148(0) <='0';
          end if;
        if(cVar2S0S17P059P063P067nsss(0)='1'  OR cVar2S1S17P059N063psss(0)='1'  OR cVar2S2S17N059P058P030nsss(0)='1'  OR cVar2S3S17P033P018nsss(0)='1'  )then
          oVar1S150(0) <='1';
          else
          oVar1S150(0) <='0';
          end if;
        if(cVar2S4S17P033N018P014nsss(0)='1'  OR cVar2S5S17P036P018nsss(0)='1'  OR cVar2S6S17P036N018P014nsss(0)='1'  OR cVar2S7S17N036P013P059nsss(0)='1'  )then
          oVar1S151(0) <='1';
          else
          oVar1S151(0) <='0';
          end if;
        if(cVar2S8S17P036P012P061nsss(0)='1'  OR cVar2S9S17P017P054nsss(0)='1'  OR cVar2S10S17P017P054P069nsss(0)='1'  OR cVar2S11S17P017P018P062nsss(0)='1'  )then
          oVar1S152(0) <='1';
          else
          oVar1S152(0) <='0';
          end if;
        if(cVar2S12S17P017P018P036nsss(0)='1'  OR cVar2S13S17P017P068nsss(0)='1'  OR cVar2S14S17P017P068P015nsss(0)='1'  OR cVar2S15S17N017P026P004nsss(0)='1'  )then
          oVar1S153(0) <='1';
          else
          oVar1S153(0) <='0';
          end if;
        if(cVar2S16S17N017N026P018nsss(0)='1'  OR cVar2S17S17P014P064P006nsss(0)='1'  OR cVar2S18S17P014P064nsss(0)='1'  OR cVar2S19S17P014N064P068nsss(0)='1'  )then
          oVar1S154(0) <='1';
          else
          oVar1S154(0) <='0';
          end if;
        if(cVar2S20S17P010P033nsss(0)='1'  OR cVar2S21S17P010N033P008nsss(0)='1'  OR cVar2S22S17N010P039nsss(0)='1'  OR cVar2S23S17N010N039P031nsss(0)='1'  )then
          oVar1S155(0) <='1';
          else
          oVar1S155(0) <='0';
          end if;
        if(cVar1S24S17P001P015P041nsss(0)='1'  OR cVar2S25S17P068P067P037nsss(0)='1'  OR cVar2S26S17P068N067P019nsss(0)='1'  OR cVar2S27S17N068P014P013nsss(0)='1'  )then
          oVar1S156(0) <='1';
          else
          oVar1S156(0) <='0';
          end if;
        if(cVar2S28S17N068N014P018nsss(0)='1'  OR cVar2S29S17P017nsss(0)='1'  OR cVar2S30S17P017P016P014nsss(0)='1'  OR cVar2S31S17P037nsss(0)='1'  )then
          oVar1S157(0) <='1';
          else
          oVar1S157(0) <='0';
          end if;
        if(cVar2S32S17P005P053P026nsss(0)='1'  )then
          oVar1S158(0) <='1';
          else
          oVar1S158(0) <='0';
          end if;
        if(cVar2S0S18P012P014nsss(0)='1'  OR cVar2S1S18P012P014P056nsss(0)='1'  OR cVar2S2S18N012P064P060nsss(0)='1'  OR cVar2S3S18N012N064P028nsss(0)='1'  )then
          oVar1S159(0) <='1';
          else
          oVar1S159(0) <='0';
          end if;
        if(cVar2S4S18P053P050nsss(0)='1'  OR cVar2S5S18P053P050P026nsss(0)='1'  OR cVar2S6S18N053P036P034nsss(0)='1'  OR cVar2S7S18N053N036psss(0)='1'  )then
          oVar1S160(0) <='1';
          else
          oVar1S160(0) <='0';
          end if;
        if(cVar2S8S18P036P063nsss(0)='1'  OR cVar2S9S18N036P019P010nsss(0)='1'  OR cVar2S10S18P064P018nsss(0)='1'  OR cVar2S11S18N064P032P014nsss(0)='1'  )then
          oVar1S161(0) <='1';
          else
          oVar1S161(0) <='0';
          end if;
        if(cVar2S12S18P068P036P010nsss(0)='1'  OR cVar2S13S18P068P036P011nsss(0)='1'  OR cVar2S14S18N068P045nsss(0)='1'  OR cVar2S15S18N068N045P066nsss(0)='1'  )then
          oVar1S162(0) <='1';
          else
          oVar1S162(0) <='0';
          end if;
        if(cVar2S16S18P033P066nsss(0)='1'  OR cVar2S17S18N033P002P032nsss(0)='1'  OR cVar2S18S18P069nsss(0)='1'  OR cVar2S19S18N069P047nsss(0)='1'  )then
          oVar1S163(0) <='1';
          else
          oVar1S163(0) <='0';
          end if;
        if(cVar2S20S18P018P055P069nsss(0)='1'  OR cVar2S21S18P018P055P013nsss(0)='1'  OR cVar2S22S18N018P017P069nsss(0)='1'  OR cVar2S23S18P018P055P063nsss(0)='1'  )then
          oVar1S164(0) <='1';
          else
          oVar1S164(0) <='0';
          end if;
        if(cVar2S24S18P018P066P062nsss(0)='1'  OR cVar2S25S18P018P066P012nsss(0)='1'  OR cVar2S26S18P066P010nsss(0)='1'  OR cVar2S27S18P066P010P018nsss(0)='1'  )then
          oVar1S165(0) <='1';
          else
          oVar1S165(0) <='0';
          end if;
        if(cVar2S28S18N066P059P033nsss(0)='1'  OR cVar2S29S18P014P028nsss(0)='1'  OR cVar2S30S18P014P034P012nsss(0)='1'  OR cVar2S31S18P015P016P063nsss(0)='1'  )then
          oVar1S166(0) <='1';
          else
          oVar1S166(0) <='0';
          end if;
        if(cVar2S32S18P015N016P068nsss(0)='1'  OR cVar1S33S18P067P007P049nsss(0)='1'  OR cVar2S34S18P017P065P037nsss(0)='1'  )then
          oVar1S167(0) <='1';
          else
          oVar1S167(0) <='0';
          end if;
        if(cVar2S0S19P054nsss(0)='1'  OR cVar2S1S19P054P013nsss(0)='1'  OR cVar2S2S19P056P062nsss(0)='1'  OR cVar2S3S19P056P062P037nsss(0)='1'  )then
          oVar1S168(0) <='1';
          else
          oVar1S168(0) <='0';
          end if;
        if(cVar2S4S19N056P055P013nsss(0)='1'  OR cVar2S5S19P056nsss(0)='1'  OR cVar2S6S19N056P016nsss(0)='1'  OR cVar2S7S19P069P062P065nsss(0)='1'  )then
          oVar1S169(0) <='1';
          else
          oVar1S169(0) <='0';
          end if;
        if(cVar2S8S19P069N062psss(0)='1'  OR cVar2S9S19P069P055nsss(0)='1'  OR cVar2S10S19P037P018nsss(0)='1'  OR cVar2S11S19P037N018P016nsss(0)='1'  )then
          oVar1S170(0) <='1';
          else
          oVar1S170(0) <='0';
          end if;
        if(cVar2S12S19P014nsss(0)='1'  OR cVar2S13S19N014P010nsss(0)='1'  OR cVar2S14S19P011P069P037nsss(0)='1'  OR cVar2S15S19N011P056P015nsss(0)='1'  )then
          oVar1S171(0) <='1';
          else
          oVar1S171(0) <='0';
          end if;
        if(cVar2S16S19P010P054P060nsss(0)='1'  OR cVar2S17S19P010P054P033nsss(0)='1'  OR cVar2S18S19P010P014P006nsss(0)='1'  OR cVar2S19S19P010P014P060nsss(0)='1'  )then
          oVar1S172(0) <='1';
          else
          oVar1S172(0) <='0';
          end if;
        if(cVar2S20S19P035P009P008nsss(0)='1'  OR cVar2S21S19P035P059nsss(0)='1'  OR cVar2S22S19P059P010P009nsss(0)='1'  OR cVar2S23S19P035P009nsss(0)='1'  )then
          oVar1S173(0) <='1';
          else
          oVar1S173(0) <='0';
          end if;
        if(cVar2S24S19N035P016P013nsss(0)='1'  OR cVar2S25S19P022nsss(0)='1'  OR cVar2S26S19N022P024nsss(0)='1'  OR cVar2S27S19N022N024P013nsss(0)='1'  )then
          oVar1S174(0) <='1';
          else
          oVar1S174(0) <='0';
          end if;
        if(cVar2S28S19P008P009nsss(0)='1'  OR cVar2S29S19P008N009P043nsss(0)='1'  OR cVar2S30S19N008P066nsss(0)='1'  OR cVar2S31S19P051P026P012nsss(0)='1'  )then
          oVar1S175(0) <='1';
          else
          oVar1S175(0) <='0';
          end if;
        if(cVar2S32S19P051N026P066nsss(0)='1'  OR cVar2S33S19N051P028P019nsss(0)='1'  OR cVar2S34S19P039P020nsss(0)='1'  OR cVar2S35S19P039N020P022nsss(0)='1'  )then
          oVar1S176(0) <='1';
          else
          oVar1S176(0) <='0';
          end if;
        if(cVar2S36S19N039P030P011nsss(0)='1'  )then
          oVar1S177(0) <='1';
          else
          oVar1S177(0) <='0';
          end if;
        if(cVar2S0S20P006P019nsss(0)='1'  OR cVar2S1S20P006P019P055nsss(0)='1'  OR cVar2S2S20P006P018nsss(0)='1'  OR cVar2S3S20P005P015nsss(0)='1'  )then
          oVar1S178(0) <='1';
          else
          oVar1S178(0) <='0';
          end if;
        if(cVar2S4S20P005P015P037nsss(0)='1'  OR cVar2S5S20P003P068P019nsss(0)='1'  OR cVar2S6S20P003P068psss(0)='1'  OR cVar2S7S20P003P059nsss(0)='1'  )then
          oVar1S179(0) <='1';
          else
          oVar1S179(0) <='0';
          end if;
        if(cVar2S8S20P014nsss(0)='1'  OR cVar2S9S20N014P019P035nsss(0)='1'  OR cVar2S10S20N014N019P054nsss(0)='1'  OR cVar2S11S20P014nsss(0)='1'  )then
          oVar1S180(0) <='1';
          else
          oVar1S180(0) <='0';
          end if;
        if(cVar2S12S20P066P010nsss(0)='1'  OR cVar2S13S20P007nsss(0)='1'  OR cVar2S14S20N007P009nsss(0)='1'  OR cVar2S15S20N007N009P069nsss(0)='1'  )then
          oVar1S181(0) <='1';
          else
          oVar1S181(0) <='0';
          end if;
        if(cVar2S16S20P010P046nsss(0)='1'  OR cVar2S17S20P010N046P064nsss(0)='1'  OR cVar2S18S20P010P025nsss(0)='1'  OR cVar2S19S20P015P059nsss(0)='1'  )then
          oVar1S182(0) <='1';
          else
          oVar1S182(0) <='0';
          end if;
        if(cVar2S20S20P015P059P034nsss(0)='1'  OR cVar2S21S20P015P061P066nsss(0)='1'  OR cVar2S22S20P015N061P060nsss(0)='1'  OR cVar2S23S20P015P061nsss(0)='1'  )then
          oVar1S183(0) <='1';
          else
          oVar1S183(0) <='0';
          end if;
        if(cVar2S24S20P015N061P018nsss(0)='1'  OR cVar2S25S20N015P016P061nsss(0)='1'  OR cVar2S26S20N015N016P010nsss(0)='1'  OR cVar2S27S20P050P042P013nsss(0)='1'  )then
          oVar1S184(0) <='1';
          else
          oVar1S184(0) <='0';
          end if;
        if(cVar2S28S20P050N042P037nsss(0)='1'  OR cVar2S29S20P050P008P067nsss(0)='1'  OR cVar2S30S20P064P067P034nsss(0)='1'  OR cVar2S31S20P064P067P011nsss(0)='1'  )then
          oVar1S185(0) <='1';
          else
          oVar1S185(0) <='0';
          end if;
        if(cVar2S32S20P030nsss(0)='1'  OR cVar2S33S20N030P067nsss(0)='1'  OR cVar2S34S20P050P013nsss(0)='1'  )then
          oVar1S186(0) <='1';
          else
          oVar1S186(0) <='0';
          end if;
        if(cVar2S0S21P035P046nsss(0)='1'  OR cVar2S1S21P035P046P049nsss(0)='1'  OR cVar2S2S21P035psss(0)='1'  OR cVar1S3S21P024P047P066P007nsss(0)='1'  )then
          oVar1S187(0) <='1';
          else
          oVar1S187(0) <='0';
          end if;
        if(cVar2S4S21P016P018nsss(0)='1'  OR cVar2S5S21P016nsss(0)='1'  OR cVar2S6S21N016P044nsss(0)='1'  OR cVar2S7S21P046P036nsss(0)='1'  )then
          oVar1S188(0) <='1';
          else
          oVar1S188(0) <='0';
          end if;
        if(cVar2S8S21N046P061P033nsss(0)='1'  OR cVar2S9S21N046N061P044nsss(0)='1'  OR cVar1S10S21P024N047P010P032nsss(0)='1'  OR cVar2S11S21P037P017nsss(0)='1'  )then
          oVar1S189(0) <='1';
          else
          oVar1S189(0) <='0';
          end if;
        if(cVar2S12S21P011nsss(0)='1'  OR cVar2S13S21P011P013nsss(0)='1'  OR cVar2S14S21P011P013P018nsss(0)='1'  OR cVar2S15S21N011P055P013nsss(0)='1'  )then
          oVar1S190(0) <='1';
          else
          oVar1S190(0) <='0';
          end if;
        if(cVar2S16S21N011P055psss(0)='1'  OR cVar2S17S21P014P040nsss(0)='1'  OR cVar2S18S21P014N040P056nsss(0)='1'  OR cVar2S19S21P014P012P011nsss(0)='1'  )then
          oVar1S191(0) <='1';
          else
          oVar1S191(0) <='0';
          end if;
        if(cVar2S20S21P014N012P060nsss(0)='1'  OR cVar2S21S21P034P012P008nsss(0)='1'  OR cVar2S22S21P034N012P059nsss(0)='1'  OR cVar2S23S21P034P007P033nsss(0)='1'  )then
          oVar1S192(0) <='1';
          else
          oVar1S192(0) <='0';
          end if;
        if(cVar2S24S21P067P056nsss(0)='1'  OR cVar2S25S21P067N056P057nsss(0)='1'  OR cVar2S26S21P067P068P012nsss(0)='1'  OR cVar2S27S21P017P014P008nsss(0)='1'  )then
          oVar1S193(0) <='1';
          else
          oVar1S193(0) <='0';
          end if;
        if(cVar2S28S21P017N014psss(0)='1'  OR cVar2S29S21N017P015P061nsss(0)='1'  OR cVar2S30S21N017N015P067nsss(0)='1'  OR cVar2S31S21P028P062P008nsss(0)='1'  )then
          oVar1S194(0) <='1';
          else
          oVar1S194(0) <='0';
          end if;
        if(cVar2S32S21P028P062P011nsss(0)='1'  OR cVar2S33S21N028P029P019nsss(0)='1'  )then
          oVar1S195(0) <='1';
          else
          oVar1S195(0) <='0';
          end if;
        if(cVar1S0S22P024P047P066nsss(0)='1'  OR cVar2S1S22P045P019nsss(0)='1'  OR cVar2S2S22P045P019P037nsss(0)='1'  OR cVar2S3S22P043nsss(0)='1'  )then
          oVar1S196(0) <='1';
          else
          oVar1S196(0) <='0';
          end if;
        if(cVar2S4S22N043P046P036nsss(0)='1'  OR cVar2S5S22N043N046P017nsss(0)='1'  OR cVar1S6S22P024N047P010P032nsss(0)='1'  OR cVar2S7S22P037P015nsss(0)='1'  )then
          oVar1S197(0) <='1';
          else
          oVar1S197(0) <='0';
          end if;
        if(cVar2S8S22P007nsss(0)='1'  OR cVar2S9S22N007P005nsss(0)='1'  OR cVar2S10S22N007N005P042nsss(0)='1'  OR cVar2S11S22P036P069nsss(0)='1'  )then
          oVar1S198(0) <='1';
          else
          oVar1S198(0) <='0';
          end if;
        if(cVar2S12S22N036psss(0)='1'  OR cVar2S13S22P066P010nsss(0)='1'  OR cVar2S14S22P066P037P055nsss(0)='1'  OR cVar2S15S22P031P012P062nsss(0)='1'  )then
          oVar1S199(0) <='1';
          else
          oVar1S199(0) <='0';
          end if;
        if(cVar2S16S22P031N012P063nsss(0)='1'  OR cVar2S17S22N031P069P063nsss(0)='1'  OR cVar2S18S22N031N069P030nsss(0)='1'  OR cVar2S19S22P036P037nsss(0)='1'  )then
          oVar1S200(0) <='1';
          else
          oVar1S200(0) <='0';
          end if;
        if(cVar2S20S22P036P037P058nsss(0)='1'  OR cVar2S21S22N036P019P062nsss(0)='1'  OR cVar2S22S22N036P019P058nsss(0)='1'  OR cVar2S23S22P003nsss(0)='1'  )then
          oVar1S201(0) <='1';
          else
          oVar1S201(0) <='0';
          end if;
        if(cVar2S24S22N003P033P014nsss(0)='1'  OR cVar2S25S22P017P046P068nsss(0)='1'  OR cVar2S26S22P017P036P018nsss(0)='1'  OR cVar2S27S22P017P036P014nsss(0)='1'  )then
          oVar1S202(0) <='1';
          else
          oVar1S202(0) <='0';
          end if;
        if(cVar2S28S22P062P018P055nsss(0)='1'  OR cVar2S29S22P062N018P023nsss(0)='1'  OR cVar2S30S22P062P019P016nsss(0)='1'  )then
          oVar1S203(0) <='1';
          else
          oVar1S203(0) <='0';
          end if;
        if(cVar1S0S23P024P047P066P063nsss(0)='1'  OR cVar1S1S23P024P047P066P007nsss(0)='1'  OR cVar2S2S23P016P018nsss(0)='1'  OR cVar2S3S23P016N018P006nsss(0)='1'  )then
          oVar1S204(0) <='1';
          else
          oVar1S204(0) <='0';
          end if;
        if(cVar2S4S23P002P061nsss(0)='1'  OR cVar2S5S23P002N061P059nsss(0)='1'  OR cVar2S6S23P002P012P018nsss(0)='1'  OR cVar2S7S23P011nsss(0)='1'  )then
          oVar1S205(0) <='1';
          else
          oVar1S205(0) <='0';
          end if;
        if(cVar2S8S23P020P040P021nsss(0)='1'  OR cVar2S9S23P020N040psss(0)='1'  OR cVar2S10S23P020P016P068nsss(0)='1'  OR cVar2S11S23P044P052nsss(0)='1'  )then
          oVar1S206(0) <='1';
          else
          oVar1S206(0) <='0';
          end if;
        if(cVar2S12S23P026nsss(0)='1'  OR cVar2S13S23N026P014nsss(0)='1'  OR cVar2S14S23N026N014P019nsss(0)='1'  OR cVar1S15S23N024N069P022P043nsss(0)='1'  )then
          oVar1S207(0) <='1';
          else
          oVar1S207(0) <='0';
          end if;
        if(cVar2S16S23P004nsss(0)='1'  OR cVar2S17S23N004P003P039nsss(0)='1'  OR cVar2S18S23P009P047P037nsss(0)='1'  OR cVar2S19S23P009P047P019nsss(0)='1'  )then
          oVar1S208(0) <='1';
          else
          oVar1S208(0) <='0';
          end if;
        if(cVar2S20S23P027P000P025nsss(0)='1'  OR cVar2S21S23N027P017P055nsss(0)='1'  OR cVar2S22S23N027N017P025nsss(0)='1'  )then
          oVar1S209(0) <='1';
          else
          oVar1S209(0) <='0';
          end if;
        if(cVar2S0S24P046nsss(0)='1'  OR cVar2S1S24P046P049nsss(0)='1'  OR cVar1S2S24P024P047P066P060psss(0)='1'  OR cVar1S3S24P024P047P066P069nsss(0)='1'  )then
          oVar1S210(0) <='1';
          else
          oVar1S210(0) <='0';
          end if;
        if(cVar2S4S24P016P018nsss(0)='1'  OR cVar2S5S24P016N018P019nsss(0)='1'  OR cVar2S6S24P045nsss(0)='1'  OR cVar2S7S24N045P037P068nsss(0)='1'  )then
          oVar1S211(0) <='1';
          else
          oVar1S211(0) <='0';
          end if;
        if(cVar2S8S24N045N037P019nsss(0)='1'  OR cVar2S9S24P059P015nsss(0)='1'  OR cVar2S10S24P059N015P032nsss(0)='1'  OR cVar2S11S24N059P006P068nsss(0)='1'  )then
          oVar1S212(0) <='1';
          else
          oVar1S212(0) <='0';
          end if;
        if(cVar1S12S24P024N047P010P025nsss(0)='1'  OR cVar2S13S24P018P011nsss(0)='1'  OR cVar1S14S24N024P040P021P035nsss(0)='1'  OR cVar2S15S24P062nsss(0)='1'  )then
          oVar1S213(0) <='1';
          else
          oVar1S213(0) <='0';
          end if;
        if(cVar2S16S24N062P012nsss(0)='1'  OR cVar2S17S24N062N012P019nsss(0)='1'  OR cVar2S18S24P023P018nsss(0)='1'  OR cVar2S19S24P023N018P004nsss(0)='1'  )then
          oVar1S214(0) <='1';
          else
          oVar1S214(0) <='0';
          end if;
        if(cVar2S20S24N023P002P038nsss(0)='1'  OR cVar2S21S24P020P005nsss(0)='1'  OR cVar2S22S24P020N005P041nsss(0)='1'  OR cVar2S23S24N020P041nsss(0)='1'  )then
          oVar1S215(0) <='1';
          else
          oVar1S215(0) <='0';
          end if;
        if(cVar2S24S24P021P026P049nsss(0)='1'  OR cVar2S25S24P021P019P036nsss(0)='1'  OR cVar2S26S24P019nsss(0)='1'  OR cVar2S27S24P048P013P046nsss(0)='1'  )then
          oVar1S216(0) <='1';
          else
          oVar1S216(0) <='0';
          end if;
        if(cVar2S28S24N048N069P020nsss(0)='1'  )then
          oVar1S217(0) <='1';
          else
          oVar1S217(0) <='0';
          end if;
        if(cVar2S0S25P017P056nsss(0)='1'  OR cVar2S1S25P017N056P060nsss(0)='1'  OR cVar2S2S25N017P018nsss(0)='1'  OR cVar2S3S25N017N018P008nsss(0)='1'  )then
          oVar1S218(0) <='1';
          else
          oVar1S218(0) <='0';
          end if;
        if(cVar2S4S25P018P064P063nsss(0)='1'  OR cVar2S5S25P062P059nsss(0)='1'  OR cVar2S6S25N062P005P030nsss(0)='1'  OR cVar2S7S25P054P014nsss(0)='1'  )then
          oVar1S219(0) <='1';
          else
          oVar1S219(0) <='0';
          end if;
        if(cVar2S8S25P054N014P034nsss(0)='1'  OR cVar2S9S25P055nsss(0)='1'  OR cVar2S10S25N055P014nsss(0)='1'  OR cVar2S11S25P059P013nsss(0)='1'  )then
          oVar1S220(0) <='1';
          else
          oVar1S220(0) <='0';
          end if;
        if(cVar2S12S25P059N013P064nsss(0)='1'  OR cVar2S13S25N059P013nsss(0)='1'  OR cVar2S14S25N059P013P069nsss(0)='1'  OR cVar2S15S25P015P068nsss(0)='1'  )then
          oVar1S221(0) <='1';
          else
          oVar1S221(0) <='0';
          end if;
        if(cVar2S16S25P015N068P035nsss(0)='1'  OR cVar2S17S25N015P049P063nsss(0)='1'  OR cVar2S18S25N015N049P047nsss(0)='1'  OR cVar2S19S25P028P051nsss(0)='1'  )then
          oVar1S222(0) <='1';
          else
          oVar1S222(0) <='0';
          end if;
        if(cVar2S20S25P028P051P010nsss(0)='1'  OR cVar2S21S25N028P032P061nsss(0)='1'  OR cVar2S22S25N028N032P029nsss(0)='1'  OR cVar2S23S25P036nsss(0)='1'  )then
          oVar1S223(0) <='1';
          else
          oVar1S223(0) <='0';
          end if;
        if(cVar2S24S25P016P019P017nsss(0)='1'  OR cVar2S25S25P016N019P068nsss(0)='1'  OR cVar1S26S25P001P023N067P041nsss(0)='1'  OR cVar2S27S25P029P019nsss(0)='1'  )then
          oVar1S224(0) <='1';
          else
          oVar1S224(0) <='0';
          end if;
        if(cVar2S28S25N029P037P013nsss(0)='1'  OR cVar2S29S25N029N037P030nsss(0)='1'  )then
          oVar1S225(0) <='1';
          else
          oVar1S225(0) <='0';
          end if;
        if(cVar2S0S26P028P051P000nsss(0)='1'  OR cVar2S1S26P069nsss(0)='1'  OR cVar2S2S26N069P063P013nsss(0)='1'  OR cVar2S3S26P047P045nsss(0)='1'  )then
          oVar1S226(0) <='1';
          else
          oVar1S226(0) <='0';
          end if;
        if(cVar2S4S26P065P035P013nsss(0)='1'  OR cVar2S5S26P065N035P036nsss(0)='1'  OR cVar2S6S26N065P067P019nsss(0)='1'  OR cVar2S7S26N065N067P057nsss(0)='1'  )then
          oVar1S227(0) <='1';
          else
          oVar1S227(0) <='0';
          end if;
        if(cVar2S8S26P002P065P016nsss(0)='1'  OR cVar2S9S26P002N065P033nsss(0)='1'  OR cVar2S10S26P002P012P011nsss(0)='1'  OR cVar2S11S26P034P036P018nsss(0)='1'  )then
          oVar1S228(0) <='1';
          else
          oVar1S228(0) <='0';
          end if;
        if(cVar2S12S26P037nsss(0)='1'  OR cVar2S13S26N037P035nsss(0)='1'  OR cVar2S14S26P024nsss(0)='1'  OR cVar2S15S26N024P025nsss(0)='1'  )then
          oVar1S229(0) <='1';
          else
          oVar1S229(0) <='0';
          end if;
        if(cVar2S16S26N024N025P031nsss(0)='1'  OR cVar2S17S26P016nsss(0)='1'  OR cVar2S18S26P016P014P019nsss(0)='1'  OR cVar2S19S26P018P069nsss(0)='1'  )then
          oVar1S230(0) <='1';
          else
          oVar1S230(0) <='0';
          end if;
        if(cVar2S20S26P018N069P056nsss(0)='1'  OR cVar2S21S26N018P010nsss(0)='1'  OR cVar2S22S26P057nsss(0)='1'  OR cVar2S23S26N057P056P018nsss(0)='1'  )then
          oVar1S231(0) <='1';
          else
          oVar1S231(0) <='0';
          end if;
        if(cVar2S24S26N057N056P058nsss(0)='1'  OR cVar2S25S26P064P054P057nsss(0)='1'  OR cVar2S26S26P064P054P037nsss(0)='1'  OR cVar2S27S26N064P010P067nsss(0)='1'  )then
          oVar1S232(0) <='1';
          else
          oVar1S232(0) <='0';
          end if;
        if(cVar2S28S26N064N010P027nsss(0)='1'  OR cVar2S29S26P013nsss(0)='1'  OR cVar2S30S26N013P014P012nsss(0)='1'  OR cVar2S31S26N013N014P011nsss(0)='1'  )then
          oVar1S233(0) <='1';
          else
          oVar1S233(0) <='0';
          end if;
        if(cVar2S32S26P063P055nsss(0)='1'  OR cVar2S33S26P063N055P036nsss(0)='1'  OR cVar2S34S26N063P060P017nsss(0)='1'  OR cVar2S35S26P047P027nsss(0)='1'  )then
          oVar1S234(0) <='1';
          else
          oVar1S234(0) <='0';
          end if;
        if(cVar2S36S26N047P046P025nsss(0)='1'  OR cVar2S37S26N047N046P022nsss(0)='1'  OR cVar2S38S26P023P042P066nsss(0)='1'  OR cVar2S39S26P023N042P064nsss(0)='1'  )then
          oVar1S235(0) <='1';
          else
          oVar1S235(0) <='0';
          end if;
        if(cVar2S40S26N023P053P068nsss(0)='1'  )then
          oVar1S236(0) <='1';
          else
          oVar1S236(0) <='0';
          end if;
        if(cVar1S0S27P002P022P043P007nsss(0)='1'  OR cVar2S1S27P003nsss(0)='1'  OR cVar2S2S27N003P005nsss(0)='1'  OR cVar2S3S27N003N005P004nsss(0)='1'  )then
          oVar1S237(0) <='1';
          else
          oVar1S237(0) <='0';
          end if;
        if(cVar2S4S27P018P004nsss(0)='1'  OR cVar2S5S27P018N004P006nsss(0)='1'  OR cVar2S6S27P003P039nsss(0)='1'  OR cVar2S7S27P003N039P057nsss(0)='1'  )then
          oVar1S238(0) <='1';
          else
          oVar1S238(0) <='0';
          end if;
        if(cVar2S8S27P017P006nsss(0)='1'  OR cVar2S9S27N017P008nsss(0)='1'  OR cVar2S10S27N017N008P006nsss(0)='1'  OR cVar2S11S27P010P069P015nsss(0)='1'  )then
          oVar1S239(0) <='1';
          else
          oVar1S239(0) <='0';
          end if;
        if(cVar2S12S27P035P060P033nsss(0)='1'  OR cVar2S13S27P035P060P033nsss(0)='1'  OR cVar2S14S27P035P016P060nsss(0)='1'  OR cVar2S15S27P059P061nsss(0)='1'  )then
          oVar1S240(0) <='1';
          else
          oVar1S240(0) <='0';
          end if;
        if(cVar2S16S27P059P061P013nsss(0)='1'  OR cVar2S17S27P059P061P064nsss(0)='1'  OR cVar2S18S27P059N061P013nsss(0)='1'  OR cVar1S19S27P002P040P021nsss(0)='1'  )then
          oVar1S241(0) <='1';
          else
          oVar1S241(0) <='0';
          end if;
        if(cVar1S20S27P002P040N021P038nsss(0)='1'  OR cVar2S21S27P019nsss(0)='1'  OR cVar2S22S27P053P019nsss(0)='1'  OR cVar2S23S27N053P069P010nsss(0)='1'  )then
          oVar1S242(0) <='1';
          else
          oVar1S242(0) <='0';
          end if;
        if(cVar2S0S28P036nsss(0)='1'  OR cVar2S1S28P036P069P063nsss(0)='1'  OR cVar2S2S28P059P058P069nsss(0)='1'  OR cVar2S3S28P059P058P012nsss(0)='1'  )then
          oVar1S244(0) <='1';
          else
          oVar1S244(0) <='0';
          end if;
        if(cVar2S4S28N059P058nsss(0)='1'  OR cVar2S5S28P034P010P059nsss(0)='1'  OR cVar2S6S28P034N010psss(0)='1'  OR cVar2S7S28P034P064nsss(0)='1'  )then
          oVar1S245(0) <='1';
          else
          oVar1S245(0) <='0';
          end if;
        if(cVar2S8S28P034N064P017nsss(0)='1'  OR cVar1S9S28P032P002P018P035nsss(0)='1'  OR cVar2S10S28P003nsss(0)='1'  OR cVar2S11S28P003P018P016nsss(0)='1'  )then
          oVar1S246(0) <='1';
          else
          oVar1S246(0) <='0';
          end if;
        if(cVar2S12S28P016P018nsss(0)='1'  OR cVar2S13S28P010P066nsss(0)='1'  OR cVar2S14S28P010N066P008nsss(0)='1'  OR cVar2S15S28P002P007P012nsss(0)='1'  )then
          oVar1S247(0) <='1';
          else
          oVar1S247(0) <='0';
          end if;
        if(cVar2S16S28P002N007psss(0)='1'  OR cVar2S17S28P002P043nsss(0)='1'  OR cVar2S18S28P035P068P015nsss(0)='1'  OR cVar2S19S28P031P057P056nsss(0)='1'  )then
          oVar1S248(0) <='1';
          else
          oVar1S248(0) <='0';
          end if;
        if(cVar2S20S28P031P019P037nsss(0)='1'  OR cVar2S21S28P031N019P065nsss(0)='1'  OR cVar2S22S28P039P020nsss(0)='1'  OR cVar2S23S28P039N020P005nsss(0)='1'  )then
          oVar1S249(0) <='1';
          else
          oVar1S249(0) <='0';
          end if;
        if(cVar2S24S28N039P025P046nsss(0)='1'  )then
          oVar1S250(0) <='1';
          else
          oVar1S250(0) <='0';
          end if;
        if(cVar1S0S29P040P021P035P002nsss(0)='1'  OR cVar2S1S29P004nsss(0)='1'  OR cVar2S2S29N004P019nsss(0)='1'  OR cVar2S3S29N004N019P038nsss(0)='1'  )then
          oVar1S251(0) <='1';
          else
          oVar1S251(0) <='0';
          end if;
        if(cVar2S4S29P062nsss(0)='1'  OR cVar2S5S29N062P012nsss(0)='1'  OR cVar2S6S29N062N012P068nsss(0)='1'  OR cVar2S7S29P036nsss(0)='1'  )then
          oVar1S252(0) <='1';
          else
          oVar1S252(0) <='0';
          end if;
        if(cVar2S8S29N036P015nsss(0)='1'  OR cVar2S9S29P046P035P000nsss(0)='1'  OR cVar2S10S29P063P062nsss(0)='1'  OR cVar2S11S29P063P062P015nsss(0)='1'  )then
          oVar1S253(0) <='1';
          else
          oVar1S253(0) <='0';
          end if;
        if(cVar2S12S29N063P064P019nsss(0)='1'  OR cVar2S13S29N063N064P068nsss(0)='1'  OR cVar2S14S29P050P016P000nsss(0)='1'  OR cVar2S15S29P050P016P003nsss(0)='1'  )then
          oVar1S254(0) <='1';
          else
          oVar1S254(0) <='0';
          end if;
        if(cVar2S16S29P050P013nsss(0)='1'  OR cVar2S17S29P051P012P011nsss(0)='1'  OR cVar2S18S29P014P003nsss(0)='1'  OR cVar1S19S29N040P038P026nsss(0)='1'  )then
          oVar1S255(0) <='1';
          else
          oVar1S255(0) <='0';
          end if;
        if(cVar2S20S29P015P036P062nsss(0)='1'  )then
          oVar1S256(0) <='1';
          else
          oVar1S256(0) <='0';
          end if;
        if(cVar2S0S30P009P048nsss(0)='1'  OR cVar2S1S30N009P062nsss(0)='1'  OR cVar2S2S30N009P062P007nsss(0)='1'  OR cVar2S3S30P006P026nsss(0)='1'  )then
          oVar1S257(0) <='1';
          else
          oVar1S257(0) <='0';
          end if;
        if(cVar2S4S30P006N026P016nsss(0)='1'  OR cVar2S5S30P045nsss(0)='1'  OR cVar2S6S30P009P018nsss(0)='1'  OR cVar2S7S30N009P048nsss(0)='1'  )then
          oVar1S258(0) <='1';
          else
          oVar1S258(0) <='0';
          end if;
        if(cVar2S8S30P029P051nsss(0)='1'  OR cVar2S9S30P029P051P011nsss(0)='1'  OR cVar2S10S30N029P028nsss(0)='1'  OR cVar2S11S30N029N028P026nsss(0)='1'  )then
          oVar1S259(0) <='1';
          else
          oVar1S259(0) <='0';
          end if;
        if(cVar2S12S30P036P015nsss(0)='1'  OR cVar2S13S30P035P017nsss(0)='1'  OR cVar2S14S30P035N017P063nsss(0)='1'  OR cVar2S15S30P035P065P017nsss(0)='1'  )then
          oVar1S260(0) <='1';
          else
          oVar1S260(0) <='0';
          end if;
        if(cVar2S16S30P053P049P066nsss(0)='1'  OR cVar2S17S30N053P057nsss(0)='1'  OR cVar2S18S30N053N057P011nsss(0)='1'  OR cVar2S19S30P065P067P066nsss(0)='1'  )then
          oVar1S261(0) <='1';
          else
          oVar1S261(0) <='0';
          end if;
        if(cVar2S20S30P065P067P037nsss(0)='1'  OR cVar2S21S30P065P036nsss(0)='1'  OR cVar2S22S30P065N036P062nsss(0)='1'  OR cVar2S23S30P024P049nsss(0)='1'  )then
          oVar1S262(0) <='1';
          else
          oVar1S262(0) <='0';
          end if;
        if(cVar2S24S30P024P049P006nsss(0)='1'  OR cVar2S25S30N024P009nsss(0)='1'  OR cVar2S26S30P064P028P013nsss(0)='1'  OR cVar2S27S30P064P028P011nsss(0)='1'  )then
          oVar1S263(0) <='1';
          else
          oVar1S263(0) <='0';
          end if;
        if(cVar2S28S30P037P029P017nsss(0)='1'  OR cVar2S29S30N037P061P035nsss(0)='1'  OR cVar2S30S30N037N061P041nsss(0)='1'  OR cVar2S31S30P053nsss(0)='1'  )then
          oVar1S264(0) <='1';
          else
          oVar1S264(0) <='0';
          end if;
        if(cVar2S32S30P069nsss(0)='1'  OR cVar2S33S30N069P011nsss(0)='1'  OR cVar2S34S30P010P019nsss(0)='1'  OR cVar2S35S30P010P019P056nsss(0)='1'  )then
          oVar1S265(0) <='1';
          else
          oVar1S265(0) <='0';
          end if;
        if(cVar2S36S30N010P017P011nsss(0)='1'  OR cVar2S37S30N010N017P003nsss(0)='1'  )then
          oVar1S266(0) <='1';
          else
          oVar1S266(0) <='0';
          end if;
        if(cVar2S0S31P019P017P034nsss(0)='1'  OR cVar2S1S31P019N017P034nsss(0)='1'  OR cVar2S2S31P019P059P066nsss(0)='1'  OR cVar2S3S31P019P059P069nsss(0)='1'  )then
          oVar1S267(0) <='1';
          else
          oVar1S267(0) <='0';
          end if;
        if(cVar2S4S31P066P019nsss(0)='1'  OR cVar2S5S31P066N019P017nsss(0)='1'  OR cVar1S6S31P036P063P005P035nsss(0)='1'  OR cVar2S7S31P067P017P015nsss(0)='1'  )then
          oVar1S268(0) <='1';
          else
          oVar1S268(0) <='0';
          end if;
        if(cVar2S8S31P017P018nsss(0)='1'  OR cVar2S9S31P017P018P014nsss(0)='1'  OR cVar2S10S31P017P015P008nsss(0)='1'  OR cVar2S11S31P017N015P014nsss(0)='1'  )then
          oVar1S269(0) <='1';
          else
          oVar1S269(0) <='0';
          end if;
        if(cVar2S12S31P062P035P069nsss(0)='1'  OR cVar2S13S31P062N035P013nsss(0)='1'  OR cVar2S14S31N062P055P067nsss(0)='1'  OR cVar2S15S31N062N055P056nsss(0)='1'  )then
          oVar1S270(0) <='1';
          else
          oVar1S270(0) <='0';
          end if;
        if(cVar2S16S31P034P015P066nsss(0)='1'  OR cVar2S17S31P034P015P021nsss(0)='1'  OR cVar2S18S31P034P068P037nsss(0)='1'  OR cVar2S19S31P034N068P012nsss(0)='1'  )then
          oVar1S271(0) <='1';
          else
          oVar1S271(0) <='0';
          end if;
        if(cVar2S20S31P067P060P033nsss(0)='1'  OR cVar2S21S31N067P058P033nsss(0)='1'  OR cVar2S22S31P051P066nsss(0)='1'  OR cVar2S23S31P051P066P019nsss(0)='1'  )then
          oVar1S272(0) <='1';
          else
          oVar1S272(0) <='0';
          end if;
        if(cVar2S24S31P051P019nsss(0)='1'  OR cVar2S25S31P051N019P064nsss(0)='1'  OR cVar2S26S31P046nsss(0)='1'  OR cVar2S27S31P056P069nsss(0)='1'  )then
          oVar1S273(0) <='1';
          else
          oVar1S273(0) <='0';
          end if;
        if(cVar2S28S31P056N069P029nsss(0)='1'  OR cVar2S29S31P067P049nsss(0)='1'  OR cVar2S30S31P067N049P058nsss(0)='1'  OR cVar2S31S31N067P066P055nsss(0)='1'  )then
          oVar1S274(0) <='1';
          else
          oVar1S274(0) <='0';
          end if;
        if(cVar2S32S31N067N066P064nsss(0)='1'  OR cVar2S33S31P037P005P066nsss(0)='1'  OR cVar2S34S31N037P059P032nsss(0)='1'  OR cVar2S35S31N037N059P045nsss(0)='1'  )then
          oVar1S275(0) <='1';
          else
          oVar1S275(0) <='0';
          end if;
        if(cVar2S36S31P015P047nsss(0)='1'  OR cVar2S37S31P015N047P013nsss(0)='1'  OR cVar2S38S31P015P016P064nsss(0)='1'  OR cVar2S39S31P015P016P011nsss(0)='1'  )then
          oVar1S276(0) <='1';
          else
          oVar1S276(0) <='0';
          end if;
        if(cVar2S40S31P016P068P037nsss(0)='1'  OR cVar2S41S31P016N068P035nsss(0)='1'  OR cVar2S42S31N016P048P042nsss(0)='1'  OR cVar2S43S31N016N048P042nsss(0)='1'  )then
          oVar1S277(0) <='1';
          else
          oVar1S277(0) <='0';
          end if;
        if(cVar2S0S32P023P019P048nsss(0)='1'  OR cVar2S1S32P023P019P064nsss(0)='1'  OR cVar2S2S32P009nsss(0)='1'  OR cVar2S3S32P018P012nsss(0)='1'  )then
          oVar1S279(0) <='1';
          else
          oVar1S279(0) <='0';
          end if;
        if(cVar2S4S32P034P047nsss(0)='1'  OR cVar2S5S32P034P059nsss(0)='1'  OR cVar2S6S32P034N059P019nsss(0)='1'  OR cVar2S7S32P003P013nsss(0)='1'  )then
          oVar1S280(0) <='1';
          else
          oVar1S280(0) <='0';
          end if;
        if(cVar2S8S32N003P008P012nsss(0)='1'  OR cVar2S9S32P017P062P037nsss(0)='1'  OR cVar2S10S32P017P062P014nsss(0)='1'  OR cVar2S11S32N017P018P050nsss(0)='1'  )then
          oVar1S281(0) <='1';
          else
          oVar1S281(0) <='0';
          end if;
        if(cVar2S12S32P019P069nsss(0)='1'  OR cVar2S13S32P033P064P004nsss(0)='1'  OR cVar2S14S32P033P064P059nsss(0)='1'  OR cVar2S15S32N033P054P012nsss(0)='1'  )then
          oVar1S282(0) <='1';
          else
          oVar1S282(0) <='0';
          end if;
        if(cVar2S16S32P035P032nsss(0)='1'  OR cVar2S17S32P035N032P065nsss(0)='1'  OR cVar2S18S32N035P017P037nsss(0)='1'  OR cVar2S19S32N035N017P068nsss(0)='1'  )then
          oVar1S283(0) <='1';
          else
          oVar1S283(0) <='0';
          end if;
        if(cVar1S20S32N036P060P048P006nsss(0)='1'  OR cVar2S21S32P009nsss(0)='1'  OR cVar2S22S32P019P067P057nsss(0)='1'  OR cVar2S23S32P019N067psss(0)='1'  )then
          oVar1S284(0) <='1';
          else
          oVar1S284(0) <='0';
          end if;
        if(cVar2S24S32P019P067P018nsss(0)='1'  OR cVar2S25S32P019P067P066nsss(0)='1'  OR cVar2S26S32P056P038P040nsss(0)='1'  OR cVar2S27S32P056N038P034nsss(0)='1'  )then
          oVar1S285(0) <='1';
          else
          oVar1S285(0) <='0';
          end if;
        if(cVar2S28S32P056P069P019nsss(0)='1'  OR cVar2S29S32P014P057nsss(0)='1'  OR cVar2S30S32N014P015P012nsss(0)='1'  OR cVar2S31S32N014N015P037nsss(0)='1'  )then
          oVar1S286(0) <='1';
          else
          oVar1S286(0) <='0';
          end if;
        if(cVar2S32S32P018P061P019nsss(0)='1'  )then
          oVar1S287(0) <='1';
          else
          oVar1S287(0) <='0';
          end if;
        if(cVar1S0S33P034P049P026P018nsss(0)='1'  OR cVar2S1S33P053P008P048nsss(0)='1'  OR cVar2S2S33P053P008P062nsss(0)='1'  OR cVar2S3S33P035P045P048nsss(0)='1'  )then
          oVar1S288(0) <='1';
          else
          oVar1S288(0) <='0';
          end if;
        if(cVar2S4S33P035P064nsss(0)='1'  OR cVar2S5S33P027P048nsss(0)='1'  OR cVar2S6S33N027P025P048nsss(0)='1'  OR cVar2S7S33N027N025P060nsss(0)='1'  )then
          oVar1S289(0) <='1';
          else
          oVar1S289(0) <='0';
          end if;
        if(cVar2S8S33P066nsss(0)='1'  OR cVar2S9S33P066P062P012nsss(0)='1'  OR cVar2S10S33P010P015nsss(0)='1'  OR cVar2S11S33P010N015P062nsss(0)='1'  )then
          oVar1S290(0) <='1';
          else
          oVar1S290(0) <='0';
          end if;
        if(cVar2S12S33N010P053P066nsss(0)='1'  OR cVar2S13S33N010N053P052nsss(0)='1'  OR cVar2S14S33P010P016P017nsss(0)='1'  OR cVar2S15S33P010N016P019nsss(0)='1'  )then
          oVar1S291(0) <='1';
          else
          oVar1S291(0) <='0';
          end if;
        if(cVar2S16S33P010P029nsss(0)='1'  OR cVar2S17S33P023P044nsss(0)='1'  OR cVar2S18S33P023N044P043nsss(0)='1'  OR cVar2S19S33N023P050nsss(0)='1'  )then
          oVar1S292(0) <='1';
          else
          oVar1S292(0) <='0';
          end if;
        if(cVar2S20S33N023N050P038nsss(0)='1'  OR cVar2S21S33P019P013nsss(0)='1'  OR cVar2S22S33P019P013P017nsss(0)='1'  OR cVar2S23S33N019P007P059nsss(0)='1'  )then
          oVar1S293(0) <='1';
          else
          oVar1S293(0) <='0';
          end if;
        if(cVar2S24S33P035P062P010nsss(0)='1'  OR cVar2S25S33P035N062P061nsss(0)='1'  OR cVar2S26S33P035P016P059nsss(0)='1'  OR cVar1S27S33P034N014P045P062nsss(0)='1'  )then
          oVar1S294(0) <='1';
          else
          oVar1S294(0) <='0';
          end if;
        if(cVar2S28S33P018P063nsss(0)='1'  OR cVar2S29S33P015P003P062nsss(0)='1'  OR cVar2S30S33N015P019P029nsss(0)='1'  OR cVar2S31S33P016P048nsss(0)='1'  )then
          oVar1S295(0) <='1';
          else
          oVar1S295(0) <='0';
          end if;
        if(cVar2S0S34P041P014nsss(0)='1'  OR cVar2S1S34N041P063P067nsss(0)='1'  OR cVar2S2S34N041N063psss(0)='1'  OR cVar2S3S34P010nsss(0)='1'  )then
          oVar1S297(0) <='1';
          else
          oVar1S297(0) <='0';
          end if;
        if(cVar2S4S34N010P058nsss(0)='1'  OR cVar2S5S34P061nsss(0)='1'  OR cVar2S6S34P061P013P065nsss(0)='1'  OR cVar2S7S34P013P035P011nsss(0)='1'  )then
          oVar1S298(0) <='1';
          else
          oVar1S298(0) <='0';
          end if;
        if(cVar2S8S34P013P035P033nsss(0)='1'  OR cVar2S9S34N013P015P052nsss(0)='1'  OR cVar2S10S34N013N015P030nsss(0)='1'  OR cVar2S11S34P066nsss(0)='1'  )then
          oVar1S299(0) <='1';
          else
          oVar1S299(0) <='0';
          end if;
        if(cVar2S12S34N066P015P006nsss(0)='1'  OR cVar2S13S34N066P015P007nsss(0)='1'  OR cVar2S14S34P017P058P035nsss(0)='1'  OR cVar2S15S34P017P058P060nsss(0)='1'  )then
          oVar1S300(0) <='1';
          else
          oVar1S300(0) <='0';
          end if;
        if(cVar2S16S34N017P015P014nsss(0)='1'  OR cVar2S17S34P016P060P011nsss(0)='1'  OR cVar2S18S34N016P012P063nsss(0)='1'  OR cVar2S19S34N016P012P010nsss(0)='1'  )then
          oVar1S301(0) <='1';
          else
          oVar1S301(0) <='0';
          end if;
        if(cVar2S20S34P066P069nsss(0)='1'  OR cVar2S21S34P066N069P016nsss(0)='1'  OR cVar2S22S34P066P011P013nsss(0)='1'  OR cVar2S23S34P066N011P055nsss(0)='1'  )then
          oVar1S302(0) <='1';
          else
          oVar1S302(0) <='0';
          end if;
        if(cVar2S24S34P035P012nsss(0)='1'  OR cVar2S25S34P035P012P019nsss(0)='1'  OR cVar2S26S34P035P019P016nsss(0)='1'  OR cVar2S27S34P014P037nsss(0)='1'  )then
          oVar1S303(0) <='1';
          else
          oVar1S303(0) <='0';
          end if;
        if(cVar2S28S34N014P069P061nsss(0)='1'  OR cVar2S29S34P059nsss(0)='1'  OR cVar2S30S34N059P037nsss(0)='1'  OR cVar2S31S34N059N037P058nsss(0)='1'  )then
          oVar1S304(0) <='1';
          else
          oVar1S304(0) <='0';
          end if;
        if(cVar2S32S34P036P015nsss(0)='1'  OR cVar2S33S34P036N015P019nsss(0)='1'  OR cVar2S34S34N036P019P035nsss(0)='1'  OR cVar2S35S34N036N019P016nsss(0)='1'  )then
          oVar1S305(0) <='1';
          else
          oVar1S305(0) <='0';
          end if;
        if(cVar2S36S34P066P060P017nsss(0)='1'  OR cVar2S37S34P066P060P011nsss(0)='1'  OR cVar2S38S34P066P017P018nsss(0)='1'  OR cVar2S39S34P061P068P015nsss(0)='1'  )then
          oVar1S306(0) <='1';
          else
          oVar1S306(0) <='0';
          end if;
        if(cVar2S40S34P061N068P016nsss(0)='1'  OR cVar2S41S34N061P060P058nsss(0)='1'  OR cVar2S42S34P016nsss(0)='1'  OR cVar2S43S34P050P065nsss(0)='1'  )then
          oVar1S307(0) <='1';
          else
          oVar1S307(0) <='0';
          end if;
        if(cVar2S44S34N050P056nsss(0)='1'  )then
          oVar1S308(0) <='1';
          else
          oVar1S308(0) <='0';
          end if;
        if(cVar1S0S35P061P064P030P013nsss(0)='1'  OR cVar2S1S35P016P057nsss(0)='1'  OR cVar2S2S35P016N057P015nsss(0)='1'  OR cVar2S3S35P033P058P032nsss(0)='1'  )then
          oVar1S309(0) <='1';
          else
          oVar1S309(0) <='0';
          end if;
        if(cVar2S4S35P033P058P063nsss(0)='1'  OR cVar2S5S35N033P056nsss(0)='1'  OR cVar2S6S35N033P056P012nsss(0)='1'  OR cVar2S7S35P037nsss(0)='1'  )then
          oVar1S310(0) <='1';
          else
          oVar1S310(0) <='0';
          end if;
        if(cVar1S8S35P061P064P058P008nsss(0)='1'  OR cVar2S9S35P018P034nsss(0)='1'  OR cVar2S10S35P018P034P014nsss(0)='1'  OR cVar2S11S35N018P068P033nsss(0)='1'  )then
          oVar1S311(0) <='1';
          else
          oVar1S311(0) <='0';
          end if;
        if(cVar2S12S35P035nsss(0)='1'  OR cVar2S13S35P056P052nsss(0)='1'  OR cVar2S14S35P056P052P012nsss(0)='1'  OR cVar2S15S35P056P054P069nsss(0)='1'  )then
          oVar1S312(0) <='1';
          else
          oVar1S312(0) <='0';
          end if;
        if(cVar2S16S35P064P016P018nsss(0)='1'  OR cVar2S17S35P017P019nsss(0)='1'  OR cVar2S18S35P033P055P029nsss(0)='1'  OR cVar2S19S35P033P055P011nsss(0)='1'  )then
          oVar1S313(0) <='1';
          else
          oVar1S313(0) <='0';
          end if;
        if(cVar2S20S35P033P017P019nsss(0)='1'  OR cVar2S21S35P033N017P016nsss(0)='1'  OR cVar2S22S35P018P015P011nsss(0)='1'  OR cVar2S23S35P018N015P063nsss(0)='1'  )then
          oVar1S314(0) <='1';
          else
          oVar1S314(0) <='0';
          end if;
        if(cVar2S24S35P035P036P065nsss(0)='1'  OR cVar2S25S35P035P036P019nsss(0)='1'  OR cVar2S26S35P049P009P048nsss(0)='1'  OR cVar2S27S35N049N067P060nsss(0)='1'  )then
          oVar1S315(0) <='1';
          else
          oVar1S315(0) <='0';
          end if;
        if(cVar2S0S36P035P019nsss(0)='1'  OR cVar2S1S36P035P019P036nsss(0)='1'  OR cVar2S2S36N035P025P058nsss(0)='1'  OR cVar2S3S36N035P025P034nsss(0)='1'  )then
          oVar1S317(0) <='1';
          else
          oVar1S317(0) <='0';
          end if;
        if(cVar2S4S36P052P059nsss(0)='1'  OR cVar2S5S36P017P061nsss(0)='1'  OR cVar2S6S36P017N061P060nsss(0)='1'  OR cVar2S7S36N017P019P015nsss(0)='1'  )then
          oVar1S318(0) <='1';
          else
          oVar1S318(0) <='0';
          end if;
        if(cVar2S8S36P034P009nsss(0)='1'  OR cVar2S9S36P012P060nsss(0)='1'  OR cVar2S10S36P012N060P055nsss(0)='1'  OR cVar2S11S36N012P040nsss(0)='1'  )then
          oVar1S319(0) <='1';
          else
          oVar1S319(0) <='0';
          end if;
        if(cVar2S12S36N012N040P047nsss(0)='1'  OR cVar2S13S36P066nsss(0)='1'  OR cVar2S14S36P035nsss(0)='1'  OR cVar2S15S36P058P066P054nsss(0)='1'  )then
          oVar1S320(0) <='1';
          else
          oVar1S320(0) <='0';
          end if;
        if(cVar2S16S36P058P066P053nsss(0)='1'  OR cVar2S17S36P058P018nsss(0)='1'  OR cVar2S18S36P058P018P013nsss(0)='1'  OR cVar2S19S36P062P018P068nsss(0)='1'  )then
          oVar1S321(0) <='1';
          else
          oVar1S321(0) <='0';
          end if;
        if(cVar2S20S36P062N018P068nsss(0)='1'  OR cVar2S21S36P062P060P066nsss(0)='1'  OR cVar2S22S36P035P034P068nsss(0)='1'  OR cVar2S23S36P035P019P017nsss(0)='1'  )then
          oVar1S322(0) <='1';
          else
          oVar1S322(0) <='0';
          end if;
        if(cVar2S24S36P014P010P018nsss(0)='1'  OR cVar2S25S36N014P016P019nsss(0)='1'  OR cVar2S26S36P052P026nsss(0)='1'  OR cVar2S27S36P052N026P060nsss(0)='1'  )then
          oVar1S323(0) <='1';
          else
          oVar1S323(0) <='0';
          end if;
        if(cVar2S28S36P052P018nsss(0)='1'  OR cVar2S29S36P026P019P018nsss(0)='1'  OR cVar2S30S36P043nsss(0)='1'  OR cVar2S31S36N043P035P026nsss(0)='1'  )then
          oVar1S324(0) <='1';
          else
          oVar1S324(0) <='0';
          end if;
        if(cVar2S32S36P068P066P039nsss(0)='1'  OR cVar2S33S36N068P069P047nsss(0)='1'  )then
          oVar1S325(0) <='1';
          else
          oVar1S325(0) <='0';
          end if;
        if(cVar2S0S37P066P036P018nsss(0)='1'  OR cVar2S1S37P066N036P015nsss(0)='1'  OR cVar2S2S37N066P064nsss(0)='1'  OR cVar2S3S37P011P016P036nsss(0)='1'  )then
          oVar1S326(0) <='1';
          else
          oVar1S326(0) <='0';
          end if;
        if(cVar2S4S37N011P062P049nsss(0)='1'  OR cVar2S5S37N011N062P059nsss(0)='1'  OR cVar2S6S37P044P041nsss(0)='1'  OR cVar2S7S37P052P060P068nsss(0)='1'  )then
          oVar1S327(0) <='1';
          else
          oVar1S327(0) <='0';
          end if;
        if(cVar2S8S37P014P034P019nsss(0)='1'  OR cVar2S9S37P014P034P011nsss(0)='1'  OR cVar2S10S37P014P047nsss(0)='1'  OR cVar2S11S37P014N047P055nsss(0)='1'  )then
          oVar1S328(0) <='1';
          else
          oVar1S328(0) <='0';
          end if;
        if(cVar2S12S37P058P014nsss(0)='1'  OR cVar2S13S37P058N014P019nsss(0)='1'  OR cVar2S14S37P058P015nsss(0)='1'  OR cVar2S15S37P019P010P064nsss(0)='1'  )then
          oVar1S329(0) <='1';
          else
          oVar1S329(0) <='0';
          end if;
        if(cVar2S16S37P019P010P066nsss(0)='1'  OR cVar2S17S37P063nsss(0)='1'  OR cVar2S18S37P012P033nsss(0)='1'  OR cVar2S19S37P012P033P016nsss(0)='1'  )then
          oVar1S330(0) <='1';
          else
          oVar1S330(0) <='0';
          end if;
        if(cVar2S20S37N012P014P036nsss(0)='1'  OR cVar2S21S37N012N014P019nsss(0)='1'  OR cVar2S22S37P015nsss(0)='1'  OR cVar2S23S37P066P069P068nsss(0)='1'  )then
          oVar1S331(0) <='1';
          else
          oVar1S331(0) <='0';
          end if;
        if(cVar2S24S37P066P036P052nsss(0)='1'  OR cVar2S25S37P066N036P069nsss(0)='1'  OR cVar2S26S37P018P057nsss(0)='1'  OR cVar2S27S37P018N057P015nsss(0)='1'  )then
          oVar1S332(0) <='1';
          else
          oVar1S332(0) <='0';
          end if;
        if(cVar2S28S37N018P000nsss(0)='1'  OR cVar2S29S37P017P018nsss(0)='1'  OR cVar2S30S37P017N018P037nsss(0)='1'  OR cVar2S31S37N017P068nsss(0)='1'  )then
          oVar1S333(0) <='1';
          else
          oVar1S333(0) <='0';
          end if;
        if(cVar2S32S37N017N068P018nsss(0)='1'  OR cVar2S33S37P058P045nsss(0)='1'  )then
          oVar1S334(0) <='1';
          else
          oVar1S334(0) <='0';
          end if;
        if(cVar2S0S38P024P029P054nsss(0)='1'  OR cVar2S1S38P024P029P016nsss(0)='1'  OR cVar2S2S38P062nsss(0)='1'  OR cVar2S3S38N062P008nsss(0)='1'  )then
          oVar1S335(0) <='1';
          else
          oVar1S335(0) <='0';
          end if;
        if(cVar2S4S38P064nsss(0)='1'  OR cVar2S5S38N064P003P063nsss(0)='1'  OR cVar2S6S38P062P058nsss(0)='1'  OR cVar2S7S38P062P058P018nsss(0)='1'  )then
          oVar1S336(0) <='1';
          else
          oVar1S336(0) <='0';
          end if;
        if(cVar2S8S38P062P067nsss(0)='1'  OR cVar2S9S38P062P067P060nsss(0)='1'  OR cVar2S10S38P011P010P028nsss(0)='1'  OR cVar2S11S38P011P010P017nsss(0)='1'  )then
          oVar1S337(0) <='1';
          else
          oVar1S337(0) <='0';
          end if;
        if(cVar2S12S38P011P027nsss(0)='1'  OR cVar2S13S38P011N027P037nsss(0)='1'  OR cVar2S14S38P007P011P018nsss(0)='1'  OR cVar2S15S38P061P015P053nsss(0)='1'  )then
          oVar1S338(0) <='1';
          else
          oVar1S338(0) <='0';
          end if;
        if(cVar2S16S38P061P015P023nsss(0)='1'  OR cVar2S17S38P061P017P034nsss(0)='1'  OR cVar2S18S38P015P061P032nsss(0)='1'  OR cVar2S19S38P015N061P018nsss(0)='1'  )then
          oVar1S339(0) <='1';
          else
          oVar1S339(0) <='0';
          end if;
        if(cVar2S20S38N015P012P017nsss(0)='1'  OR cVar2S21S38P056P057P016nsss(0)='1'  OR cVar2S22S38P056P057P031nsss(0)='1'  OR cVar2S23S38N056P018nsss(0)='1'  )then
          oVar1S340(0) <='1';
          else
          oVar1S340(0) <='0';
          end if;
        if(cVar2S24S38N056N018P032nsss(0)='1'  OR cVar2S25S38P066P007P017nsss(0)='1'  OR cVar2S26S38P020P005nsss(0)='1'  OR cVar2S27S38P020N005P040nsss(0)='1'  )then
          oVar1S341(0) <='1';
          else
          oVar1S341(0) <='0';
          end if;
        if(cVar2S28S38N020P013P062nsss(0)='1'  OR cVar2S29S38P011P060P028nsss(0)='1'  OR cVar2S30S38P011N060psss(0)='1'  OR cVar2S31S38N011P024P026nsss(0)='1'  )then
          oVar1S342(0) <='1';
          else
          oVar1S342(0) <='0';
          end if;
        if(cVar2S32S38P064P015nsss(0)='1'  OR cVar2S33S38P064P015P059nsss(0)='1'  OR cVar2S34S38P064P065nsss(0)='1'  OR cVar2S35S38P054P036nsss(0)='1'  )then
          oVar1S343(0) <='1';
          else
          oVar1S343(0) <='0';
          end if;
        if(cVar2S36S38P054P036P018nsss(0)='1'  OR cVar2S37S38P065P063P017nsss(0)='1'  OR cVar2S38S38N065P035P010nsss(0)='1'  )then
          oVar1S344(0) <='1';
          else
          oVar1S344(0) <='0';
          end if;
        if(cVar2S0S39P019P059P009nsss(0)='1'  OR cVar2S1S39P019N059P033nsss(0)='1'  OR cVar2S2S39P019P068P032nsss(0)='1'  OR cVar2S3S39P019N068P065nsss(0)='1'  )then
          oVar1S345(0) <='1';
          else
          oVar1S345(0) <='0';
          end if;
        if(cVar2S4S39P068P065P037nsss(0)='1'  OR cVar2S5S39P068P065P036nsss(0)='1'  OR cVar2S6S39N068P047nsss(0)='1'  OR cVar2S7S39N068N047P045nsss(0)='1'  )then
          oVar1S346(0) <='1';
          else
          oVar1S346(0) <='0';
          end if;
        if(cVar2S8S39P056P057nsss(0)='1'  OR cVar2S9S39P056P057P014nsss(0)='1'  OR cVar2S10S39N056P054P060nsss(0)='1'  OR cVar2S11S39P015P035P034nsss(0)='1'  )then
          oVar1S347(0) <='1';
          else
          oVar1S347(0) <='0';
          end if;
        if(cVar2S12S39P015N035P016nsss(0)='1'  OR cVar2S13S39P037P018P033nsss(0)='1'  OR cVar2S14S39P037N018P014nsss(0)='1'  OR cVar2S15S39P037P036P018nsss(0)='1'  )then
          oVar1S348(0) <='1';
          else
          oVar1S348(0) <='0';
          end if;
        if(cVar2S16S39P037P036P012nsss(0)='1'  OR cVar2S17S39P046P018nsss(0)='1'  OR cVar2S18S39N046P015P033nsss(0)='1'  OR cVar2S19S39P063nsss(0)='1'  )then
          oVar1S349(0) <='1';
          else
          oVar1S349(0) <='0';
          end if;
        if(cVar2S20S39P067P001nsss(0)='1'  OR cVar2S21S39N067P019P066nsss(0)='1'  OR cVar2S22S39P057nsss(0)='1'  OR cVar2S23S39N057P036nsss(0)='1'  )then
          oVar1S350(0) <='1';
          else
          oVar1S350(0) <='0';
          end if;
        if(cVar2S24S39N057N036P017nsss(0)='1'  OR cVar2S25S39P009P069nsss(0)='1'  OR cVar2S26S39P009N069P037nsss(0)='1'  OR cVar2S27S39P009P018P066nsss(0)='1'  )then
          oVar1S351(0) <='1';
          else
          oVar1S351(0) <='0';
          end if;
        if(cVar2S28S39P037P069nsss(0)='1'  OR cVar2S29S39P037N069P055nsss(0)='1'  OR cVar2S30S39N037P061P014nsss(0)='1'  OR cVar2S31S39P014P015P037nsss(0)='1'  )then
          oVar1S352(0) <='1';
          else
          oVar1S352(0) <='0';
          end if;
        if(cVar2S32S39P034nsss(0)='1'  OR cVar2S33S39N034P018nsss(0)='1'  OR cVar2S34S39N034N018P032nsss(0)='1'  OR cVar2S35S39P026P057nsss(0)='1'  )then
          oVar1S353(0) <='1';
          else
          oVar1S353(0) <='0';
          end if;
        if(cVar2S36S39P026N057P063nsss(0)='1'  OR cVar2S37S39P026nsss(0)='1'  OR cVar2S38S39N026P066nsss(0)='1'  OR cVar2S39S39P067P054P032nsss(0)='1'  )then
          oVar1S354(0) <='1';
          else
          oVar1S354(0) <='0';
          end if;
        if(cVar2S40S39P067P055P018nsss(0)='1'  )then
          oVar1S355(0) <='1';
          else
          oVar1S355(0) <='0';
          end if;
        if(cVar2S0S40P058nsss(0)='1'  OR cVar2S1S40P058P012P065nsss(0)='1'  OR cVar2S2S40P058N012P063nsss(0)='1'  OR cVar2S3S40P019P047nsss(0)='1'  )then
          oVar1S356(0) <='1';
          else
          oVar1S356(0) <='0';
          end if;
        if(cVar2S4S40N019P063nsss(0)='1'  OR cVar2S5S40P068P063nsss(0)='1'  OR cVar2S6S40P068N063P013nsss(0)='1'  OR cVar2S7S40P068P037nsss(0)='1'  )then
          oVar1S357(0) <='1';
          else
          oVar1S357(0) <='0';
          end if;
        if(cVar2S8S40P068P017nsss(0)='1'  OR cVar2S9S40P068N017P019nsss(0)='1'  OR cVar2S10S40N068P060P065nsss(0)='1'  OR cVar2S11S40N068N060P052nsss(0)='1'  )then
          oVar1S358(0) <='1';
          else
          oVar1S358(0) <='0';
          end if;
        if(cVar1S12S40P069P053P059P060nsss(0)='1'  OR cVar2S13S40P057P006P054nsss(0)='1'  OR cVar2S14S40P030P059nsss(0)='1'  OR cVar2S15S40P030P059P012nsss(0)='1'  )then
          oVar1S359(0) <='1';
          else
          oVar1S359(0) <='0';
          end if;
        if(cVar2S16S40P030P011P010nsss(0)='1'  OR cVar2S17S40P011nsss(0)='1'  OR cVar2S18S40N011P056P057nsss(0)='1'  OR cVar2S19S40N011P056P018nsss(0)='1'  )then
          oVar1S360(0) <='1';
          else
          oVar1S360(0) <='0';
          end if;
        if(cVar2S20S40P033nsss(0)='1'  OR cVar2S21S40P033P054nsss(0)='1'  OR cVar2S22S40P054P035nsss(0)='1'  OR cVar2S23S40N054P011P014nsss(0)='1'  )then
          oVar1S361(0) <='1';
          else
          oVar1S361(0) <='0';
          end if;
        if(cVar2S24S40N054N011P029nsss(0)='1'  OR cVar2S25S40P013nsss(0)='1'  OR cVar2S26S40N013P062nsss(0)='1'  OR cVar2S27S40P045nsss(0)='1'  )then
          oVar1S362(0) <='1';
          else
          oVar1S362(0) <='0';
          end if;
        if(cVar2S28S40N045P064P013nsss(0)='1'  OR cVar2S29S40N045P064P037nsss(0)='1'  OR cVar2S30S40P058P013P026nsss(0)='1'  OR cVar2S31S40P058P013P059nsss(0)='1'  )then
          oVar1S363(0) <='1';
          else
          oVar1S363(0) <='0';
          end if;
        if(cVar2S32S40P058P014P016nsss(0)='1'  OR cVar2S33S40P062P035nsss(0)='1'  OR cVar2S34S40P062N035P033nsss(0)='1'  OR cVar2S35S40N062P059P015nsss(0)='1'  )then
          oVar1S364(0) <='1';
          else
          oVar1S364(0) <='0';
          end if;
        if(cVar2S36S40N062N059P020nsss(0)='1'  )then
          oVar1S365(0) <='1';
          else
          oVar1S365(0) <='0';
          end if;
        if(cVar1S0S41P025P004P048nsss(0)='1'  OR cVar1S1S41P025P004N048P008nsss(0)='1'  OR cVar2S2S41P065P003nsss(0)='1'  OR cVar2S3S41P065P016nsss(0)='1'  )then
          oVar1S366(0) <='1';
          else
          oVar1S366(0) <='0';
          end if;
        if(cVar2S4S41P044P036nsss(0)='1'  OR cVar2S5S41P015P016nsss(0)='1'  OR cVar2S6S41N015P017nsss(0)='1'  OR cVar2S7S41P033P012nsss(0)='1'  )then
          oVar1S367(0) <='1';
          else
          oVar1S367(0) <='0';
          end if;
        if(cVar2S8S41N033P006nsss(0)='1'  OR cVar2S9S41N033N006P009nsss(0)='1'  OR cVar2S10S41P067P006nsss(0)='1'  OR cVar2S11S41P067P006P056nsss(0)='1'  )then
          oVar1S368(0) <='1';
          else
          oVar1S368(0) <='0';
          end if;
        if(cVar2S12S41P067P046P018nsss(0)='1'  OR cVar2S13S41P013P031P054nsss(0)='1'  OR cVar2S14S41P013N031P018nsss(0)='1'  OR cVar2S15S41N013P068nsss(0)='1'  )then
          oVar1S369(0) <='1';
          else
          oVar1S369(0) <='0';
          end if;
        if(cVar2S16S41N013N068P056nsss(0)='1'  OR cVar2S17S41P048P063P059nsss(0)='1'  OR cVar2S18S41P048N063P035nsss(0)='1'  OR cVar2S19S41P046P008nsss(0)='1'  )then
          oVar1S370(0) <='1';
          else
          oVar1S370(0) <='0';
          end if;
        if(cVar2S20S41P046N008P036nsss(0)='1'  OR cVar2S21S41N046P069nsss(0)='1'  OR cVar2S22S41N046P069P048nsss(0)='1'  OR cVar2S23S41P009nsss(0)='1'  )then
          oVar1S371(0) <='1';
          else
          oVar1S371(0) <='0';
          end if;
        if(cVar2S24S41P056P033P008nsss(0)='1'  OR cVar2S25S41P056N033P054nsss(0)='1'  OR cVar2S26S41N056P068P064nsss(0)='1'  OR cVar2S27S41N056N068P055nsss(0)='1'  )then
          oVar1S372(0) <='1';
          else
          oVar1S372(0) <='0';
          end if;
        if(cVar2S28S41P069P010nsss(0)='1'  OR cVar2S29S41P069N010P024nsss(0)='1'  )then
          oVar1S373(0) <='1';
          else
          oVar1S373(0) <='0';
          end if;
        if(cVar1S0S42P068P004P025P048nsss(0)='1'  OR cVar2S1S42P012nsss(0)='1'  OR cVar2S2S42P021nsss(0)='1'  OR cVar2S3S42N021P020nsss(0)='1'  )then
          oVar1S374(0) <='1';
          else
          oVar1S374(0) <='0';
          end if;
        if(cVar2S4S42N021N020P023nsss(0)='1'  OR cVar2S5S42P044nsss(0)='1'  OR cVar2S6S42N044P048P022nsss(0)='1'  OR cVar2S7S42P057nsss(0)='1'  )then
          oVar1S375(0) <='1';
          else
          oVar1S375(0) <='0';
          end if;
        if(cVar2S8S42P057P035P059nsss(0)='1'  OR cVar2S9S42P058P005nsss(0)='1'  OR cVar2S10S42N058P052P010nsss(0)='1'  OR cVar2S11S42N058N052P030nsss(0)='1'  )then
          oVar1S376(0) <='1';
          else
          oVar1S376(0) <='0';
          end if;
        if(cVar2S12S42P057P019P036nsss(0)='1'  OR cVar2S13S42P057N019P064nsss(0)='1'  OR cVar2S14S42N057P069P061nsss(0)='1'  OR cVar2S15S42N057N069P014nsss(0)='1'  )then
          oVar1S377(0) <='1';
          else
          oVar1S377(0) <='0';
          end if;
        if(cVar2S16S42P065nsss(0)='1'  OR cVar2S17S42P032P007nsss(0)='1'  OR cVar2S18S42P032P037nsss(0)='1'  OR cVar2S19S42P032P037P014nsss(0)='1'  )then
          oVar1S378(0) <='1';
          else
          oVar1S378(0) <='0';
          end if;
        if(cVar2S20S42P014nsss(0)='1'  OR cVar2S21S42N014P013nsss(0)='1'  OR cVar1S22S42P068P015N061P025nsss(0)='1'  OR cVar2S23S42P016P037P001nsss(0)='1'  )then
          oVar1S379(0) <='1';
          else
          oVar1S379(0) <='0';
          end if;
        if(cVar2S24S42P016N037P036nsss(0)='1'  OR cVar2S25S42N016P066P052nsss(0)='1'  OR cVar2S26S42P033P063P036nsss(0)='1'  OR cVar2S27S42P033P034nsss(0)='1'  )then
          oVar1S380(0) <='1';
          else
          oVar1S380(0) <='0';
          end if;
        if(cVar2S28S42P019P063P008nsss(0)='1'  OR cVar2S29S42P019P009nsss(0)='1'  OR cVar2S30S42P019N009P033nsss(0)='1'  OR cVar2S31S42P060P057nsss(0)='1'  )then
          oVar1S381(0) <='1';
          else
          oVar1S381(0) <='0';
          end if;
        if(cVar2S32S42P060N057P016nsss(0)='1'  OR cVar2S33S42P060P017nsss(0)='1'  OR cVar2S34S42P060N017P012nsss(0)='1'  OR cVar2S35S42P062P036P064nsss(0)='1'  )then
          oVar1S382(0) <='1';
          else
          oVar1S382(0) <='0';
          end if;
        if(cVar2S36S42N062P069P014nsss(0)='1'  )then
          oVar1S383(0) <='1';
          else
          oVar1S383(0) <='0';
          end if;
        if(cVar2S0S43P043P019P013nsss(0)='1'  OR cVar2S1S43P043P019P004nsss(0)='1'  OR cVar2S2S43N043P024nsss(0)='1'  OR cVar2S3S43N043P024P056nsss(0)='1'  )then
          oVar1S384(0) <='1';
          else
          oVar1S384(0) <='0';
          end if;
        if(cVar2S4S43P024P049nsss(0)='1'  OR cVar2S5S43P024P049P006nsss(0)='1'  OR cVar2S6S43N024P064P013nsss(0)='1'  OR cVar2S7S43P037nsss(0)='1'  )then
          oVar1S385(0) <='1';
          else
          oVar1S385(0) <='0';
          end if;
        if(cVar2S8S43P018P012nsss(0)='1'  OR cVar2S9S43N018P017P010nsss(0)='1'  OR cVar2S10S43P022P015P029nsss(0)='1'  OR cVar2S11S43P022P015P009nsss(0)='1'  )then
          oVar1S386(0) <='1';
          else
          oVar1S386(0) <='0';
          end if;
        if(cVar2S12S43P064P017nsss(0)='1'  OR cVar2S13S43P064P017P016nsss(0)='1'  OR cVar2S14S43N064P066P012nsss(0)='1'  OR cVar1S15S43N068P004P025P048nsss(0)='1'  )then
          oVar1S387(0) <='1';
          else
          oVar1S387(0) <='0';
          end if;
        if(cVar2S16S43P012nsss(0)='1'  OR cVar2S17S43P019nsss(0)='1'  OR cVar2S18S43N019P021nsss(0)='1'  OR cVar2S19S43N019N021P020nsss(0)='1'  )then
          oVar1S388(0) <='1';
          else
          oVar1S388(0) <='0';
          end if;
        if(cVar2S20S43P042P017nsss(0)='1'  OR cVar2S21S43P042N017P036nsss(0)='1'  OR cVar2S22S43N042P021P018nsss(0)='1'  OR cVar2S23S43P023P057nsss(0)='1'  )then
          oVar1S389(0) <='1';
          else
          oVar1S389(0) <='0';
          end if;
        if(cVar2S24S43P023N057P036nsss(0)='1'  OR cVar2S25S43P066P052P065nsss(0)='1'  OR cVar2S26S43P066N052P058nsss(0)='1'  OR cVar2S27S43P066P067P015nsss(0)='1'  )then
          oVar1S390(0) <='1';
          else
          oVar1S390(0) <='0';
          end if;
        if(cVar2S28S43P052P035P017nsss(0)='1'  OR cVar2S29S43P052P035P016nsss(0)='1'  OR cVar2S30S43P052P010nsss(0)='1'  OR cVar2S31S43P052N010P059nsss(0)='1'  )then
          oVar1S391(0) <='1';
          else
          oVar1S391(0) <='0';
          end if;
        if(cVar2S32S43P024P007nsss(0)='1'  OR cVar2S33S43P024N007P006nsss(0)='1'  )then
          oVar1S392(0) <='1';
          else
          oVar1S392(0) <='0';
          end if;
        if(cVar2S0S44P026P029P060nsss(0)='1'  OR cVar2S1S44P054P035P069nsss(0)='1'  OR cVar2S2S44P054P035P049nsss(0)='1'  OR cVar2S3S44P054P012P037nsss(0)='1'  )then
          oVar1S393(0) <='1';
          else
          oVar1S393(0) <='0';
          end if;
        if(cVar2S4S44P054N012P010nsss(0)='1'  OR cVar2S5S44P042P047P065nsss(0)='1'  OR cVar2S6S44P042P047P017nsss(0)='1'  OR cVar2S7S44P038P002nsss(0)='1'  )then
          oVar1S394(0) <='1';
          else
          oVar1S394(0) <='0';
          end if;
        if(cVar2S8S44P038N002P004nsss(0)='1'  OR cVar2S9S44N038P044nsss(0)='1'  OR cVar2S10S44N038N044P014nsss(0)='1'  OR cVar2S11S44P033P014P015nsss(0)='1'  )then
          oVar1S395(0) <='1';
          else
          oVar1S395(0) <='0';
          end if;
        if(cVar2S12S44P033N014P040nsss(0)='1'  OR cVar2S13S44P033P009P017nsss(0)='1'  OR cVar2S14S44P067P018nsss(0)='1'  OR cVar2S15S44P038nsss(0)='1'  )then
          oVar1S396(0) <='1';
          else
          oVar1S396(0) <='0';
          end if;
        if(cVar1S16S44P068P067P057P032nsss(0)='1'  OR cVar2S17S44P035nsss(0)='1'  OR cVar2S18S44N035P037P030nsss(0)='1'  OR cVar2S19S44P037nsss(0)='1'  )then
          oVar1S397(0) <='1';
          else
          oVar1S397(0) <='0';
          end if;
        if(cVar2S20S44N037P017nsss(0)='1'  OR cVar2S21S44N037N017P013nsss(0)='1'  OR cVar2S22S44P015P018nsss(0)='1'  OR cVar2S23S44P015P059P032nsss(0)='1'  )then
          oVar1S398(0) <='1';
          else
          oVar1S398(0) <='0';
          end if;
        if(cVar2S24S44P003P012P016nsss(0)='1'  OR cVar2S25S44P003P012P014nsss(0)='1'  )then
          oVar1S399(0) <='1';
          else
          oVar1S399(0) <='0';
          end if;
        if(cVar2S0S45P062P066P064nsss(0)='1'  OR cVar2S1S45P062N066P064nsss(0)='1'  OR cVar2S2S45P062psss(0)='1'  OR cVar2S3S45P024nsss(0)='1'  )then
          oVar1S400(0) <='1';
          else
          oVar1S400(0) <='0';
          end if;
        if(cVar2S4S45N024P066P042nsss(0)='1'  OR cVar2S5S45P019P034P054nsss(0)='1'  OR cVar2S6S45P019P034P060nsss(0)='1'  OR cVar2S7S45N019P029P059nsss(0)='1'  )then
          oVar1S401(0) <='1';
          else
          oVar1S401(0) <='0';
          end if;
        if(cVar2S8S45N019N029P012nsss(0)='1'  OR cVar2S9S45P017P045P060nsss(0)='1'  OR cVar2S10S45N017P019P034nsss(0)='1'  OR cVar2S11S45N017N019P060nsss(0)='1'  )then
          oVar1S402(0) <='1';
          else
          oVar1S402(0) <='0';
          end if;
        if(cVar2S12S45P008nsss(0)='1'  OR cVar2S13S45N008P036nsss(0)='1'  OR cVar2S14S45P027P065nsss(0)='1'  OR cVar2S15S45N027P009P010nsss(0)='1'  )then
          oVar1S403(0) <='1';
          else
          oVar1S403(0) <='0';
          end if;
        if(cVar2S16S45N027P009P004nsss(0)='1'  OR cVar2S17S45P062nsss(0)='1'  OR cVar2S18S45N062P015P016nsss(0)='1'  OR cVar2S19S45P008nsss(0)='1'  )then
          oVar1S404(0) <='1';
          else
          oVar1S404(0) <='0';
          end if;
        if(cVar2S20S45P008P065P035nsss(0)='1'  OR cVar2S21S45P010P060nsss(0)='1'  OR cVar2S22S45P010N060P029nsss(0)='1'  OR cVar2S23S45N010P005P053nsss(0)='1'  )then
          oVar1S405(0) <='1';
          else
          oVar1S405(0) <='0';
          end if;
        if(cVar2S24S45P017nsss(0)='1'  OR cVar2S25S45P010P012P032nsss(0)='1'  OR cVar2S26S45P066nsss(0)='1'  OR cVar2S27S45N066P016P034nsss(0)='1'  )then
          oVar1S406(0) <='1';
          else
          oVar1S406(0) <='0';
          end if;
        if(cVar2S28S45P065P059P013nsss(0)='1'  OR cVar2S29S45N065P046P062nsss(0)='1'  OR cVar2S30S45P053nsss(0)='1'  )then
          oVar1S407(0) <='1';
          else
          oVar1S407(0) <='0';
          end if;
        if(cVar1S0S46P016P038P021nsss(0)='1'  OR cVar2S1S46P058nsss(0)='1'  OR cVar2S2S46N058P007nsss(0)='1'  OR cVar2S3S46N058N007P065nsss(0)='1'  )then
          oVar1S408(0) <='1';
          else
          oVar1S408(0) <='0';
          end if;
        if(cVar2S4S46N069N037P014nsss(0)='1'  OR cVar2S5S46P034P011nsss(0)='1'  OR cVar2S6S46P034P011P066nsss(0)='1'  OR cVar2S7S46P034P014P065nsss(0)='1'  )then
          oVar1S409(0) <='1';
          else
          oVar1S409(0) <='0';
          end if;
        if(cVar2S8S46P034P014P033nsss(0)='1'  OR cVar2S9S46P019P050nsss(0)='1'  OR cVar2S10S46P019N050P015nsss(0)='1'  OR cVar2S11S46P046P034nsss(0)='1'  )then
          oVar1S410(0) <='1';
          else
          oVar1S410(0) <='0';
          end if;
        if(cVar2S12S46N046P017P002nsss(0)='1'  OR cVar2S13S46N046N017P054nsss(0)='1'  OR cVar2S14S46P067P029P050nsss(0)='1'  OR cVar2S15S46N067P064P068nsss(0)='1'  )then
          oVar1S411(0) <='1';
          else
          oVar1S411(0) <='0';
          end if;
        if(cVar2S16S46N067N064P006nsss(0)='1'  OR cVar2S17S46P005P037nsss(0)='1'  OR cVar2S18S46P005N037P015nsss(0)='1'  OR cVar2S19S46P011P014nsss(0)='1'  )then
          oVar1S412(0) <='1';
          else
          oVar1S412(0) <='0';
          end if;
        if(cVar2S20S46P056P037P048nsss(0)='1'  OR cVar2S21S46P056P037P064nsss(0)='1'  OR cVar2S22S46P056P065P031nsss(0)='1'  OR cVar2S23S46P056P065P029nsss(0)='1'  )then
          oVar1S413(0) <='1';
          else
          oVar1S413(0) <='0';
          end if;
        if(cVar2S24S46P064P012nsss(0)='1'  OR cVar2S25S46P064P062P009nsss(0)='1'  OR cVar2S26S46P062P015P060nsss(0)='1'  OR cVar2S27S46P062P015P035nsss(0)='1'  )then
          oVar1S414(0) <='1';
          else
          oVar1S414(0) <='0';
          end if;
        if(cVar2S28S46P062P068P064nsss(0)='1'  OR cVar2S29S46P015P066P029nsss(0)='1'  OR cVar2S30S46P015P066P063nsss(0)='1'  OR cVar2S31S46N015P019P062nsss(0)='1'  )then
          oVar1S415(0) <='1';
          else
          oVar1S415(0) <='0';
          end if;
        if(cVar2S32S46N015N019P009nsss(0)='1'  )then
          oVar1S416(0) <='1';
          else
          oVar1S416(0) <='0';
          end if;
        if(cVar2S0S47P048P031nsss(0)='1'  OR cVar2S1S47P048P018nsss(0)='1'  OR cVar2S2S47P048N018P019nsss(0)='1'  OR cVar2S3S47P027P048P034nsss(0)='1'  )then
          oVar1S417(0) <='1';
          else
          oVar1S417(0) <='0';
          end if;
        if(cVar2S4S47P027N048P068nsss(0)='1'  OR cVar2S5S47N027P051nsss(0)='1'  OR cVar2S6S47N027N051P026nsss(0)='1'  OR cVar2S7S47P047P013P056nsss(0)='1'  )then
          oVar1S418(0) <='1';
          else
          oVar1S418(0) <='0';
          end if;
        if(cVar2S8S47P047N013P055nsss(0)='1'  OR cVar2S9S47P047P035P066nsss(0)='1'  OR cVar2S10S47P046P025nsss(0)='1'  OR cVar2S11S47P046N025P017nsss(0)='1'  )then
          oVar1S419(0) <='1';
          else
          oVar1S419(0) <='0';
          end if;
        if(cVar2S12S47P001P036nsss(0)='1'  OR cVar2S13S47P001N036P032nsss(0)='1'  OR cVar2S14S47P065P014nsss(0)='1'  OR cVar2S15S47P065N014P036nsss(0)='1'  )then
          oVar1S420(0) <='1';
          else
          oVar1S420(0) <='0';
          end if;
        if(cVar2S16S47N065P035P014nsss(0)='1'  OR cVar2S17S47P055nsss(0)='1'  OR cVar2S18S47N055P010P013nsss(0)='1'  OR cVar2S19S47P018P036nsss(0)='1'  )then
          oVar1S421(0) <='1';
          else
          oVar1S421(0) <='0';
          end if;
        if(cVar2S20S47P018N036P015nsss(0)='1'  OR cVar2S21S47P018P019nsss(0)='1'  OR cVar2S22S47P018P012P060nsss(0)='1'  OR cVar2S23S47P018N012P032nsss(0)='1'  )then
          oVar1S422(0) <='1';
          else
          oVar1S422(0) <='0';
          end if;
        if(cVar2S24S47N018P013nsss(0)='1'  OR cVar2S25S47P032P061nsss(0)='1'  OR cVar2S26S47P032N061P066nsss(0)='1'  OR cVar2S27S47N032P059P030nsss(0)='1'  )then
          oVar1S423(0) <='1';
          else
          oVar1S423(0) <='0';
          end if;
        if(cVar2S28S47P018P032P010nsss(0)='1'  OR cVar2S29S47N018P061nsss(0)='1'  OR cVar2S30S47P064P037nsss(0)='1'  OR cVar2S31S47P064P019P017nsss(0)='1'  )then
          oVar1S424(0) <='1';
          else
          oVar1S424(0) <='0';
          end if;
        if(cVar2S32S47P037P010nsss(0)='1'  OR cVar2S33S47N037P013P068nsss(0)='1'  )then
          oVar1S425(0) <='1';
          else
          oVar1S425(0) <='0';
          end if;
        if(cVar2S0S48P012P063P007nsss(0)='1'  OR cVar2S1S48P012P019nsss(0)='1'  OR cVar2S2S48P069P041P036nsss(0)='1'  OR cVar2S3S48P069N041P005nsss(0)='1'  )then
          oVar1S426(0) <='1';
          else
          oVar1S426(0) <='0';
          end if;
        if(cVar2S4S48N069P046P016nsss(0)='1'  OR cVar2S5S48P066P059P063nsss(0)='1'  OR cVar2S6S48P066P059P014nsss(0)='1'  OR cVar2S7S48P066P059nsss(0)='1'  )then
          oVar1S427(0) <='1';
          else
          oVar1S427(0) <='0';
          end if;
        if(cVar2S8S48P066N059P014nsss(0)='1'  OR cVar2S9S48P030P019nsss(0)='1'  OR cVar2S10S48P030nsss(0)='1'  OR cVar2S11S48N030P053nsss(0)='1'  )then
          oVar1S428(0) <='1';
          else
          oVar1S428(0) <='0';
          end if;
        if(cVar2S12S48N030P053P009nsss(0)='1'  OR cVar2S13S48P008P065P048nsss(0)='1'  OR cVar2S14S48N008P066P018nsss(0)='1'  OR cVar2S15S48P002P006nsss(0)='1'  )then
          oVar1S429(0) <='1';
          else
          oVar1S429(0) <='0';
          end if;
        if(cVar2S16S48P002P006P051nsss(0)='1'  OR cVar2S17S48P002P030nsss(0)='1'  OR cVar2S18S48P025P007P042nsss(0)='1'  OR cVar2S19S48P025N007P061nsss(0)='1'  )then
          oVar1S430(0) <='1';
          else
          oVar1S430(0) <='0';
          end if;
        if(cVar2S20S48N025P048P026nsss(0)='1'  OR cVar2S21S48N025P048P006nsss(0)='1'  OR cVar2S22S48P016nsss(0)='1'  OR cVar2S23S48N016P018nsss(0)='1'  )then
          oVar1S431(0) <='1';
          else
          oVar1S431(0) <='0';
          end if;
        if(cVar2S24S48P041P033P007nsss(0)='1'  OR cVar1S25S48N067P036P005P032nsss(0)='1'  OR cVar2S26S48P061nsss(0)='1'  OR cVar2S27S48N061P033P010nsss(0)='1'  )then
          oVar1S432(0) <='1';
          else
          oVar1S432(0) <='0';
          end if;
        if(cVar2S0S49P028P019nsss(0)='1'  OR cVar2S1S49P028N019P064nsss(0)='1'  OR cVar2S2S49N028psss(0)='1'  OR cVar2S3S49P015P032P059nsss(0)='1'  )then
          oVar1S434(0) <='1';
          else
          oVar1S434(0) <='0';
          end if;
        if(cVar2S4S49P015N032P068nsss(0)='1'  OR cVar2S5S49N015P007P035nsss(0)='1'  OR cVar1S6S49P036P011P010P042nsss(0)='1'  OR cVar2S7S49P066P005P017nsss(0)='1'  )then
          oVar1S435(0) <='1';
          else
          oVar1S435(0) <='0';
          end if;
        if(cVar2S8S49P066P056P069nsss(0)='1'  OR cVar2S9S49P020nsss(0)='1'  OR cVar2S10S49N020P016nsss(0)='1'  OR cVar2S11S49N020N016P021nsss(0)='1'  )then
          oVar1S436(0) <='1';
          else
          oVar1S436(0) <='0';
          end if;
        if(cVar2S12S49P050P019nsss(0)='1'  OR cVar2S13S49N050P055P061nsss(0)='1'  OR cVar2S14S49P015P054nsss(0)='1'  OR cVar2S15S49P015N054P013nsss(0)='1'  )then
          oVar1S437(0) <='1';
          else
          oVar1S437(0) <='0';
          end if;
        if(cVar2S16S49N015P009P064nsss(0)='1'  OR cVar2S17S49N015N009P013nsss(0)='1'  OR cVar2S18S49P067P068nsss(0)='1'  OR cVar2S19S49P067N068P056nsss(0)='1'  )then
          oVar1S438(0) <='1';
          else
          oVar1S438(0) <='0';
          end if;
        if(cVar2S20S49N067P002P004nsss(0)='1'  OR cVar1S21S49P036P043P022nsss(0)='1'  OR cVar2S22S49P016nsss(0)='1'  OR cVar2S23S49N016P019nsss(0)='1'  )then
          oVar1S439(0) <='1';
          else
          oVar1S439(0) <='0';
          end if;
        if(cVar2S24S49N016N019P069nsss(0)='1'  OR cVar2S25S49P065P022P038nsss(0)='1'  OR cVar2S26S49P065P032P019nsss(0)='1'  OR cVar2S27S49P014P065nsss(0)='1'  )then
          oVar1S440(0) <='1';
          else
          oVar1S440(0) <='0';
          end if;
        if(cVar2S28S49P014N065P035nsss(0)='1'  OR cVar2S29S49N014P068P033nsss(0)='1'  OR cVar2S30S49P037nsss(0)='1'  )then
          oVar1S441(0) <='1';
          else
          oVar1S441(0) <='0';
          end if;
        if(cVar2S0S50P002nsss(0)='1'  OR cVar2S1S50N002P004P021nsss(0)='1'  OR cVar2S2S50N002N004P039nsss(0)='1'  OR cVar2S3S50P023P042P040nsss(0)='1'  )then
          oVar1S442(0) <='1';
          else
          oVar1S442(0) <='0';
          end if;
        if(cVar2S4S50P023N042P045nsss(0)='1'  OR cVar2S5S50N023P044nsss(0)='1'  OR cVar2S6S50N023P044P053nsss(0)='1'  OR cVar2S7S50P028P010nsss(0)='1'  )then
          oVar1S443(0) <='1';
          else
          oVar1S443(0) <='0';
          end if;
        if(cVar2S8S50P028N010P011nsss(0)='1'  OR cVar2S9S50N028P063nsss(0)='1'  OR cVar2S10S50N028N063P013nsss(0)='1'  OR cVar2S11S50P007nsss(0)='1'  )then
          oVar1S444(0) <='1';
          else
          oVar1S444(0) <='0';
          end if;
        if(cVar2S12S50N007P047P009nsss(0)='1'  OR cVar2S13S50P056P008P055nsss(0)='1'  OR cVar2S14S50N056P031P003nsss(0)='1'  OR cVar2S15S50N056P031P034nsss(0)='1'  )then
          oVar1S445(0) <='1';
          else
          oVar1S445(0) <='0';
          end if;
        if(cVar2S16S50P009P058nsss(0)='1'  OR cVar1S17S50P036P033P026P047nsss(0)='1'  OR cVar2S18S50P054P004P018nsss(0)='1'  OR cVar2S19S50P050P026P012nsss(0)='1'  )then
          oVar1S446(0) <='1';
          else
          oVar1S446(0) <='0';
          end if;
        if(cVar2S20S50P012nsss(0)='1'  OR cVar2S21S50N012P016P058nsss(0)='1'  OR cVar2S22S50N012N016P033nsss(0)='1'  OR cVar2S23S50P037P066P067nsss(0)='1'  )then
          oVar1S447(0) <='1';
          else
          oVar1S447(0) <='0';
          end if;
        if(cVar2S24S50P037N066P069nsss(0)='1'  OR cVar2S25S50P000P010P069nsss(0)='1'  OR cVar2S26S50N000P008P009nsss(0)='1'  OR cVar1S27S50P036P068P019P025nsss(0)='1'  )then
          oVar1S448(0) <='1';
          else
          oVar1S448(0) <='0';
          end if;
        if(cVar2S28S50P005P054nsss(0)='1'  OR cVar2S29S50P005N054P018nsss(0)='1'  OR cVar2S30S50P037P018nsss(0)='1'  OR cVar2S31S50P037N018P017nsss(0)='1'  )then
          oVar1S449(0) <='1';
          else
          oVar1S449(0) <='0';
          end if;
        if(cVar2S32S50N037P012P017nsss(0)='1'  OR cVar2S33S50N037P012P035nsss(0)='1'  OR cVar2S34S50P065P069nsss(0)='1'  )then
          oVar1S450(0) <='1';
          else
          oVar1S450(0) <='0';
          end if;
        if(cVar2S0S51P068P050nsss(0)='1'  OR cVar2S1S51P068P060nsss(0)='1'  OR cVar2S2S51P061P064nsss(0)='1'  OR cVar2S3S51P061N064P016nsss(0)='1'  )then
          oVar1S451(0) <='1';
          else
          oVar1S451(0) <='0';
          end if;
        if(cVar2S4S51P061P068nsss(0)='1'  OR cVar2S5S51P014nsss(0)='1'  OR cVar2S6S51P014P037P029nsss(0)='1'  OR cVar2S7S51P006P051P062nsss(0)='1'  )then
          oVar1S452(0) <='1';
          else
          oVar1S452(0) <='0';
          end if;
        if(cVar2S8S51P006N051P056nsss(0)='1'  OR cVar2S9S51P006P067P019nsss(0)='1'  OR cVar2S10S51P018P014nsss(0)='1'  OR cVar2S11S51P018P014P068nsss(0)='1'  )then
          oVar1S453(0) <='1';
          else
          oVar1S453(0) <='0';
          end if;
        if(cVar2S12S51N018P007P016nsss(0)='1'  OR cVar2S13S51N018N007P009nsss(0)='1'  OR cVar2S14S51P046P042P052nsss(0)='1'  OR cVar2S15S51N046P040nsss(0)='1'  )then
          oVar1S454(0) <='1';
          else
          oVar1S454(0) <='0';
          end if;
        if(cVar2S16S51N046N040P044nsss(0)='1'  OR cVar2S17S51P062P017P057nsss(0)='1'  OR cVar2S18S51P062N017P014nsss(0)='1'  OR cVar2S19S51P062P069nsss(0)='1'  )then
          oVar1S455(0) <='1';
          else
          oVar1S455(0) <='0';
          end if;
        if(cVar2S20S51P030P055nsss(0)='1'  OR cVar2S21S51P030P055P012nsss(0)='1'  OR cVar2S22S51N030P034P060nsss(0)='1'  OR cVar2S23S51N030N034P008nsss(0)='1'  )then
          oVar1S456(0) <='1';
          else
          oVar1S456(0) <='0';
          end if;
        if(cVar2S24S51P011P030nsss(0)='1'  OR cVar2S25S51P011P054nsss(0)='1'  OR cVar2S26S51P057P013nsss(0)='1'  OR cVar2S27S51P057N013P054nsss(0)='1'  )then
          oVar1S457(0) <='1';
          else
          oVar1S457(0) <='0';
          end if;
        if(cVar2S28S51P065P017nsss(0)='1'  OR cVar1S29S51P033N056P006P042nsss(0)='1'  OR cVar2S30S51P028nsss(0)='1'  OR cVar2S31S51N028P012P059nsss(0)='1'  )then
          oVar1S458(0) <='1';
          else
          oVar1S458(0) <='0';
          end if;
        if(cVar2S0S52P049P056nsss(0)='1'  OR cVar2S1S52P049P056P035nsss(0)='1'  OR cVar2S2S52P003P069nsss(0)='1'  OR cVar2S3S52N003P046nsss(0)='1'  )then
          oVar1S460(0) <='1';
          else
          oVar1S460(0) <='0';
          end if;
        if(cVar2S4S52N003N046P062nsss(0)='1'  OR cVar2S5S52P013P030nsss(0)='1'  OR cVar2S6S52P013P030P062nsss(0)='1'  OR cVar2S7S52P013P003P031nsss(0)='1'  )then
          oVar1S461(0) <='1';
          else
          oVar1S461(0) <='0';
          end if;
        if(cVar2S8S52P027nsss(0)='1'  OR cVar2S9S52N027P024nsss(0)='1'  OR cVar2S10S52P014P015nsss(0)='1'  OR cVar2S11S52P014P015P058nsss(0)='1'  )then
          oVar1S462(0) <='1';
          else
          oVar1S462(0) <='0';
          end if;
        if(cVar2S12S52N014P007P015nsss(0)='1'  OR cVar2S13S52N014N007P016nsss(0)='1'  OR cVar2S14S52P004P036P045nsss(0)='1'  OR cVar2S15S52N004P005P067nsss(0)='1'  )then
          oVar1S463(0) <='1';
          else
          oVar1S463(0) <='0';
          end if;
        if(cVar2S16S52P033nsss(0)='1'  OR cVar2S17S52N033P032P049nsss(0)='1'  OR cVar2S18S52P064P012P054nsss(0)='1'  OR cVar2S19S52P064P014P015nsss(0)='1'  )then
          oVar1S464(0) <='1';
          else
          oVar1S464(0) <='0';
          end if;
        if(cVar1S20S52P006P042P044nsss(0)='1'  OR cVar1S21S52P006P042N044P019nsss(0)='1'  OR cVar2S22S52P009nsss(0)='1'  OR cVar2S23S52N009P024P046nsss(0)='1'  )then
          oVar1S465(0) <='1';
          else
          oVar1S465(0) <='0';
          end if;
        if(cVar2S24S52N009N024P048nsss(0)='1'  OR cVar2S25S52P045nsss(0)='1'  OR cVar2S26S52P051P036P037nsss(0)='1'  OR cVar2S27S52N051P033P058nsss(0)='1'  )then
          oVar1S466(0) <='1';
          else
          oVar1S466(0) <='0';
          end if;
        if(cVar2S0S53P029P030nsss(0)='1'  OR cVar2S1S53P029P030P012nsss(0)='1'  OR cVar2S2S53N029P019P044nsss(0)='1'  OR cVar2S3S53N029N019psss(0)='1'  )then
          oVar1S468(0) <='1';
          else
          oVar1S468(0) <='0';
          end if;
        if(cVar2S4S53P018P010P036nsss(0)='1'  OR cVar2S5S53N018P054nsss(0)='1'  OR cVar2S6S53N018N054P053nsss(0)='1'  OR cVar2S7S53P019P018P035nsss(0)='1'  )then
          oVar1S469(0) <='1';
          else
          oVar1S469(0) <='0';
          end if;
        if(cVar2S8S53P019N018P037nsss(0)='1'  OR cVar2S9S53P019P018nsss(0)='1'  OR cVar2S10S53P019P018P004nsss(0)='1'  OR cVar2S11S53P066P034nsss(0)='1'  )then
          oVar1S470(0) <='1';
          else
          oVar1S470(0) <='0';
          end if;
        if(cVar2S12S53P066P034P012nsss(0)='1'  OR cVar2S13S53N066P053nsss(0)='1'  OR cVar2S14S53N066N053P049nsss(0)='1'  OR cVar2S15S53P033nsss(0)='1'  )then
          oVar1S471(0) <='1';
          else
          oVar1S471(0) <='0';
          end if;
        if(cVar2S16S53N033P061nsss(0)='1'  OR cVar2S17S53N033N061P018nsss(0)='1'  OR cVar2S18S53P058P069nsss(0)='1'  OR cVar2S19S53P058P069P013nsss(0)='1'  )then
          oVar1S472(0) <='1';
          else
          oVar1S472(0) <='0';
          end if;
        if(cVar2S20S53P058P034P037nsss(0)='1'  OR cVar2S21S53P062P061nsss(0)='1'  OR cVar2S22S53P062N061P050nsss(0)='1'  OR cVar2S23S53P062P013P032nsss(0)='1'  )then
          oVar1S473(0) <='1';
          else
          oVar1S473(0) <='0';
          end if;
        if(cVar2S24S53P062N013P011nsss(0)='1'  OR cVar2S25S53P014P061nsss(0)='1'  OR cVar2S26S53P054P060P035nsss(0)='1'  OR cVar2S27S53P054N060P037nsss(0)='1'  )then
          oVar1S474(0) <='1';
          else
          oVar1S474(0) <='0';
          end if;
        if(cVar2S28S53P054P035P056nsss(0)='1'  OR cVar2S29S53P054N035P010nsss(0)='1'  OR cVar2S30S53P026P005P066nsss(0)='1'  OR cVar2S31S53P033P065nsss(0)='1'  )then
          oVar1S475(0) <='1';
          else
          oVar1S475(0) <='0';
          end if;
        if(cVar2S32S53P033N065P007nsss(0)='1'  OR cVar2S33S53P062P063nsss(0)='1'  OR cVar2S34S53N062P061P008nsss(0)='1'  OR cVar2S35S53P008nsss(0)='1'  )then
          oVar1S476(0) <='1';
          else
          oVar1S476(0) <='0';
          end if;
        if(cVar2S36S53N008P069nsss(0)='1'  OR cVar2S37S53N008N069P066nsss(0)='1'  )then
          oVar1S477(0) <='1';
          else
          oVar1S477(0) <='0';
          end if;
        if(cVar2S0S54P036P044P012nsss(0)='1'  OR cVar2S1S54N036P004P040nsss(0)='1'  OR cVar2S2S54N036P004P042nsss(0)='1'  OR cVar2S3S54P024P023nsss(0)='1'  )then
          oVar1S478(0) <='1';
          else
          oVar1S478(0) <='0';
          end if;
        if(cVar2S4S54P024N023P029nsss(0)='1'  OR cVar2S5S54P069nsss(0)='1'  OR cVar2S6S54N069P040P018nsss(0)='1'  OR cVar2S7S54P032P002nsss(0)='1'  )then
          oVar1S479(0) <='1';
          else
          oVar1S479(0) <='0';
          end if;
        if(cVar2S8S54P032P015P014nsss(0)='1'  OR cVar2S9S54P048P052nsss(0)='1'  OR cVar2S10S54P020P005nsss(0)='1'  OR cVar2S11S54P020N005P038nsss(0)='1'  )then
          oVar1S480(0) <='1';
          else
          oVar1S480(0) <='0';
          end if;
        if(cVar2S12S54N020P008P067nsss(0)='1'  OR cVar2S13S54P051P064nsss(0)='1'  OR cVar2S14S54N051P017P018nsss(0)='1'  OR cVar2S15S54P000P009nsss(0)='1'  )then
          oVar1S481(0) <='1';
          else
          oVar1S481(0) <='0';
          end if;
        if(cVar2S16S54N000P016P017nsss(0)='1'  OR cVar2S17S54N000P016P069nsss(0)='1'  OR cVar2S18S54P013P062nsss(0)='1'  OR cVar2S19S54P013N062P015nsss(0)='1'  )then
          oVar1S482(0) <='1';
          else
          oVar1S482(0) <='0';
          end if;
        if(cVar2S20S54N013P019P015nsss(0)='1'  OR cVar2S21S54P059nsss(0)='1'  OR cVar2S22S54N059P063nsss(0)='1'  OR cVar2S23S54N059N063P009nsss(0)='1'  )then
          oVar1S483(0) <='1';
          else
          oVar1S483(0) <='0';
          end if;
        if(cVar2S24S54P014P015nsss(0)='1'  OR cVar2S25S54P036P007P004nsss(0)='1'  OR cVar2S26S54P036P007P066nsss(0)='1'  OR cVar2S27S54P036P010P019nsss(0)='1'  )then
          oVar1S484(0) <='1';
          else
          oVar1S484(0) <='0';
          end if;
        if(cVar2S28S54P012P066nsss(0)='1'  OR cVar2S29S54P012N066P014nsss(0)='1'  OR cVar2S30S54N012P010nsss(0)='1'  OR cVar2S31S54N012N010P032nsss(0)='1'  )then
          oVar1S485(0) <='1';
          else
          oVar1S485(0) <='0';
          end if;
        if(cVar2S32S54P034P006P005nsss(0)='1'  OR cVar2S33S54N034P063P069nsss(0)='1'  OR cVar2S34S54P025nsss(0)='1'  OR cVar2S35S54N025P004P014nsss(0)='1'  )then
          oVar1S486(0) <='1';
          else
          oVar1S486(0) <='0';
          end if;
        if(cVar2S0S55P041P065nsss(0)='1'  OR cVar2S1S55P041P065P018nsss(0)='1'  OR cVar2S2S55N041P003P020nsss(0)='1'  OR cVar2S3S55N041P003P043nsss(0)='1'  )then
          oVar1S488(0) <='1';
          else
          oVar1S488(0) <='0';
          end if;
        if(cVar2S4S55P067P010P065nsss(0)='1'  OR cVar2S5S55P035P024nsss(0)='1'  OR cVar2S6S55N035P058P033nsss(0)='1'  OR cVar2S7S55P026nsss(0)='1'  )then
          oVar1S489(0) <='1';
          else
          oVar1S489(0) <='0';
          end if;
        if(cVar1S8S55P016P037P017P008nsss(0)='1'  OR cVar2S9S55P067P035P068nsss(0)='1'  OR cVar2S10S55P067N035P068nsss(0)='1'  OR cVar2S11S55P067P062P064nsss(0)='1'  )then
          oVar1S490(0) <='1';
          else
          oVar1S490(0) <='0';
          end if;
        if(cVar2S12S55P067N062P014nsss(0)='1'  OR cVar2S13S55P063P048nsss(0)='1'  OR cVar2S14S55P063P034P066nsss(0)='1'  OR cVar2S15S55P019P015P034nsss(0)='1'  )then
          oVar1S491(0) <='1';
          else
          oVar1S491(0) <='0';
          end if;
        if(cVar2S16S55P019P015P013nsss(0)='1'  OR cVar2S17S55N019P065P004nsss(0)='1'  OR cVar2S18S55P046P055P034nsss(0)='1'  OR cVar2S19S55P046N055P027nsss(0)='1'  )then
          oVar1S492(0) <='1';
          else
          oVar1S492(0) <='0';
          end if;
        if(cVar2S20S55P046P019nsss(0)='1'  OR cVar2S21S55P010P065nsss(0)='1'  OR cVar2S22S55P010N065P067nsss(0)='1'  OR cVar2S23S55N010P029P062nsss(0)='1'  )then
          oVar1S493(0) <='1';
          else
          oVar1S493(0) <='0';
          end if;
        if(cVar1S24S55P016N036P046P024nsss(0)='1'  OR cVar2S25S55P047P018nsss(0)='1'  OR cVar2S26S55P047P018P037nsss(0)='1'  OR cVar2S27S55P054P000P042nsss(0)='1'  )then
          oVar1S494(0) <='1';
          else
          oVar1S494(0) <='0';
          end if;
        if(cVar2S28S55P054P035P013nsss(0)='1'  OR cVar2S29S55P054N035P010nsss(0)='1'  OR cVar2S30S55P006nsss(0)='1'  OR cVar2S31S55N006P008nsss(0)='1'  )then
          oVar1S495(0) <='1';
          else
          oVar1S495(0) <='0';
          end if;
        if(cVar2S0S56P060P040P048nsss(0)='1'  OR cVar2S1S56N060P058P031nsss(0)='1'  OR cVar2S2S56N060P058P057nsss(0)='1'  OR cVar2S3S56P062P017nsss(0)='1'  )then
          oVar1S497(0) <='1';
          else
          oVar1S497(0) <='0';
          end if;
        if(cVar2S4S56N062P065P037nsss(0)='1'  OR cVar2S5S56P037P065nsss(0)='1'  OR cVar2S6S56P037P065P018nsss(0)='1'  OR cVar2S7S56P037P065nsss(0)='1'  )then
          oVar1S498(0) <='1';
          else
          oVar1S498(0) <='0';
          end if;
        if(cVar2S8S56P066P013nsss(0)='1'  OR cVar2S9S56P066N013P019nsss(0)='1'  OR cVar1S10S56P016P036P043P015nsss(0)='1'  OR cVar2S11S56P020P055P059nsss(0)='1'  )then
          oVar1S499(0) <='1';
          else
          oVar1S499(0) <='0';
          end if;
        if(cVar2S12S56P062P014nsss(0)='1'  OR cVar2S13S56N062P003nsss(0)='1'  OR cVar2S14S56P060nsss(0)='1'  OR cVar2S15S56P060P011nsss(0)='1'  )then
          oVar1S500(0) <='1';
          else
          oVar1S500(0) <='0';
          end if;
        if(cVar2S16S56P056P066nsss(0)='1'  OR cVar2S17S56P056N066P064nsss(0)='1'  OR cVar2S18S56P059nsss(0)='1'  OR cVar2S19S56N059P018P049nsss(0)='1'  )then
          oVar1S501(0) <='1';
          else
          oVar1S501(0) <='0';
          end if;
        if(cVar2S20S56P060P013nsss(0)='1'  OR cVar2S21S56P060N013P052nsss(0)='1'  OR cVar2S22S56P060P015nsss(0)='1'  OR cVar2S23S56P051nsss(0)='1'  )then
          oVar1S502(0) <='1';
          else
          oVar1S502(0) <='0';
          end if;
        if(cVar2S24S56P051P017nsss(0)='1'  OR cVar2S25S56P051P069nsss(0)='1'  OR cVar2S26S56N051P036nsss(0)='1'  OR cVar2S27S56N051N036P034nsss(0)='1'  )then
          oVar1S503(0) <='1';
          else
          oVar1S503(0) <='0';
          end if;
        if(cVar2S28S56P049P026P011nsss(0)='1'  OR cVar2S29S56P049N026P034nsss(0)='1'  )then
          oVar1S504(0) <='1';
          else
          oVar1S504(0) <='0';
          end if;
        if(cVar2S0S57P020P005P013nsss(0)='1'  OR cVar2S1S57P020N005P017nsss(0)='1'  OR cVar2S2S57N020P019P041nsss(0)='1'  OR cVar2S3S57N020N019P017nsss(0)='1'  )then
          oVar1S505(0) <='1';
          else
          oVar1S505(0) <='0';
          end if;
        if(cVar2S4S57P028P055P057nsss(0)='1'  OR cVar2S5S57N028P029P018nsss(0)='1'  OR cVar2S6S57P005P020P019nsss(0)='1'  OR cVar2S7S57P005P062P014nsss(0)='1'  )then
          oVar1S506(0) <='1';
          else
          oVar1S506(0) <='0';
          end if;
        if(cVar2S8S57P005N062P010nsss(0)='1'  OR cVar2S9S57P054P060P008nsss(0)='1'  OR cVar2S10S57P054N060P057nsss(0)='1'  OR cVar2S11S57P054P014P017nsss(0)='1'  )then
          oVar1S507(0) <='1';
          else
          oVar1S507(0) <='0';
          end if;
        if(cVar2S12S57P054N014P034nsss(0)='1'  OR cVar2S13S57P026nsss(0)='1'  OR cVar2S14S57N026P019nsss(0)='1'  OR cVar2S15S57P067nsss(0)='1'  )then
          oVar1S508(0) <='1';
          else
          oVar1S508(0) <='0';
          end if;
        if(cVar2S16S57N067P055nsss(0)='1'  OR cVar2S17S57N067N055P059nsss(0)='1'  OR cVar2S18S57P016P059P033nsss(0)='1'  OR cVar2S19S57N016P015P018nsss(0)='1'  )then
          oVar1S509(0) <='1';
          else
          oVar1S509(0) <='0';
          end if;
        if(cVar2S20S57P068P035P013nsss(0)='1'  OR cVar2S21S57P068N035P026nsss(0)='1'  OR cVar2S22S57P005P035nsss(0)='1'  OR cVar2S23S57P005N035P033nsss(0)='1'  )then
          oVar1S510(0) <='1';
          else
          oVar1S510(0) <='0';
          end if;
        if(cVar2S24S57P005P009P064nsss(0)='1'  OR cVar2S25S57P035nsss(0)='1'  OR cVar1S26S57P056P052P009nsss(0)='1'  OR cVar1S27S57P056P052N009P008nsss(0)='1'  )then
          oVar1S511(0) <='1';
          else
          oVar1S511(0) <='0';
          end if;
        if(cVar2S28S57P012P050nsss(0)='1'  )then
          oVar1S512(0) <='1';
          else
          oVar1S512(0) <='0';
          end if;
        if(cVar2S0S58P005nsss(0)='1'  OR cVar2S1S58N005P023nsss(0)='1'  OR cVar2S2S58N005N023P004nsss(0)='1'  OR cVar2S3S58P039nsss(0)='1'  )then
          oVar1S513(0) <='1';
          else
          oVar1S513(0) <='0';
          end if;
        if(cVar2S4S58P002nsss(0)='1'  OR cVar2S5S58N002P021nsss(0)='1'  OR cVar2S6S58P015P036nsss(0)='1'  OR cVar2S7S58P015P036P061nsss(0)='1'  )then
          oVar1S514(0) <='1';
          else
          oVar1S514(0) <='0';
          end if;
        if(cVar2S8S58N015P058nsss(0)='1'  OR cVar2S9S58P035P034P013nsss(0)='1'  OR cVar2S10S58P035P034P014nsss(0)='1'  OR cVar2S11S58N035P013nsss(0)='1'  )then
          oVar1S515(0) <='1';
          else
          oVar1S515(0) <='0';
          end if;
        if(cVar2S12S58N035N013P014nsss(0)='1'  OR cVar2S13S58P064P016nsss(0)='1'  OR cVar2S14S58P064P016P013nsss(0)='1'  OR cVar2S15S58N064P037nsss(0)='1'  )then
          oVar1S516(0) <='1';
          else
          oVar1S516(0) <='0';
          end if;
        if(cVar2S16S58P018nsss(0)='1'  OR cVar2S17S58P030P059nsss(0)='1'  OR cVar2S18S58N030P015P036nsss(0)='1'  OR cVar2S19S58N030N015P009nsss(0)='1'  )then
          oVar1S517(0) <='1';
          else
          oVar1S517(0) <='0';
          end if;
        if(cVar2S20S58P035P014P033nsss(0)='1'  OR cVar2S21S58P035N014P063nsss(0)='1'  OR cVar2S22S58N035P014P054nsss(0)='1'  OR cVar2S23S58N035P014P068nsss(0)='1'  )then
          oVar1S518(0) <='1';
          else
          oVar1S518(0) <='0';
          end if;
        if(cVar2S24S58P013P069P062nsss(0)='1'  OR cVar2S25S58P013P069psss(0)='1'  OR cVar2S26S58P013P016nsss(0)='1'  OR cVar2S27S58P046nsss(0)='1'  )then
          oVar1S519(0) <='1';
          else
          oVar1S519(0) <='0';
          end if;
        if(cVar2S28S58P019P033nsss(0)='1'  OR cVar2S29S58P019P033P061nsss(0)='1'  OR cVar2S30S58P019P069P018nsss(0)='1'  OR cVar2S31S58P018P036nsss(0)='1'  )then
          oVar1S520(0) <='1';
          else
          oVar1S520(0) <='0';
          end if;
        if(cVar2S32S58N018P069P016nsss(0)='1'  OR cVar2S33S58P045nsss(0)='1'  OR cVar2S34S58P045P018nsss(0)='1'  OR cVar2S35S58P037P015P004nsss(0)='1'  )then
          oVar1S521(0) <='1';
          else
          oVar1S521(0) <='0';
          end if;
        if(cVar2S36S58N037P047P014nsss(0)='1'  OR cVar2S37S58N037N047P031nsss(0)='1'  )then
          oVar1S522(0) <='1';
          else
          oVar1S522(0) <='0';
          end if;
        if(cVar2S0S59P066P068nsss(0)='1'  OR cVar2S1S59P066N068P056nsss(0)='1'  OR cVar2S2S59P066P019nsss(0)='1'  OR cVar2S3S59P034P017P018nsss(0)='1'  )then
          oVar1S523(0) <='1';
          else
          oVar1S523(0) <='0';
          end if;
        if(cVar2S4S59P034P017P062nsss(0)='1'  OR cVar2S5S59P012P067P010nsss(0)='1'  OR cVar2S6S59P012P067P034nsss(0)='1'  OR cVar2S7S59N012P031P062nsss(0)='1'  )then
          oVar1S524(0) <='1';
          else
          oVar1S524(0) <='0';
          end if;
        if(cVar2S8S59N012P031P065nsss(0)='1'  OR cVar2S9S59P010P054P013nsss(0)='1'  OR cVar2S10S59P017nsss(0)='1'  OR cVar2S11S59P019P035nsss(0)='1'  )then
          oVar1S525(0) <='1';
          else
          oVar1S525(0) <='0';
          end if;
        if(cVar2S12S59P019P035P066nsss(0)='1'  OR cVar2S13S59P019P034P018nsss(0)='1'  OR cVar2S14S59P019N034P033nsss(0)='1'  OR cVar2S15S59P055P061P069nsss(0)='1'  )then
          oVar1S526(0) <='1';
          else
          oVar1S526(0) <='0';
          end if;
        if(cVar2S16S59P067P035nsss(0)='1'  OR cVar2S17S59P010P036nsss(0)='1'  OR cVar2S18S59P051P058P037nsss(0)='1'  OR cVar2S19S59P041P016nsss(0)='1'  )then
          oVar1S527(0) <='1';
          else
          oVar1S527(0) <='0';
          end if;
        if(cVar2S20S59P041P016P013nsss(0)='1'  OR cVar2S21S59N041P038nsss(0)='1'  OR cVar2S22S59P008P019P018nsss(0)='1'  OR cVar2S23S59P008N019P013nsss(0)='1'  )then
          oVar1S528(0) <='1';
          else
          oVar1S528(0) <='0';
          end if;
        if(cVar2S24S59N008P011P017nsss(0)='1'  )then
          oVar1S529(0) <='1';
          else
          oVar1S529(0) <='0';
          end if;
        if(cVar2S0S60P007P035P020nsss(0)='1'  OR cVar2S1S60P007N035P066nsss(0)='1'  OR cVar2S2S60P007P057P064nsss(0)='1'  OR cVar2S3S60P012P048P066nsss(0)='1'  )then
          oVar1S530(0) <='1';
          else
          oVar1S530(0) <='0';
          end if;
        if(cVar2S4S60N012P004nsss(0)='1'  OR cVar2S5S60N012N004P026nsss(0)='1'  OR cVar2S6S60P015P013nsss(0)='1'  OR cVar2S7S60N015P013nsss(0)='1'  )then
          oVar1S531(0) <='1';
          else
          oVar1S531(0) <='0';
          end if;
        if(cVar2S8S60P067P062P060nsss(0)='1'  OR cVar2S9S60P067N062P011nsss(0)='1'  OR cVar2S10S60N067P058P012nsss(0)='1'  OR cVar2S11S60P014P016nsss(0)='1'  )then
          oVar1S532(0) <='1';
          else
          oVar1S532(0) <='0';
          end if;
        if(cVar2S12S60P014N016P017nsss(0)='1'  OR cVar2S13S60P014P011nsss(0)='1'  OR cVar2S14S60P067P065P015nsss(0)='1'  OR cVar2S15S60P067P065P066nsss(0)='1'  )then
          oVar1S533(0) <='1';
          else
          oVar1S533(0) <='0';
          end if;
        if(cVar2S16S60P067P064P016nsss(0)='1'  OR cVar1S17S60P037P063P068P052nsss(0)='1'  OR cVar2S18S60P012P013nsss(0)='1'  OR cVar2S19S60N012P059P033nsss(0)='1'  )then
          oVar1S534(0) <='1';
          else
          oVar1S534(0) <='0';
          end if;
        if(cVar2S20S60P007nsss(0)='1'  OR cVar2S21S60N007P056nsss(0)='1'  OR cVar2S22S60P014P024nsss(0)='1'  OR cVar2S23S60P014N024P015nsss(0)='1'  )then
          oVar1S535(0) <='1';
          else
          oVar1S535(0) <='0';
          end if;
        if(cVar2S24S60P014P023P069nsss(0)='1'  OR cVar2S25S60P036P064nsss(0)='1'  OR cVar2S26S60P036N064P017nsss(0)='1'  OR cVar2S27S60P069P034P017nsss(0)='1'  )then
          oVar1S536(0) <='1';
          else
          oVar1S536(0) <='0';
          end if;
        if(cVar2S28S60P067P036nsss(0)='1'  OR cVar2S29S60P067P036P034nsss(0)='1'  OR cVar2S30S60N067P051P066nsss(0)='1'  OR cVar2S31S60P010nsss(0)='1'  )then
          oVar1S537(0) <='1';
          else
          oVar1S537(0) <='0';
          end if;
        if(cVar2S32S60N010P031P015nsss(0)='1'  OR cVar2S33S60N010N031P062nsss(0)='1'  OR cVar2S34S60P033P060P012nsss(0)='1'  OR cVar2S35S60P033N060P055nsss(0)='1'  )then
          oVar1S538(0) <='1';
          else
          oVar1S538(0) <='0';
          end if;
        if(cVar2S36S60N033P055P031nsss(0)='1'  )then
          oVar1S539(0) <='1';
          else
          oVar1S539(0) <='0';
          end if;
        if(cVar2S0S61P065P055nsss(0)='1'  OR cVar2S1S61P065P055P056nsss(0)='1'  OR cVar2S2S61P065P030nsss(0)='1'  OR cVar2S3S61P065N030P009nsss(0)='1'  )then
          oVar1S540(0) <='1';
          else
          oVar1S540(0) <='0';
          end if;
        if(cVar2S4S61P067P064P068nsss(0)='1'  OR cVar2S5S61P067N064psss(0)='1'  OR cVar2S6S61N067P033P069nsss(0)='1'  OR cVar2S7S61N067P033P028nsss(0)='1'  )then
          oVar1S541(0) <='1';
          else
          oVar1S541(0) <='0';
          end if;
        if(cVar2S8S61P046nsss(0)='1'  OR cVar2S9S61N046P068P019nsss(0)='1'  OR cVar2S10S61P064P061nsss(0)='1'  OR cVar2S11S61P064P037P069nsss(0)='1'  )then
          oVar1S542(0) <='1';
          else
          oVar1S542(0) <='0';
          end if;
        if(cVar2S12S61P064N037P056nsss(0)='1'  OR cVar2S13S61P059P062P055nsss(0)='1'  OR cVar2S14S61P059N062P015nsss(0)='1'  OR cVar2S15S61P059P018P032nsss(0)='1'  )then
          oVar1S543(0) <='1';
          else
          oVar1S543(0) <='0';
          end if;
        if(cVar2S16S61P012P032nsss(0)='1'  OR cVar2S17S61P012P032P016nsss(0)='1'  OR cVar2S18S61P012P018nsss(0)='1'  OR cVar2S19S61P062P056nsss(0)='1'  )then
          oVar1S544(0) <='1';
          else
          oVar1S544(0) <='0';
          end if;
        if(cVar2S20S61N062P049P047nsss(0)='1'  OR cVar2S21S61N062N049P052nsss(0)='1'  OR cVar1S22S61P063P062P068P060nsss(0)='1'  OR cVar2S23S61P067P017nsss(0)='1'  )then
          oVar1S545(0) <='1';
          else
          oVar1S545(0) <='0';
          end if;
        if(cVar2S24S61P067N017P034nsss(0)='1'  OR cVar2S25S61N067P014P018nsss(0)='1'  OR cVar2S26S61P037P034P014nsss(0)='1'  OR cVar2S27S61P037N034P014nsss(0)='1'  )then
          oVar1S546(0) <='1';
          else
          oVar1S546(0) <='0';
          end if;
        if(cVar2S28S61N037P069P067nsss(0)='1'  OR cVar2S29S61N037N069P012nsss(0)='1'  OR cVar2S30S61P007P053P036nsss(0)='1'  OR cVar2S31S61P066P045P025nsss(0)='1'  )then
          oVar1S547(0) <='1';
          else
          oVar1S547(0) <='0';
          end if;
        if(cVar2S32S61P066P052P054nsss(0)='1'  OR cVar2S33S61P019nsss(0)='1'  OR cVar2S34S61P067P066P015nsss(0)='1'  )then
          oVar1S548(0) <='1';
          else
          oVar1S548(0) <='0';
          end if;
        if(cVar2S0S62P016P065nsss(0)='1'  OR cVar2S1S62P016N065P007nsss(0)='1'  OR cVar2S2S62N016P025nsss(0)='1'  OR cVar2S3S62N016N025P010nsss(0)='1'  )then
          oVar1S549(0) <='1';
          else
          oVar1S549(0) <='0';
          end if;
        if(cVar1S4S62P062P017P048P046nsss(0)='1'  OR cVar2S5S62P016P035nsss(0)='1'  OR cVar2S6S62P045P012nsss(0)='1'  OR cVar2S7S62N045P015P049nsss(0)='1'  )then
          oVar1S550(0) <='1';
          else
          oVar1S550(0) <='0';
          end if;
        if(cVar2S8S62N045N015P066nsss(0)='1'  OR cVar2S9S62P039nsss(0)='1'  OR cVar2S10S62N039P014P060nsss(0)='1'  OR cVar1S11S62P062N017P047P026nsss(0)='1'  )then
          oVar1S551(0) <='1';
          else
          oVar1S551(0) <='0';
          end if;
        if(cVar2S12S62P007nsss(0)='1'  OR cVar2S13S62P033P015nsss(0)='1'  OR cVar2S14S62P033P015P035nsss(0)='1'  OR cVar2S15S62P033P058P007nsss(0)='1'  )then
          oVar1S552(0) <='1';
          else
          oVar1S552(0) <='0';
          end if;
        if(cVar2S16S62P015P032P058nsss(0)='1'  OR cVar2S17S62P015P032P012nsss(0)='1'  OR cVar2S18S62N015P032P060nsss(0)='1'  OR cVar2S19S62N015N032P030nsss(0)='1'  )then
          oVar1S553(0) <='1';
          else
          oVar1S553(0) <='0';
          end if;
        if(cVar2S20S62P036P034P015nsss(0)='1'  OR cVar2S21S62P036P034P018nsss(0)='1'  OR cVar2S22S62P036P051nsss(0)='1'  OR cVar2S23S62P058P061P068nsss(0)='1'  )then
          oVar1S554(0) <='1';
          else
          oVar1S554(0) <='0';
          end if;
        if(cVar2S24S62P058P061P032nsss(0)='1'  OR cVar2S25S62N058P055P017nsss(0)='1'  OR cVar2S26S62P063P064P060nsss(0)='1'  OR cVar2S27S62P063P029nsss(0)='1'  )then
          oVar1S555(0) <='1';
          else
          oVar1S555(0) <='0';
          end if;
        if(cVar2S28S62P063N029P053nsss(0)='1'  OR cVar2S29S62P012P048nsss(0)='1'  OR cVar2S30S62P012P048P015nsss(0)='1'  OR cVar2S31S62N012P008P032nsss(0)='1'  )then
          oVar1S556(0) <='1';
          else
          oVar1S556(0) <='0';
          end if;
        if(cVar2S32S62P060P069P042nsss(0)='1'  OR cVar2S33S62P060P011nsss(0)='1'  OR cVar2S34S62P060N011P032nsss(0)='1'  OR cVar2S35S62P067P065nsss(0)='1'  )then
          oVar1S557(0) <='1';
          else
          oVar1S557(0) <='0';
          end if;
        if(cVar2S36S62P067N065P061nsss(0)='1'  OR cVar2S37S62N067P068P019nsss(0)='1'  )then
          oVar1S558(0) <='1';
          else
          oVar1S558(0) <='0';
          end if;
        if(cVar2S0S63P028P017nsss(0)='1'  OR cVar2S1S63P028P017P060nsss(0)='1'  OR cVar2S2S63P028P011P066nsss(0)='1'  OR cVar2S3S63P019P012P010nsss(0)='1'  )then
          oVar1S559(0) <='1';
          else
          oVar1S559(0) <='0';
          end if;
        if(cVar2S4S63N019P013P064nsss(0)='1'  OR cVar2S5S63P017nsss(0)='1'  OR cVar2S6S63P068P029nsss(0)='1'  OR cVar2S7S63P068N029P052nsss(0)='1'  )then
          oVar1S560(0) <='1';
          else
          oVar1S560(0) <='0';
          end if;
        if(cVar2S8S63P040P030P021nsss(0)='1'  OR cVar2S9S63P040P030P015nsss(0)='1'  OR cVar2S10S63P034P064nsss(0)='1'  OR cVar2S11S63P034P064P017nsss(0)='1'  )then
          oVar1S561(0) <='1';
          else
          oVar1S561(0) <='0';
          end if;
        if(cVar2S12S63P034P069P062nsss(0)='1'  OR cVar2S13S63P017P069P003nsss(0)='1'  OR cVar2S14S63N017P045nsss(0)='1'  OR cVar2S15S63N017N045P038nsss(0)='1'  )then
          oVar1S562(0) <='1';
          else
          oVar1S562(0) <='0';
          end if;
        if(cVar1S16S63N067P044P028nsss(0)='1'  OR cVar2S17S63P012nsss(0)='1'  OR cVar2S18S63P025P062nsss(0)='1'  OR cVar2S19S63P025N062P042nsss(0)='1'  )then
          oVar1S563(0) <='1';
          else
          oVar1S563(0) <='0';
          end if;
        if(cVar2S20S63N025P065P017nsss(0)='1'  OR cVar2S21S63N025N065P006nsss(0)='1'  OR cVar2S22S63P010P055P054nsss(0)='1'  OR cVar2S23S63P010P055P034nsss(0)='1'  )then
          oVar1S564(0) <='1';
          else
          oVar1S564(0) <='0';
          end if;
        if(cVar2S24S63P010P024P015nsss(0)='1'  OR cVar2S25S63P051nsss(0)='1'  OR cVar2S26S63P030P013nsss(0)='1'  OR cVar2S27S63P030N013P058nsss(0)='1'  )then
          oVar1S565(0) <='1';
          else
          oVar1S565(0) <='0';
          end if;
        if(cVar2S28S63P030P009P065nsss(0)='1'  OR cVar2S29S63P034P008P062nsss(0)='1'  OR cVar2S30S63P034P008P053nsss(0)='1'  OR cVar2S31S63N034P025P051nsss(0)='1'  )then
          oVar1S566(0) <='1';
          else
          oVar1S566(0) <='0';
          end if;
        if(cVar2S0S64P030P067P018nsss(0)='1'  OR cVar2S1S64P030P067P017nsss(0)='1'  OR cVar2S2S64P062P047P066nsss(0)='1'  OR cVar2S3S64P062N047P026nsss(0)='1'  )then
          oVar1S568(0) <='1';
          else
          oVar1S568(0) <='0';
          end if;
        if(cVar2S4S64P062P006P030nsss(0)='1'  OR cVar2S5S64P060nsss(0)='1'  OR cVar2S6S64P060P062P064nsss(0)='1'  OR cVar2S7S64P032P060P062nsss(0)='1'  )then
          oVar1S569(0) <='1';
          else
          oVar1S569(0) <='0';
          end if;
        if(cVar2S8S64P032N060P055nsss(0)='1'  OR cVar1S9S64P059P061P067P069nsss(0)='1'  OR cVar2S10S64P065P007nsss(0)='1'  OR cVar2S11S64P019nsss(0)='1'  )then
          oVar1S570(0) <='1';
          else
          oVar1S570(0) <='0';
          end if;
        if(cVar2S12S64P013P035nsss(0)='1'  OR cVar2S13S64N013P056nsss(0)='1'  OR cVar2S14S64N013N056P060nsss(0)='1'  OR cVar2S15S64P011P060P061nsss(0)='1'  )then
          oVar1S571(0) <='1';
          else
          oVar1S571(0) <='0';
          end if;
        if(cVar2S16S64P011N060P036nsss(0)='1'  OR cVar2S17S64N011N014P031nsss(0)='1'  OR cVar2S18S64P060nsss(0)='1'  OR cVar2S19S64N060P003nsss(0)='1'  )then
          oVar1S572(0) <='1';
          else
          oVar1S572(0) <='0';
          end if;
        if(cVar1S20S64P059P049P055P051nsss(0)='1'  OR cVar2S21S64P033nsss(0)='1'  )then
          oVar1S573(0) <='1';
          else
          oVar1S573(0) <='0';
          end if;
        if(cVar1S0S65P058P054P047P026nsss(0)='1'  OR cVar2S1S65P037P024P016nsss(0)='1'  OR cVar2S2S65P019P037P035nsss(0)='1'  OR cVar2S3S65P019P037P036nsss(0)='1'  )then
          oVar1S574(0) <='1';
          else
          oVar1S574(0) <='0';
          end if;
        if(cVar2S4S65N019P007P028nsss(0)='1'  OR cVar2S5S65P003P065nsss(0)='1'  OR cVar2S6S65P003N065P009nsss(0)='1'  OR cVar2S7S65N003P009nsss(0)='1'  )then
          oVar1S575(0) <='1';
          else
          oVar1S575(0) <='0';
          end if;
        if(cVar1S8S65P058P054P015P013nsss(0)='1'  OR cVar2S9S65P012P056P033nsss(0)='1'  OR cVar2S10S65P011nsss(0)='1'  OR cVar2S11S65N011P031P013nsss(0)='1'  )then
          oVar1S576(0) <='1';
          else
          oVar1S576(0) <='0';
          end if;
        if(cVar2S12S65P036P068P013nsss(0)='1'  OR cVar1S13S65N058P043P022P003nsss(0)='1'  OR cVar2S14S65P034nsss(0)='1'  OR cVar2S15S65N034P069P064nsss(0)='1'  )then
          oVar1S577(0) <='1';
          else
          oVar1S577(0) <='0';
          end if;
        if(cVar2S16S65P007P016nsss(0)='1'  OR cVar2S17S65P007N016P045nsss(0)='1'  OR cVar2S18S65N007P021nsss(0)='1'  OR cVar2S19S65P036P021nsss(0)='1'  )then
          oVar1S578(0) <='1';
          else
          oVar1S578(0) <='0';
          end if;
        if(cVar2S20S65P036N021P020nsss(0)='1'  OR cVar2S21S65P036psss(0)='1'  OR cVar2S22S65P004P068nsss(0)='1'  OR cVar2S23S65N004P037P062nsss(0)='1'  )then
          oVar1S579(0) <='1';
          else
          oVar1S579(0) <='0';
          end if;
        if(cVar2S24S65P039P020nsss(0)='1'  OR cVar2S25S65P039N020P021nsss(0)='1'  OR cVar2S26S65N039P021P047nsss(0)='1'  OR cVar2S27S65P037P069P066nsss(0)='1'  )then
          oVar1S580(0) <='1';
          else
          oVar1S580(0) <='0';
          end if;
        if(cVar1S0S66P015P044P025nsss(0)='1'  OR cVar1S1S66P015P044N025P023nsss(0)='1'  OR cVar2S2S66P058P022nsss(0)='1'  OR cVar2S3S66P058N022P068nsss(0)='1'  )then
          oVar1S582(0) <='1';
          else
          oVar1S582(0) <='0';
          end if;
        if(cVar2S4S66P035nsss(0)='1'  OR cVar2S5S66P007P005nsss(0)='1'  OR cVar2S6S66P007N005P011nsss(0)='1'  OR cVar2S7S66P007P013P066nsss(0)='1'  )then
          oVar1S583(0) <='1';
          else
          oVar1S583(0) <='0';
          end if;
        if(cVar2S8S66P026P025nsss(0)='1'  OR cVar2S9S66P039P048P006nsss(0)='1'  OR cVar2S10S66P039P048P061nsss(0)='1'  OR cVar2S11S66P039P067nsss(0)='1'  )then
          oVar1S584(0) <='1';
          else
          oVar1S584(0) <='0';
          end if;
        if(cVar2S12S66P032P019nsss(0)='1'  OR cVar2S13S66P032N019P014nsss(0)='1'  OR cVar2S14S66N032psss(0)='1'  OR cVar2S15S66P011P066nsss(0)='1'  )then
          oVar1S585(0) <='1';
          else
          oVar1S585(0) <='0';
          end if;
        if(cVar2S16S66N011P018P035nsss(0)='1'  OR cVar2S17S66P052P059P019nsss(0)='1'  OR cVar2S18S66P052P059P019nsss(0)='1'  OR cVar2S19S66P052P029P050nsss(0)='1'  )then
          oVar1S586(0) <='1';
          else
          oVar1S586(0) <='0';
          end if;
        if(cVar2S20S66P068P018nsss(0)='1'  OR cVar2S21S66P068P018P013nsss(0)='1'  OR cVar2S22S66N068P036P053nsss(0)='1'  OR cVar2S23S66P036P037P055nsss(0)='1'  )then
          oVar1S587(0) <='1';
          else
          oVar1S587(0) <='0';
          end if;
        if(cVar2S24S66P036P037P009nsss(0)='1'  OR cVar2S25S66P036P011nsss(0)='1'  OR cVar2S26S66P036N011P009nsss(0)='1'  OR cVar2S27S66P017P051P033nsss(0)='1'  )then
          oVar1S588(0) <='1';
          else
          oVar1S588(0) <='0';
          end if;
        if(cVar2S28S66P043nsss(0)='1'  OR cVar2S29S66N043P039nsss(0)='1'  OR cVar2S30S66P050P011P014nsss(0)='1'  OR cVar2S31S66P050P011P031nsss(0)='1'  )then
          oVar1S589(0) <='1';
          else
          oVar1S589(0) <='0';
          end if;
        if(cVar2S32S66P050P027P017nsss(0)='1'  OR cVar2S33S66P050N027P026nsss(0)='1'  )then
          oVar1S590(0) <='1';
          else
          oVar1S590(0) <='0';
          end if;
        if(cVar2S0S67P028P034nsss(0)='1'  OR cVar2S1S67P028P034P069nsss(0)='1'  OR cVar2S2S67P028P018nsss(0)='1'  OR cVar2S3S67P028P018P035nsss(0)='1'  )then
          oVar1S591(0) <='1';
          else
          oVar1S591(0) <='0';
          end if;
        if(cVar2S4S67P035P009P010nsss(0)='1'  OR cVar2S5S67N035P020nsss(0)='1'  OR cVar2S6S67N035N020P031nsss(0)='1'  OR cVar2S7S67P035P012nsss(0)='1'  )then
          oVar1S592(0) <='1';
          else
          oVar1S592(0) <='0';
          end if;
        if(cVar2S8S67P035N012P054nsss(0)='1'  OR cVar2S9S67P010P019nsss(0)='1'  OR cVar2S10S67P010N019P054nsss(0)='1'  OR cVar2S11S67N010P027P007nsss(0)='1'  )then
          oVar1S593(0) <='1';
          else
          oVar1S593(0) <='0';
          end if;
        if(cVar2S12S67P033P019P051nsss(0)='1'  OR cVar2S13S67P033P019P056nsss(0)='1'  OR cVar2S14S67N033P057nsss(0)='1'  OR cVar2S15S67N033N057P050nsss(0)='1'  )then
          oVar1S594(0) <='1';
          else
          oVar1S594(0) <='0';
          end if;
        if(cVar2S16S67P009P068nsss(0)='1'  OR cVar2S17S67P009N068P062nsss(0)='1'  OR cVar2S18S67P010P032nsss(0)='1'  OR cVar2S19S67P010N032P008nsss(0)='1'  )then
          oVar1S595(0) <='1';
          else
          oVar1S595(0) <='0';
          end if;
        if(cVar1S20S67P015P044P031P006nsss(0)='1'  OR cVar2S21S67P068nsss(0)='1'  OR cVar2S22S67N068P004nsss(0)='1'  OR cVar1S23S67P015N044P003P055nsss(0)='1'  )then
          oVar1S596(0) <='1';
          else
          oVar1S596(0) <='0';
          end if;
        if(cVar2S24S67P007P005nsss(0)='1'  OR cVar2S25S67P007N005P068nsss(0)='1'  OR cVar2S26S67P007P013P066nsss(0)='1'  OR cVar2S27S67P026P025nsss(0)='1'  )then
          oVar1S597(0) <='1';
          else
          oVar1S597(0) <='0';
          end if;
        if(cVar2S28S67P026P019nsss(0)='1'  OR cVar2S29S67P039P023P018nsss(0)='1'  OR cVar2S30S67P039P023P014nsss(0)='1'  OR cVar2S31S67P039P067nsss(0)='1'  )then
          oVar1S598(0) <='1';
          else
          oVar1S598(0) <='0';
          end if;
        if(cVar2S0S68P062P051nsss(0)='1'  OR cVar2S1S68P062P019nsss(0)='1'  OR cVar2S2S68P062N019P066nsss(0)='1'  OR cVar2S3S68P018P060nsss(0)='1'  )then
          oVar1S600(0) <='1';
          else
          oVar1S600(0) <='0';
          end if;
        if(cVar2S4S68P018N060P009nsss(0)='1'  OR cVar2S5S68P018P023P013nsss(0)='1'  OR cVar2S6S68P018N023P019nsss(0)='1'  OR cVar2S7S68P066P017nsss(0)='1'  )then
          oVar1S601(0) <='1';
          else
          oVar1S601(0) <='0';
          end if;
        if(cVar1S8S68P014P012P001P010nsss(0)='1'  OR cVar2S9S68P034nsss(0)='1'  OR cVar2S10S68N034P009nsss(0)='1'  OR cVar2S11S68P051P066nsss(0)='1'  )then
          oVar1S602(0) <='1';
          else
          oVar1S602(0) <='0';
          end if;
        if(cVar2S12S68P051N066P056nsss(0)='1'  OR cVar2S13S68P051P066P018nsss(0)='1'  OR cVar2S14S68P004P011nsss(0)='1'  OR cVar2S15S68P067P049nsss(0)='1'  )then
          oVar1S603(0) <='1';
          else
          oVar1S603(0) <='0';
          end if;
        if(cVar2S16S68P067N049P018nsss(0)='1'  OR cVar2S17S68N067psss(0)='1'  OR cVar2S18S68P034nsss(0)='1'  OR cVar2S19S68P023P005nsss(0)='1'  )then
          oVar1S604(0) <='1';
          else
          oVar1S604(0) <='0';
          end if;
        if(cVar2S20S68P023N005P008nsss(0)='1'  OR cVar2S21S68P010P015P068nsss(0)='1'  OR cVar2S22S68P001P068nsss(0)='1'  OR cVar2S23S68P001N068P019nsss(0)='1'  )then
          oVar1S605(0) <='1';
          else
          oVar1S605(0) <='0';
          end if;
        if(cVar2S24S68N001P066P013nsss(0)='1'  OR cVar2S25S68N001P066P064nsss(0)='1'  OR cVar2S26S68P062P067P018nsss(0)='1'  OR cVar2S27S68P062P015P013nsss(0)='1'  )then
          oVar1S606(0) <='1';
          else
          oVar1S606(0) <='0';
          end if;
        if(cVar2S28S68P062N015P013nsss(0)='1'  OR cVar2S29S68P005P042P006nsss(0)='1'  OR cVar2S30S68P005P018nsss(0)='1'  OR cVar2S31S68P044P033nsss(0)='1'  )then
          oVar1S607(0) <='1';
          else
          oVar1S607(0) <='0';
          end if;
        if(cVar2S32S68N044P023P045nsss(0)='1'  OR cVar2S33S68N044P023P065nsss(0)='1'  )then
          oVar1S608(0) <='1';
          else
          oVar1S608(0) <='0';
          end if;
        if(cVar2S0S69P063P065nsss(0)='1'  OR cVar2S1S69P063N065P055nsss(0)='1'  OR cVar2S2S69P063P005nsss(0)='1'  OR cVar2S3S69P063N005P048nsss(0)='1'  )then
          oVar1S609(0) <='1';
          else
          oVar1S609(0) <='0';
          end if;
        if(cVar2S4S69P065P019P067nsss(0)='1'  OR cVar2S5S69N065P035P032nsss(0)='1'  OR cVar2S6S69N065N035P030nsss(0)='1'  OR cVar2S7S69P059nsss(0)='1'  )then
          oVar1S610(0) <='1';
          else
          oVar1S610(0) <='0';
          end if;
        if(cVar2S8S69N059P015nsss(0)='1'  OR cVar2S9S69P009P014nsss(0)='1'  OR cVar2S10S69P009P014P016nsss(0)='1'  OR cVar2S11S69N009P036P069nsss(0)='1'  )then
          oVar1S611(0) <='1';
          else
          oVar1S611(0) <='0';
          end if;
        if(cVar2S12S69N009N036P069nsss(0)='1'  OR cVar2S13S69P012P031nsss(0)='1'  OR cVar2S14S69P012N031P029nsss(0)='1'  OR cVar2S15S69N012P026P029nsss(0)='1'  )then
          oVar1S612(0) <='1';
          else
          oVar1S612(0) <='0';
          end if;
        if(cVar2S16S69P040P002nsss(0)='1'  OR cVar2S17S69P040N002P069nsss(0)='1'  OR cVar2S18S69N040P038P047nsss(0)='1'  OR cVar2S19S69P025P068nsss(0)='1'  )then
          oVar1S613(0) <='1';
          else
          oVar1S613(0) <='0';
          end if;
        if(cVar2S20S69P025N068P018nsss(0)='1'  OR cVar2S21S69N025P039P058nsss(0)='1'  OR cVar2S22S69P068P066P007nsss(0)='1'  OR cVar2S23S69P068P016P015nsss(0)='1'  )then
          oVar1S614(0) <='1';
          else
          oVar1S614(0) <='0';
          end if;
        if(cVar2S24S69P051P064nsss(0)='1'  OR cVar2S25S69P051P064P068nsss(0)='1'  OR cVar2S26S69N051P026nsss(0)='1'  OR cVar2S27S69P030P013P018nsss(0)='1'  )then
          oVar1S615(0) <='1';
          else
          oVar1S615(0) <='0';
          end if;
        if(cVar2S28S69P030N013P011nsss(0)='1'  OR cVar2S29S69N030P032nsss(0)='1'  OR cVar2S30S69N030N032P007nsss(0)='1'  OR cVar2S31S69P068P051P055nsss(0)='1'  )then
          oVar1S616(0) <='1';
          else
          oVar1S616(0) <='0';
          end if;
        if(cVar2S32S69P051P026nsss(0)='1'  OR cVar2S33S69P051N026P018nsss(0)='1'  OR cVar2S34S69P051P008nsss(0)='1'  OR cVar2S35S69P024P045nsss(0)='1'  )then
          oVar1S617(0) <='1';
          else
          oVar1S617(0) <='0';
          end if;
        if(cVar2S36S69N024P025nsss(0)='1'  OR cVar2S37S69N024N025P051nsss(0)='1'  OR cVar2S38S69P016nsss(0)='1'  OR cVar2S39S69N016P060nsss(0)='1'  )then
          oVar1S618(0) <='1';
          else
          oVar1S618(0) <='0';
          end if;
        if(cVar2S40S69P042P067P030nsss(0)='1'  OR cVar2S41S69P042N067P046nsss(0)='1'  OR cVar2S42S69P042P021P040nsss(0)='1'  OR cVar2S43S69P042N021P006nsss(0)='1'  )then
          oVar1S619(0) <='1';
          else
          oVar1S619(0) <='0';
          end if;
        if(cVar2S0S70P020P047nsss(0)='1'  OR cVar2S1S70P020N047P012nsss(0)='1'  OR cVar2S2S70P047P007nsss(0)='1'  OR cVar2S3S70P047P006nsss(0)='1'  )then
          oVar1S621(0) <='1';
          else
          oVar1S621(0) <='0';
          end if;
        if(cVar2S4S70P047N006P009nsss(0)='1'  OR cVar2S5S70P010nsss(0)='1'  OR cVar2S6S70P023P040P038nsss(0)='1'  OR cVar2S7S70P023N040P016nsss(0)='1'  )then
          oVar1S622(0) <='1';
          else
          oVar1S622(0) <='0';
          end if;
        if(cVar1S8S70P017P014P012P041nsss(0)='1'  OR cVar2S9S70P039P069P062nsss(0)='1'  OR cVar2S10S70P001nsss(0)='1'  OR cVar2S11S70N001P018P010nsss(0)='1'  )then
          oVar1S623(0) <='1';
          else
          oVar1S623(0) <='0';
          end if;
        if(cVar2S12S70N001N018P019nsss(0)='1'  OR cVar2S13S70P020P052P068nsss(0)='1'  OR cVar2S14S70P020P052P059nsss(0)='1'  OR cVar2S15S70P020P059nsss(0)='1'  )then
          oVar1S624(0) <='1';
          else
          oVar1S624(0) <='0';
          end if;
        if(cVar2S16S70P069P012P067nsss(0)='1'  OR cVar2S17S70N069P029P000nsss(0)='1'  OR cVar2S18S70N069N029P015nsss(0)='1'  OR cVar2S19S70P048P037nsss(0)='1'  )then
          oVar1S625(0) <='1';
          else
          oVar1S625(0) <='0';
          end if;
        if(cVar2S20S70P048N037P023nsss(0)='1'  OR cVar2S21S70P048P046nsss(0)='1'  OR cVar2S22S70P020P032P010nsss(0)='1'  OR cVar2S23S70P020P068nsss(0)='1'  )then
          oVar1S626(0) <='1';
          else
          oVar1S626(0) <='0';
          end if;
        if(cVar2S24S70N020P065P036nsss(0)='1'  OR cVar1S25S70N017P066P004P061nsss(0)='1'  OR cVar2S26S70P042nsss(0)='1'  OR cVar2S27S70N042P037P009nsss(0)='1'  )then
          oVar1S627(0) <='1';
          else
          oVar1S627(0) <='0';
          end if;
        if(cVar2S0S71P016P060nsss(0)='1'  OR cVar2S1S71P016P060P013nsss(0)='1'  OR cVar2S2S71P016P055P007nsss(0)='1'  OR cVar2S3S71P016P055P065nsss(0)='1'  )then
          oVar1S629(0) <='1';
          else
          oVar1S629(0) <='0';
          end if;
        if(cVar2S4S71P019P066P037nsss(0)='1'  OR cVar2S5S71N019P063P016nsss(0)='1'  OR cVar2S6S71P033P021P040nsss(0)='1'  OR cVar2S7S71P033N021P061nsss(0)='1'  )then
          oVar1S630(0) <='1';
          else
          oVar1S630(0) <='0';
          end if;
        if(cVar2S8S71P014P007P013nsss(0)='1'  OR cVar2S9S71P014P007P024nsss(0)='1'  OR cVar2S10S71N014P016P007nsss(0)='1'  OR cVar2S11S71N014N016P012nsss(0)='1'  )then
          oVar1S631(0) <='1';
          else
          oVar1S631(0) <='0';
          end if;
        if(cVar2S12S71P013P019P012nsss(0)='1'  OR cVar2S13S71P013N019P018nsss(0)='1'  OR cVar2S14S71P013P019nsss(0)='1'  OR cVar2S15S71P028P019P035nsss(0)='1'  )then
          oVar1S632(0) <='1';
          else
          oVar1S632(0) <='0';
          end if;
        if(cVar2S16S71P028P019P010nsss(0)='1'  OR cVar2S17S71N028P013nsss(0)='1'  OR cVar2S18S71N028N013P022nsss(0)='1'  OR cVar2S19S71P034P006P008nsss(0)='1'  )then
          oVar1S633(0) <='1';
          else
          oVar1S633(0) <='0';
          end if;
        if(cVar2S20S71P034N006P019nsss(0)='1'  OR cVar2S21S71P034P027nsss(0)='1'  OR cVar2S22S71P055P004P009nsss(0)='1'  OR cVar2S23S71P034nsss(0)='1'  )then
          oVar1S634(0) <='1';
          else
          oVar1S634(0) <='0';
          end if;
        if(cVar2S24S71N034P012P036nsss(0)='1'  OR cVar2S25S71N034N012P009nsss(0)='1'  OR cVar2S26S71P019P017nsss(0)='1'  OR cVar2S27S71P042P013P011nsss(0)='1'  )then
          oVar1S635(0) <='1';
          else
          oVar1S635(0) <='0';
          end if;
        if(cVar2S28S71P042P013P034nsss(0)='1'  OR cVar2S29S71P009P019P015nsss(0)='1'  OR cVar2S30S71N009P000P036nsss(0)='1'  OR cVar2S31S71P018P019nsss(0)='1'  )then
          oVar1S636(0) <='1';
          else
          oVar1S636(0) <='0';
          end if;
        if(cVar2S32S71P018P047P007nsss(0)='1'  )then
          oVar1S637(0) <='1';
          else
          oVar1S637(0) <='0';
          end if;
        if(cVar2S0S72P006nsss(0)='1'  OR cVar2S1S72P013P021nsss(0)='1'  OR cVar2S2S72N013P006nsss(0)='1'  OR cVar2S3S72N013N006P044nsss(0)='1'  )then
          oVar1S638(0) <='1';
          else
          oVar1S638(0) <='0';
          end if;
        if(cVar2S4S72P054P018nsss(0)='1'  OR cVar2S5S72P054P018P036nsss(0)='1'  OR cVar2S6S72N054P060nsss(0)='1'  OR cVar2S7S72N054N060P053nsss(0)='1'  )then
          oVar1S639(0) <='1';
          else
          oVar1S639(0) <='0';
          end if;
        if(cVar1S8S72P069P045P018P006nsss(0)='1'  OR cVar2S9S72P067nsss(0)='1'  OR cVar2S10S72P015P019nsss(0)='1'  OR cVar2S11S72P006P017nsss(0)='1'  )then
          oVar1S640(0) <='1';
          else
          oVar1S640(0) <='0';
          end if;
        if(cVar2S12S72P006P017P035nsss(0)='1'  OR cVar2S13S72P012P025nsss(0)='1'  OR cVar2S14S72P012P010P009nsss(0)='1'  OR cVar2S15S72P020P050nsss(0)='1'  )then
          oVar1S641(0) <='1';
          else
          oVar1S641(0) <='0';
          end if;
        if(cVar2S16S72N020P016nsss(0)='1'  OR cVar2S17S72N020P016P053nsss(0)='1'  OR cVar2S18S72P031nsss(0)='1'  OR cVar2S19S72N031P053P030nsss(0)='1'  )then
          oVar1S642(0) <='1';
          else
          oVar1S642(0) <='0';
          end if;
        if(cVar2S20S72P059P057P013nsss(0)='1'  OR cVar2S21S72P059N057P010nsss(0)='1'  OR cVar2S22S72P059P033nsss(0)='1'  OR cVar2S23S72P039P044nsss(0)='1'  )then
          oVar1S643(0) <='1';
          else
          oVar1S643(0) <='0';
          end if;
        if(cVar2S24S72P039P003nsss(0)='1'  OR cVar2S25S72P039N003P035nsss(0)='1'  OR cVar2S26S72P016P061nsss(0)='1'  OR cVar2S27S72P016P033P008nsss(0)='1'  )then
          oVar1S644(0) <='1';
          else
          oVar1S644(0) <='0';
          end if;
        if(cVar2S0S73P003nsss(0)='1'  OR cVar2S1S73P065nsss(0)='1'  OR cVar2S2S73N065P068nsss(0)='1'  OR cVar2S3S73N065N068P012nsss(0)='1'  )then
          oVar1S646(0) <='1';
          else
          oVar1S646(0) <='0';
          end if;
        if(cVar2S4S73P018P005nsss(0)='1'  OR cVar2S5S73P018P005P002nsss(0)='1'  OR cVar2S6S73N018P059P000nsss(0)='1'  OR cVar2S7S73N018P059P034nsss(0)='1'  )then
          oVar1S647(0) <='1';
          else
          oVar1S647(0) <='0';
          end if;
        if(cVar2S8S73P011P014nsss(0)='1'  OR cVar2S9S73N011P009nsss(0)='1'  OR cVar2S10S73N011N009P033nsss(0)='1'  OR cVar2S11S73P066nsss(0)='1'  )then
          oVar1S648(0) <='1';
          else
          oVar1S648(0) <='0';
          end if;
        if(cVar2S12S73N066P012nsss(0)='1'  OR cVar2S13S73P009nsss(0)='1'  OR cVar2S14S73N009P067P048nsss(0)='1'  OR cVar2S15S73N009P067P019nsss(0)='1'  )then
          oVar1S649(0) <='1';
          else
          oVar1S649(0) <='0';
          end if;
        if(cVar2S16S73P048nsss(0)='1'  OR cVar2S17S73N048P051nsss(0)='1'  OR cVar2S18S73N048N051P011nsss(0)='1'  OR cVar2S19S73P002nsss(0)='1'  )then
          oVar1S650(0) <='1';
          else
          oVar1S650(0) <='0';
          end if;
        if(cVar2S20S73N002P000nsss(0)='1'  OR cVar2S21S73N002N000P021nsss(0)='1'  OR cVar2S22S73P028P043nsss(0)='1'  OR cVar2S23S73P028N043P030nsss(0)='1'  )then
          oVar1S651(0) <='1';
          else
          oVar1S651(0) <='0';
          end if;
        if(cVar2S24S73N028P067P034nsss(0)='1'  OR cVar2S25S73N028N067P035nsss(0)='1'  OR cVar2S26S73P013P009nsss(0)='1'  OR cVar2S27S73N013P047P049nsss(0)='1'  )then
          oVar1S652(0) <='1';
          else
          oVar1S652(0) <='0';
          end if;
        if(cVar2S28S73P066P064P059nsss(0)='1'  OR cVar2S29S73N066P019P069nsss(0)='1'  OR cVar2S30S73P067nsss(0)='1'  )then
          oVar1S653(0) <='1';
          else
          oVar1S653(0) <='0';
          end if;
        if(cVar2S0S74P049P058nsss(0)='1'  OR cVar2S1S74P049N058P024nsss(0)='1'  OR cVar2S2S74N049P050nsss(0)='1'  OR cVar2S3S74N049N050P048nsss(0)='1'  )then
          oVar1S654(0) <='1';
          else
          oVar1S654(0) <='0';
          end if;
        if(cVar2S4S74P055P015nsss(0)='1'  OR cVar2S5S74P055N015P051nsss(0)='1'  OR cVar2S6S74N055P057P022nsss(0)='1'  OR cVar2S7S74P010nsss(0)='1'  )then
          oVar1S655(0) <='1';
          else
          oVar1S655(0) <='0';
          end if;
        if(cVar2S8S74N010P008nsss(0)='1'  OR cVar2S9S74N010N008P014nsss(0)='1'  OR cVar2S10S74P026P037P013nsss(0)='1'  OR cVar2S11S74P028nsss(0)='1'  )then
          oVar1S656(0) <='1';
          else
          oVar1S656(0) <='0';
          end if;
        if(cVar2S12S74N028P051nsss(0)='1'  OR cVar2S13S74N028N051P055nsss(0)='1'  OR cVar2S14S74P057P011P010nsss(0)='1'  OR cVar2S15S74P057P066P051nsss(0)='1'  )then
          oVar1S657(0) <='1';
          else
          oVar1S657(0) <='0';
          end if;
        if(cVar2S16S74P035nsss(0)='1'  OR cVar1S17S74P016P043P062nsss(0)='1'  OR cVar1S18S74P016P043N062P022nsss(0)='1'  OR cVar2S19S74P006nsss(0)='1'  )then
          oVar1S658(0) <='1';
          else
          oVar1S658(0) <='0';
          end if;
        if(cVar2S20S74N006P068P019nsss(0)='1'  OR cVar2S21S74P010P052nsss(0)='1'  OR cVar2S22S74P010N052P029nsss(0)='1'  OR cVar2S23S74N010P054P014nsss(0)='1'  )then
          oVar1S659(0) <='1';
          else
          oVar1S659(0) <='0';
          end if;
        if(cVar2S24S74P011P026P067nsss(0)='1'  OR cVar2S25S74P011P010P055nsss(0)='1'  OR cVar2S26S74P018P066nsss(0)='1'  OR cVar2S27S74P018N066P017nsss(0)='1'  )then
          oVar1S660(0) <='1';
          else
          oVar1S660(0) <='0';
          end if;
        if(cVar2S0S75P037P048nsss(0)='1'  OR cVar2S1S75P037N048P052nsss(0)='1'  OR cVar2S2S75P045P014nsss(0)='1'  OR cVar2S3S75P045P014P046nsss(0)='1'  )then
          oVar1S662(0) <='1';
          else
          oVar1S662(0) <='0';
          end if;
        if(cVar2S4S75P009nsss(0)='1'  OR cVar2S5S75P056P031P033nsss(0)='1'  OR cVar2S6S75P056N031P004nsss(0)='1'  OR cVar2S7S75P056P032nsss(0)='1'  )then
          oVar1S663(0) <='1';
          else
          oVar1S663(0) <='0';
          end if;
        if(cVar2S8S75P056N032P013nsss(0)='1'  OR cVar2S9S75P011P066nsss(0)='1'  OR cVar2S10S75N011P067P012nsss(0)='1'  OR cVar2S11S75P007P008nsss(0)='1'  )then
          oVar1S664(0) <='1';
          else
          oVar1S664(0) <='0';
          end if;
        if(cVar2S12S75N007P016P045nsss(0)='1'  OR cVar2S13S75P065P037P069nsss(0)='1'  OR cVar2S14S75P065N037P066nsss(0)='1'  OR cVar2S15S75N065P030P019nsss(0)='1'  )then
          oVar1S665(0) <='1';
          else
          oVar1S665(0) <='0';
          end if;
        if(cVar2S16S75N065N030P051nsss(0)='1'  OR cVar2S17S75P012nsss(0)='1'  OR cVar2S18S75P009P033nsss(0)='1'  OR cVar2S19S75N009P014P062nsss(0)='1'  )then
          oVar1S666(0) <='1';
          else
          oVar1S666(0) <='0';
          end if;
        if(cVar2S20S75N009N014P032nsss(0)='1'  OR cVar2S21S75P017P068P063nsss(0)='1'  OR cVar2S22S75P017P068P062nsss(0)='1'  OR cVar2S23S75P017P063nsss(0)='1'  )then
          oVar1S667(0) <='1';
          else
          oVar1S667(0) <='0';
          end if;
        if(cVar2S24S75P017P063P067nsss(0)='1'  OR cVar2S25S75P019P012nsss(0)='1'  OR cVar2S26S75P019N012P016nsss(0)='1'  OR cVar2S27S75P019P015P011nsss(0)='1'  )then
          oVar1S668(0) <='1';
          else
          oVar1S668(0) <='0';
          end if;
        if(cVar2S28S75P035nsss(0)='1'  OR cVar2S29S75N035P067P063nsss(0)='1'  OR cVar2S30S75N035P067P014nsss(0)='1'  OR cVar2S31S75P055P024nsss(0)='1'  )then
          oVar1S669(0) <='1';
          else
          oVar1S669(0) <='0';
          end if;
        if(cVar2S32S75P055P068nsss(0)='1'  OR cVar2S33S75P055N068P056nsss(0)='1'  )then
          oVar1S670(0) <='1';
          else
          oVar1S670(0) <='0';
          end if;
        if(cVar2S0S76P033P065P068nsss(0)='1'  OR cVar2S1S76P033N065P059nsss(0)='1'  OR cVar2S2S76N033P025nsss(0)='1'  OR cVar2S3S76P052P029nsss(0)='1'  )then
          oVar1S671(0) <='1';
          else
          oVar1S671(0) <='0';
          end if;
        if(cVar2S4S76P052N029P015nsss(0)='1'  OR cVar2S5S76N052P029nsss(0)='1'  OR cVar2S6S76P026P018nsss(0)='1'  OR cVar2S7S76P026N018P030nsss(0)='1'  )then
          oVar1S672(0) <='1';
          else
          oVar1S672(0) <='0';
          end if;
        if(cVar2S8S76P010P057nsss(0)='1'  OR cVar2S9S76P037nsss(0)='1'  OR cVar2S10S76P037P035P019nsss(0)='1'  OR cVar2S11S76P037N035P034nsss(0)='1'  )then
          oVar1S673(0) <='1';
          else
          oVar1S673(0) <='0';
          end if;
        if(cVar2S12S76P066P058nsss(0)='1'  OR cVar2S13S76N066P033nsss(0)='1'  OR cVar2S14S76P036P008P035nsss(0)='1'  OR cVar2S15S76P036P066P019nsss(0)='1'  )then
          oVar1S674(0) <='1';
          else
          oVar1S674(0) <='0';
          end if;
        if(cVar2S16S76P001P068nsss(0)='1'  OR cVar2S17S76P001N068P037nsss(0)='1'  OR cVar2S18S76N001P011nsss(0)='1'  OR cVar2S19S76P032P037nsss(0)='1'  )then
          oVar1S675(0) <='1';
          else
          oVar1S675(0) <='0';
          end if;
        if(cVar2S20S76P032P037P017nsss(0)='1'  OR cVar2S21S76N032P052nsss(0)='1'  OR cVar2S22S76P025nsss(0)='1'  OR cVar2S23S76N025P066P019nsss(0)='1'  )then
          oVar1S676(0) <='1';
          else
          oVar1S676(0) <='0';
          end if;
        if(cVar2S24S76P037nsss(0)='1'  OR cVar2S25S76P031P030nsss(0)='1'  OR cVar2S26S76P031N030P008nsss(0)='1'  OR cVar2S27S76P035P053P007nsss(0)='1'  )then
          oVar1S677(0) <='1';
          else
          oVar1S677(0) <='0';
          end if;
        if(cVar2S28S76P035P053P018nsss(0)='1'  OR cVar2S29S76P035P033P004nsss(0)='1'  OR cVar2S30S76P015P011P033nsss(0)='1'  OR cVar2S31S76P015N011P054nsss(0)='1'  )then
          oVar1S678(0) <='1';
          else
          oVar1S678(0) <='0';
          end if;
        if(cVar2S32S76N015P010P056nsss(0)='1'  OR cVar2S33S76N015N010P014nsss(0)='1'  )then
          oVar1S679(0) <='1';
          else
          oVar1S679(0) <='0';
          end if;
        if(cVar2S0S77P064P018nsss(0)='1'  OR cVar2S1S77P064P018P062nsss(0)='1'  OR cVar2S2S77P064P000P044nsss(0)='1'  OR cVar2S3S77P064P000P033nsss(0)='1'  )then
          oVar1S680(0) <='1';
          else
          oVar1S680(0) <='0';
          end if;
        if(cVar2S4S77P051P018nsss(0)='1'  OR cVar2S5S77P051N018P011nsss(0)='1'  OR cVar2S6S77P014P030nsss(0)='1'  OR cVar2S7S77P014P030P062nsss(0)='1'  )then
          oVar1S681(0) <='1';
          else
          oVar1S681(0) <='0';
          end if;
        if(cVar2S8S77N014P011P020nsss(0)='1'  OR cVar2S9S77N014P011P033nsss(0)='1'  OR cVar2S10S77P013P037P019nsss(0)='1'  OR cVar2S11S77P011nsss(0)='1'  )then
          oVar1S682(0) <='1';
          else
          oVar1S682(0) <='0';
          end if;
        if(cVar2S12S77N011P015nsss(0)='1'  OR cVar2S13S77N011N015P010nsss(0)='1'  OR cVar2S14S77P000P047P009nsss(0)='1'  OR cVar2S15S77P015P010P028nsss(0)='1'  )then
          oVar1S683(0) <='1';
          else
          oVar1S683(0) <='0';
          end if;
        if(cVar2S16S77P015N010P011nsss(0)='1'  OR cVar2S17S77N015P001nsss(0)='1'  OR cVar2S18S77N015N001P031nsss(0)='1'  OR cVar2S19S77P069P060P032nsss(0)='1'  )then
          oVar1S684(0) <='1';
          else
          oVar1S684(0) <='0';
          end if;
        if(cVar1S20S77P035P052P012P029nsss(0)='1'  OR cVar2S21S77P060P067nsss(0)='1'  OR cVar2S22S77P060N067P027nsss(0)='1'  OR cVar1S23S77P035P052P012P064nsss(0)='1'  )then
          oVar1S685(0) <='1';
          else
          oVar1S685(0) <='0';
          end if;
        if(cVar2S24S77P019nsss(0)='1'  OR cVar2S25S77P019P016nsss(0)='1'  OR cVar2S26S77P037nsss(0)='1'  OR cVar2S27S77N037P053nsss(0)='1'  )then
          oVar1S686(0) <='1';
          else
          oVar1S686(0) <='0';
          end if;
        if(cVar2S28S77P007P006P064nsss(0)='1'  OR cVar2S29S77P007P006P045nsss(0)='1'  OR cVar2S30S77P007P057P047nsss(0)='1'  )then
          oVar1S687(0) <='1';
          else
          oVar1S687(0) <='0';
          end if;
        if(cVar1S0S78P035P064P052P036nsss(0)='1'  OR cVar2S1S78P015nsss(0)='1'  OR cVar2S2S78N015P029nsss(0)='1'  OR cVar2S3S78N015N029P017nsss(0)='1'  )then
          oVar1S688(0) <='1';
          else
          oVar1S688(0) <='0';
          end if;
        if(cVar2S4S78P034P067nsss(0)='1'  OR cVar2S5S78P034P067P019nsss(0)='1'  OR cVar2S6S78P034P012nsss(0)='1'  OR cVar2S7S78P034N012P013nsss(0)='1'  )then
          oVar1S689(0) <='1';
          else
          oVar1S689(0) <='0';
          end if;
        if(cVar2S8S78P062P020nsss(0)='1'  OR cVar2S9S78P062N020P001nsss(0)='1'  OR cVar2S10S78N062P068nsss(0)='1'  OR cVar2S11S78P013P031nsss(0)='1'  )then
          oVar1S690(0) <='1';
          else
          oVar1S690(0) <='0';
          end if;
        if(cVar2S12S78P013P015P019nsss(0)='1'  OR cVar2S13S78P013P015P063nsss(0)='1'  OR cVar2S14S78P026P009P069nsss(0)='1'  OR cVar2S15S78P026P009P067nsss(0)='1'  )then
          oVar1S691(0) <='1';
          else
          oVar1S691(0) <='0';
          end if;
        if(cVar2S16S78P056P054nsss(0)='1'  OR cVar2S17S78P018P007P049nsss(0)='1'  OR cVar2S18S78P018P063P011nsss(0)='1'  OR cVar2S19S78P017P056P060nsss(0)='1'  )then
          oVar1S692(0) <='1';
          else
          oVar1S692(0) <='0';
          end if;
        if(cVar2S20S78P017N056P006nsss(0)='1'  OR cVar2S21S78N017P065P020nsss(0)='1'  OR cVar2S22S78P051P057P060nsss(0)='1'  OR cVar2S23S78P051N057P040nsss(0)='1'  )then
          oVar1S693(0) <='1';
          else
          oVar1S693(0) <='0';
          end if;
        if(cVar2S24S78P051P026nsss(0)='1'  OR cVar2S25S78P058P008nsss(0)='1'  OR cVar2S26S78P028P011nsss(0)='1'  OR cVar2S27S78P028N011P037nsss(0)='1'  )then
          oVar1S694(0) <='1';
          else
          oVar1S694(0) <='0';
          end if;
        if(cVar2S28S78N028P047P000nsss(0)='1'  OR cVar2S29S78P014P019P059nsss(0)='1'  OR cVar2S30S78P014N019P061nsss(0)='1'  OR cVar2S31S78N014P045P064nsss(0)='1'  )then
          oVar1S695(0) <='1';
          else
          oVar1S695(0) <='0';
          end if;
        if(cVar2S32S78N014N045P057nsss(0)='1'  OR cVar2S33S78P013P065P069nsss(0)='1'  )then
          oVar1S696(0) <='1';
          else
          oVar1S696(0) <='0';
          end if;
        if(cVar1S0S79P064P035P052P053nsss(0)='1'  OR cVar2S1S79P046P019nsss(0)='1'  OR cVar2S2S79N046P057P059nsss(0)='1'  OR cVar2S3S79N046N057psss(0)='1'  )then
          oVar1S697(0) <='1';
          else
          oVar1S697(0) <='0';
          end if;
        if(cVar2S4S79P056nsss(0)='1'  OR cVar2S5S79N056P013P016nsss(0)='1'  OR cVar2S6S79P009nsss(0)='1'  OR cVar2S7S79N009P050nsss(0)='1'  )then
          oVar1S698(0) <='1';
          else
          oVar1S698(0) <='0';
          end if;
        if(cVar2S8S79N009P050P008nsss(0)='1'  OR cVar2S9S79P058P034P017nsss(0)='1'  OR cVar2S10S79P019P026nsss(0)='1'  OR cVar2S11S79P050nsss(0)='1'  )then
          oVar1S699(0) <='1';
          else
          oVar1S699(0) <='0';
          end if;
        if(cVar2S12S79N050P029P044nsss(0)='1'  OR cVar2S13S79P015P003nsss(0)='1'  OR cVar2S14S79P015P003P045nsss(0)='1'  OR cVar2S15S79P015P055P033nsss(0)='1'  )then
          oVar1S700(0) <='1';
          else
          oVar1S700(0) <='0';
          end if;
        if(cVar2S16S79P015N055P058nsss(0)='1'  OR cVar2S17S79P029nsss(0)='1'  OR cVar2S18S79N029P027nsss(0)='1'  OR cVar2S19S79N029N027P028nsss(0)='1'  )then
          oVar1S701(0) <='1';
          else
          oVar1S701(0) <='0';
          end if;
        if(cVar2S20S79P065P069P060nsss(0)='1'  OR cVar2S21S79N065P037P063nsss(0)='1'  OR cVar2S22S79P029P017P010nsss(0)='1'  OR cVar2S23S79P032P059P014nsss(0)='1'  )then
          oVar1S702(0) <='1';
          else
          oVar1S702(0) <='0';
          end if;
        if(cVar2S24S79P032P059P060nsss(0)='1'  OR cVar2S25S79P032P059P063nsss(0)='1'  OR cVar2S26S79P057nsss(0)='1'  OR cVar2S27S79N057P012nsss(0)='1'  )then
          oVar1S703(0) <='1';
          else
          oVar1S703(0) <='0';
          end if;
        if(cVar2S28S79P015P059P068nsss(0)='1'  OR cVar2S29S79P015P063P016nsss(0)='1'  )then
          oVar1S704(0) <='1';
          else
          oVar1S704(0) <='0';
          end if;
        if(cVar2S0S80P032P010nsss(0)='1'  OR cVar2S1S80P032P010P027nsss(0)='1'  OR cVar2S2S80P032P061P014nsss(0)='1'  OR cVar2S3S80P014P031nsss(0)='1'  )then
          oVar1S705(0) <='1';
          else
          oVar1S705(0) <='0';
          end if;
        if(cVar2S4S80P014N031P009nsss(0)='1'  OR cVar2S5S80P014P031P015nsss(0)='1'  OR cVar2S6S80P016nsss(0)='1'  OR cVar2S7S80N016P030nsss(0)='1'  )then
          oVar1S706(0) <='1';
          else
          oVar1S706(0) <='0';
          end if;
        if(cVar2S8S80P012P035nsss(0)='1'  OR cVar2S9S80P044nsss(0)='1'  OR cVar2S10S80N044P011nsss(0)='1'  OR cVar2S11S80N044P011P058nsss(0)='1'  )then
          oVar1S707(0) <='1';
          else
          oVar1S707(0) <='0';
          end if;
        if(cVar2S12S80P031P062nsss(0)='1'  OR cVar2S13S80N031P032P009nsss(0)='1'  OR cVar2S14S80P061P013nsss(0)='1'  OR cVar2S15S80P061P031P058nsss(0)='1'  )then
          oVar1S708(0) <='1';
          else
          oVar1S708(0) <='0';
          end if;
        if(cVar2S16S80P061P031P013nsss(0)='1'  OR cVar2S17S80P032P005nsss(0)='1'  OR cVar2S18S80N032P058P031nsss(0)='1'  OR cVar2S19S80N032P058P016nsss(0)='1'  )then
          oVar1S709(0) <='1';
          else
          oVar1S709(0) <='0';
          end if;
        if(cVar1S20S80P037P015P052P029nsss(0)='1'  OR cVar2S21S80P018P016nsss(0)='1'  OR cVar2S22S80P016P068nsss(0)='1'  OR cVar2S23S80P016N068P018nsss(0)='1'  )then
          oVar1S710(0) <='1';
          else
          oVar1S710(0) <='0';
          end if;
        if(cVar2S24S80P026P047P024nsss(0)='1'  OR cVar2S25S80P026P053P068nsss(0)='1'  OR cVar2S26S80P034P035nsss(0)='1'  OR cVar2S27S80P034P035P017nsss(0)='1'  )then
          oVar1S711(0) <='1';
          else
          oVar1S711(0) <='0';
          end if;
        if(cVar2S28S80N034P062P061nsss(0)='1'  OR cVar2S29S80N034P062P059nsss(0)='1'  OR cVar2S30S80P053P062nsss(0)='1'  OR cVar2S31S80P040P062nsss(0)='1'  )then
          oVar1S712(0) <='1';
          else
          oVar1S712(0) <='0';
          end if;
        if(cVar2S32S80P040N062P038nsss(0)='1'  OR cVar2S33S80N040P055P008nsss(0)='1'  OR cVar2S34S80N040N055P035nsss(0)='1'  OR cVar2S35S80P060P069nsss(0)='1'  )then
          oVar1S713(0) <='1';
          else
          oVar1S713(0) <='0';
          end if;
        if(cVar2S36S80P060N069P019nsss(0)='1'  OR cVar2S37S80N060P030nsss(0)='1'  )then
          oVar1S714(0) <='1';
          else
          oVar1S714(0) <='0';
          end if;
        if(cVar2S0S81P029P030P052nsss(0)='1'  OR cVar2S1S81N029P054nsss(0)='1'  OR cVar2S2S81N029P054P028nsss(0)='1'  OR cVar2S3S81P013P065P028nsss(0)='1'  )then
          oVar1S715(0) <='1';
          else
          oVar1S715(0) <='0';
          end if;
        if(cVar2S4S81N013P052P014nsss(0)='1'  OR cVar2S5S81N013P052P009nsss(0)='1'  OR cVar2S6S81P069P061P018nsss(0)='1'  OR cVar2S7S81N069P062P014nsss(0)='1'  )then
          oVar1S716(0) <='1';
          else
          oVar1S716(0) <='0';
          end if;
        if(cVar2S8S81P069P026P031nsss(0)='1'  OR cVar2S9S81P069P029nsss(0)='1'  OR cVar2S10S81P027P045P014nsss(0)='1'  OR cVar2S11S81P027P045P043nsss(0)='1'  )then
          oVar1S717(0) <='1';
          else
          oVar1S717(0) <='0';
          end if;
        if(cVar2S12S81P010nsss(0)='1'  OR cVar2S13S81N010P019nsss(0)='1'  OR cVar2S14S81P030nsss(0)='1'  OR cVar2S15S81N030P015P036nsss(0)='1'  )then
          oVar1S718(0) <='1';
          else
          oVar1S718(0) <='0';
          end if;
        if(cVar2S16S81N030P015P019nsss(0)='1'  OR cVar2S17S81P012P058nsss(0)='1'  OR cVar2S18S81P012N058P065nsss(0)='1'  OR cVar1S19S81P037P052P008P013nsss(0)='1'  )then
          oVar1S719(0) <='1';
          else
          oVar1S719(0) <='0';
          end if;
        if(cVar2S20S81P027nsss(0)='1'  OR cVar2S21S81N027P017nsss(0)='1'  OR cVar2S22S81N027N017P068nsss(0)='1'  OR cVar2S23S81P017nsss(0)='1'  )then
          oVar1S720(0) <='1';
          else
          oVar1S720(0) <='0';
          end if;
        if(cVar2S24S81N017P067nsss(0)='1'  OR cVar2S25S81N017N067P010nsss(0)='1'  OR cVar2S26S81P033nsss(0)='1'  OR cVar2S27S81N033P065nsss(0)='1'  )then
          oVar1S721(0) <='1';
          else
          oVar1S721(0) <='0';
          end if;
        if(cVar2S28S81N033N065P011nsss(0)='1'  OR cVar1S29S81P037N052P025P044nsss(0)='1'  OR cVar2S30S81P036P016nsss(0)='1'  OR cVar2S31S81N036P062P066nsss(0)='1'  )then
          oVar1S722(0) <='1';
          else
          oVar1S722(0) <='0';
          end if;
        if(cVar2S32S81P021nsss(0)='1'  OR cVar2S33S81N021P066nsss(0)='1'  OR cVar2S34S81N021P066P005nsss(0)='1'  OR cVar2S35S81P047P007P054nsss(0)='1'  )then
          oVar1S723(0) <='1';
          else
          oVar1S723(0) <='0';
          end if;
        if(cVar2S36S81P047P007P022nsss(0)='1'  OR cVar2S37S81P047P026P008nsss(0)='1'  OR cVar2S38S81P047N026P010nsss(0)='1'  )then
          oVar1S724(0) <='1';
          else
          oVar1S724(0) <='0';
          end if;
        if(cVar2S0S82P044P007nsss(0)='1'  OR cVar2S1S82N044P067nsss(0)='1'  OR cVar2S2S82N044P067P063nsss(0)='1'  OR cVar2S3S82P035P036nsss(0)='1'  )then
          oVar1S725(0) <='1';
          else
          oVar1S725(0) <='0';
          end if;
        if(cVar2S4S82P035P007nsss(0)='1'  OR cVar2S5S82P035N007P012nsss(0)='1'  OR cVar2S6S82P012nsss(0)='1'  OR cVar2S7S82P067P029nsss(0)='1'  )then
          oVar1S726(0) <='1';
          else
          oVar1S726(0) <='0';
          end if;
        if(cVar2S8S82P067N029P012nsss(0)='1'  OR cVar2S9S82N067P019P010nsss(0)='1'  OR cVar2S10S82P054nsss(0)='1'  OR cVar2S11S82P018P068nsss(0)='1'  )then
          oVar1S727(0) <='1';
          else
          oVar1S727(0) <='0';
          end if;
        if(cVar2S12S82P018P068P010nsss(0)='1'  OR cVar2S13S82P013P011P057nsss(0)='1'  OR cVar2S14S82P010nsss(0)='1'  OR cVar2S15S82P019P042nsss(0)='1'  )then
          oVar1S728(0) <='1';
          else
          oVar1S728(0) <='0';
          end if;
        if(cVar2S16S82N019P069P036nsss(0)='1'  OR cVar2S17S82N019P069P018nsss(0)='1'  OR cVar2S18S82P005nsss(0)='1'  OR cVar2S19S82N005P014P018nsss(0)='1'  )then
          oVar1S729(0) <='1';
          else
          oVar1S729(0) <='0';
          end if;
        if(cVar2S20S82P067P036nsss(0)='1'  OR cVar2S21S82P067P036nsss(0)='1'  OR cVar2S22S82P056P030nsss(0)='1'  OR cVar2S23S82P056P052P031nsss(0)='1'  )then
          oVar1S730(0) <='1';
          else
          oVar1S730(0) <='0';
          end if;
        if(cVar2S24S82P026nsss(0)='1'  OR cVar2S25S82P000P044P010nsss(0)='1'  )then
          oVar1S731(0) <='1';
          else
          oVar1S731(0) <='0';
          end if;
        if(cVar2S0S83P006P046nsss(0)='1'  OR cVar2S1S83N006P060P049nsss(0)='1'  OR cVar2S2S83N006N060P018nsss(0)='1'  OR cVar2S3S83P024P049nsss(0)='1'  )then
          oVar1S732(0) <='1';
          else
          oVar1S732(0) <='0';
          end if;
        if(cVar2S4S83P024P049P051nsss(0)='1'  OR cVar2S5S83P024P002P020nsss(0)='1'  OR cVar1S6S83P017P037P000P021nsss(0)='1'  OR cVar2S7S83P003P069nsss(0)='1'  )then
          oVar1S733(0) <='1';
          else
          oVar1S733(0) <='0';
          end if;
        if(cVar2S8S83P005nsss(0)='1'  OR cVar2S9S83P029nsss(0)='1'  OR cVar2S10S83N029P067P061nsss(0)='1'  OR cVar2S11S83N029P067P056nsss(0)='1'  )then
          oVar1S734(0) <='1';
          else
          oVar1S734(0) <='0';
          end if;
        if(cVar2S12S83P062P067P000nsss(0)='1'  OR cVar2S13S83P062N067P034nsss(0)='1'  OR cVar2S14S83P062P066P030nsss(0)='1'  OR cVar2S15S83P050nsss(0)='1'  )then
          oVar1S735(0) <='1';
          else
          oVar1S735(0) <='0';
          end if;
        if(cVar2S16S83P015nsss(0)='1'  OR cVar2S17S83P069nsss(0)='1'  OR cVar2S18S83N069P010P012nsss(0)='1'  OR cVar2S19S83P063P005nsss(0)='1'  )then
          oVar1S736(0) <='1';
          else
          oVar1S736(0) <='0';
          end if;
        if(cVar2S20S83P063N005P035nsss(0)='1'  OR cVar2S21S83N063P064P008nsss(0)='1'  OR cVar1S22S83P017N044P023P065nsss(0)='1'  OR cVar2S23S83P005nsss(0)='1'  )then
          oVar1S737(0) <='1';
          else
          oVar1S737(0) <='0';
          end if;
        if(cVar2S0S84P035nsss(0)='1'  OR cVar2S1S84P035P067P068nsss(0)='1'  OR cVar2S2S84P001nsss(0)='1'  OR cVar2S3S84N001P036P062nsss(0)='1'  )then
          oVar1S739(0) <='1';
          else
          oVar1S739(0) <='0';
          end if;
        if(cVar2S4S84N001P036P003nsss(0)='1'  OR cVar2S5S84P014nsss(0)='1'  OR cVar2S6S84P068P036P037nsss(0)='1'  OR cVar2S7S84P068P036P030nsss(0)='1'  )then
          oVar1S740(0) <='1';
          else
          oVar1S740(0) <='0';
          end if;
        if(cVar2S8S84P068P037P011nsss(0)='1'  OR cVar2S9S84P030P057nsss(0)='1'  OR cVar2S10S84P030N057P068nsss(0)='1'  OR cVar2S11S84N030P031nsss(0)='1'  )then
          oVar1S741(0) <='1';
          else
          oVar1S741(0) <='0';
          end if;
        if(cVar2S12S84P065P058nsss(0)='1'  OR cVar2S13S84P065N058P012nsss(0)='1'  OR cVar2S14S84N065P036P017nsss(0)='1'  OR cVar2S15S84N065N036P025nsss(0)='1'  )then
          oVar1S742(0) <='1';
          else
          oVar1S742(0) <='0';
          end if;
        if(cVar2S16S84P067nsss(0)='1'  OR cVar2S17S84P067P037nsss(0)='1'  OR cVar2S18S84P067N037P060nsss(0)='1'  OR cVar2S19S84P059P012nsss(0)='1'  )then
          oVar1S743(0) <='1';
          else
          oVar1S743(0) <='0';
          end if;
        if(cVar2S20S84N059P034P060nsss(0)='1'  OR cVar2S21S84P046P008nsss(0)='1'  OR cVar2S22S84P046P049nsss(0)='1'  OR cVar2S23S84P049P046P051nsss(0)='1'  )then
          oVar1S744(0) <='1';
          else
          oVar1S744(0) <='0';
          end if;
        if(cVar2S24S84N049P046nsss(0)='1'  OR cVar2S25S84N049N046P024nsss(0)='1'  OR cVar2S26S84P069P036nsss(0)='1'  OR cVar2S27S84N069P018P026nsss(0)='1'  )then
          oVar1S745(0) <='1';
          else
          oVar1S745(0) <='0';
          end if;
        if(cVar2S28S84P012P069nsss(0)='1'  OR cVar2S29S84P012P069P068nsss(0)='1'  OR cVar2S30S84P012P018nsss(0)='1'  OR cVar2S31S84P017nsss(0)='1'  )then
          oVar1S746(0) <='1';
          else
          oVar1S746(0) <='0';
          end if;
        if(cVar2S32S84P005P051P050nsss(0)='1'  OR cVar2S33S84P005P039nsss(0)='1'  OR cVar2S34S84P005N039P042nsss(0)='1'  OR cVar2S35S84P059P010nsss(0)='1'  )then
          oVar1S747(0) <='1';
          else
          oVar1S747(0) <='0';
          end if;
        if(cVar2S36S84N059P046P013nsss(0)='1'  OR cVar2S37S84N059N046P041nsss(0)='1'  )then
          oVar1S748(0) <='1';
          else
          oVar1S748(0) <='0';
          end if;
        if(cVar2S0S85P021P058nsss(0)='1'  OR cVar2S1S85P021N058P060nsss(0)='1'  OR cVar2S2S85P021P010P017nsss(0)='1'  OR cVar2S3S85P065P011nsss(0)='1'  )then
          oVar1S749(0) <='1';
          else
          oVar1S749(0) <='0';
          end if;
        if(cVar2S4S85P065N011P016nsss(0)='1'  OR cVar2S5S85N065P012P036nsss(0)='1'  OR cVar2S6S85N065N012P009nsss(0)='1'  OR cVar2S7S85P017P004nsss(0)='1'  )then
          oVar1S750(0) <='1';
          else
          oVar1S750(0) <='0';
          end if;
        if(cVar2S8S85P017P004P065nsss(0)='1'  OR cVar2S9S85N017P069P044nsss(0)='1'  OR cVar2S10S85N017P069P016nsss(0)='1'  OR cVar2S11S85P014P010nsss(0)='1'  )then
          oVar1S751(0) <='1';
          else
          oVar1S751(0) <='0';
          end if;
        if(cVar2S12S85P014N010P060nsss(0)='1'  OR cVar2S13S85N014P061nsss(0)='1'  OR cVar1S14S85P019P051P008P027nsss(0)='1'  OR cVar2S15S85P007P050nsss(0)='1'  )then
          oVar1S752(0) <='1';
          else
          oVar1S752(0) <='0';
          end if;
        if(cVar2S16S85P007P050P026nsss(0)='1'  OR cVar2S17S85P026P069nsss(0)='1'  OR cVar2S18S85N026P006nsss(0)='1'  OR cVar2S19S85N026N006P030nsss(0)='1'  )then
          oVar1S753(0) <='1';
          else
          oVar1S753(0) <='0';
          end if;
        if(cVar2S20S85P030nsss(0)='1'  OR cVar2S21S85P034P036P053nsss(0)='1'  OR cVar2S22S85P034P036P047nsss(0)='1'  OR cVar2S23S85P034P015P068nsss(0)='1'  )then
          oVar1S754(0) <='1';
          else
          oVar1S754(0) <='0';
          end if;
        if(cVar2S24S85P013P063nsss(0)='1'  OR cVar2S25S85P013N063P011nsss(0)='1'  OR cVar2S26S85N013P059nsss(0)='1'  OR cVar2S27S85P013nsss(0)='1'  )then
          oVar1S755(0) <='1';
          else
          oVar1S755(0) <='0';
          end if;
        if(cVar2S28S85P034P069nsss(0)='1'  OR cVar2S29S85P034N069P017nsss(0)='1'  OR cVar2S30S85N034P068P065nsss(0)='1'  OR cVar2S31S85N034N068P035nsss(0)='1'  )then
          oVar1S756(0) <='1';
          else
          oVar1S756(0) <='0';
          end if;
        if(cVar2S32S85P014P065nsss(0)='1'  OR cVar2S33S85P014P068P037nsss(0)='1'  OR cVar2S34S85P002P047nsss(0)='1'  OR cVar2S35S85P002N047P063nsss(0)='1'  )then
          oVar1S757(0) <='1';
          else
          oVar1S757(0) <='0';
          end if;
        if(cVar2S36S85P050nsss(0)='1'  OR cVar2S37S85N050P017P009nsss(0)='1'  OR cVar2S38S85N050N017P047nsss(0)='1'  OR cVar2S39S85P052P058P037nsss(0)='1'  )then
          oVar1S758(0) <='1';
          else
          oVar1S758(0) <='0';
          end if;
        if(cVar2S40S85P052P013P015nsss(0)='1'  OR cVar2S41S85P052N013P026nsss(0)='1'  )then
          oVar1S759(0) <='1';
          else
          oVar1S759(0) <='0';
          end if;
        if(cVar2S0S86P056nsss(0)='1'  OR cVar2S1S86N056P003nsss(0)='1'  OR cVar2S2S86N056N003P008nsss(0)='1'  OR cVar2S3S86P068P013P059nsss(0)='1'  )then
          oVar1S760(0) <='1';
          else
          oVar1S760(0) <='0';
          end if;
        if(cVar2S4S86P068P013P015nsss(0)='1'  OR cVar2S5S86N068P066P015nsss(0)='1'  OR cVar2S6S86P006P005nsss(0)='1'  OR cVar2S7S86P006N005P016nsss(0)='1'  )then
          oVar1S761(0) <='1';
          else
          oVar1S761(0) <='0';
          end if;
        if(cVar2S8S86P006P001nsss(0)='1'  OR cVar2S9S86P006N001P021nsss(0)='1'  OR cVar2S10S86P020nsss(0)='1'  OR cVar2S11S86N020P002nsss(0)='1'  )then
          oVar1S762(0) <='1';
          else
          oVar1S762(0) <='0';
          end if;
        if(cVar2S12S86P037nsss(0)='1'  OR cVar2S13S86P037P013nsss(0)='1'  OR cVar2S14S86P011P066nsss(0)='1'  OR cVar2S15S86N011P061nsss(0)='1'  )then
          oVar1S763(0) <='1';
          else
          oVar1S763(0) <='0';
          end if;
        if(cVar2S16S86N011N061P069nsss(0)='1'  OR cVar2S17S86P033P057P062nsss(0)='1'  OR cVar2S18S86P033P057P059nsss(0)='1'  OR cVar2S19S86P033P013P067nsss(0)='1'  )then
          oVar1S764(0) <='1';
          else
          oVar1S764(0) <='0';
          end if;
        if(cVar2S20S86P025nsss(0)='1'  OR cVar2S21S86P020P005P017nsss(0)='1'  OR cVar2S22S86P020P005P062nsss(0)='1'  OR cVar2S23S86P020P066nsss(0)='1'  )then
          oVar1S765(0) <='1';
          else
          oVar1S765(0) <='0';
          end if;
        if(cVar2S24S86P059P013nsss(0)='1'  OR cVar2S25S86N059P012P056nsss(0)='1'  OR cVar1S26S86N019P067P002P064nsss(0)='1'  OR cVar2S27S86P063P017P018nsss(0)='1'  )then
          oVar1S766(0) <='1';
          else
          oVar1S766(0) <='0';
          end if;
        if(cVar2S28S86P039P059nsss(0)='1'  OR cVar2S29S86P039N059P032nsss(0)='1'  OR cVar2S30S86P029P050nsss(0)='1'  OR cVar2S31S86P029N050P002nsss(0)='1'  )then
          oVar1S767(0) <='1';
          else
          oVar1S767(0) <='0';
          end if;
        if(cVar2S32S86P029P026P035nsss(0)='1'  OR cVar2S33S86P027P050nsss(0)='1'  OR cVar2S34S86P027N050P008nsss(0)='1'  OR cVar2S35S86N027P048P010nsss(0)='1'  )then
          oVar1S768(0) <='1';
          else
          oVar1S768(0) <='0';
          end if;
        if(cVar2S36S86N027P048P025nsss(0)='1'  OR cVar2S37S86P065P036nsss(0)='1'  OR cVar2S38S86P065N036P016nsss(0)='1'  OR cVar2S39S86N065P047nsss(0)='1'  )then
          oVar1S769(0) <='1';
          else
          oVar1S769(0) <='0';
          end if;
        if(cVar2S40S86N065N047P057nsss(0)='1'  )then
          oVar1S770(0) <='1';
          else
          oVar1S770(0) <='0';
          end if;
        if(cVar2S0S87P009P008nsss(0)='1'  OR cVar2S1S87P009P008P016nsss(0)='1'  OR cVar2S2S87N009P069nsss(0)='1'  OR cVar2S3S87N009N069P018nsss(0)='1'  )then
          oVar1S771(0) <='1';
          else
          oVar1S771(0) <='0';
          end if;
        if(cVar2S4S87P009P068P018nsss(0)='1'  OR cVar2S5S87P009P050P012nsss(0)='1'  OR cVar2S6S87P009N050P047nsss(0)='1'  OR cVar1S7S87P017P002P038P004nsss(0)='1'  )then
          oVar1S772(0) <='1';
          else
          oVar1S772(0) <='0';
          end if;
        if(cVar2S8S87N064P009nsss(0)='1'  OR cVar1S9S87P017P002P040nsss(0)='1'  OR cVar2S10S87P036nsss(0)='1'  OR cVar2S11S87N036P019P014nsss(0)='1'  )then
          oVar1S773(0) <='1';
          else
          oVar1S773(0) <='0';
          end if;
        if(cVar2S12S87P035P067nsss(0)='1'  OR cVar2S13S87P035N067P018nsss(0)='1'  OR cVar2S14S87N035P037P019nsss(0)='1'  OR cVar2S15S87P057nsss(0)='1'  )then
          oVar1S774(0) <='1';
          else
          oVar1S774(0) <='0';
          end if;
        if(cVar2S16S87N057P037P053nsss(0)='1'  OR cVar2S17S87N057N037P051nsss(0)='1'  OR cVar2S18S87P042P063nsss(0)='1'  OR cVar2S19S87N042P056P053nsss(0)='1'  )then
          oVar1S775(0) <='1';
          else
          oVar1S775(0) <='0';
          end if;
        if(cVar2S20S87N042N056P010nsss(0)='1'  OR cVar2S21S87P029nsss(0)='1'  OR cVar2S22S87N029P018nsss(0)='1'  OR cVar2S23S87P010P050nsss(0)='1'  )then
          oVar1S776(0) <='1';
          else
          oVar1S776(0) <='0';
          end if;
        if(cVar2S24S87N010P026P008nsss(0)='1'  OR cVar2S25S87N010N026P013nsss(0)='1'  OR cVar2S26S87P018P056nsss(0)='1'  OR cVar2S27S87P018N056P010nsss(0)='1'  )then
          oVar1S777(0) <='1';
          else
          oVar1S777(0) <='0';
          end if;
        if(cVar2S28S87N018P021nsss(0)='1'  OR cVar2S29S87N018N021P014nsss(0)='1'  OR cVar2S30S87P032P059nsss(0)='1'  OR cVar2S31S87N032P047nsss(0)='1'  )then
          oVar1S778(0) <='1';
          else
          oVar1S778(0) <='0';
          end if;
        if(cVar2S32S87N032N047P045nsss(0)='1'  OR cVar2S33S87P018P037P016nsss(0)='1'  OR cVar2S34S87P018P037P015nsss(0)='1'  OR cVar2S35S87P018P036P015nsss(0)='1'  )then
          oVar1S779(0) <='1';
          else
          oVar1S779(0) <='0';
          end if;
        if(cVar2S36S87P018N036P014nsss(0)='1'  OR cVar2S37S87P062P037P024nsss(0)='1'  OR cVar2S38S87P062N037P058nsss(0)='1'  OR cVar2S39S87P062P011nsss(0)='1'  )then
          oVar1S780(0) <='1';
          else
          oVar1S780(0) <='0';
          end if;
        if(cVar2S0S88P019P017nsss(0)='1'  OR cVar2S1S88P019P015nsss(0)='1'  OR cVar2S2S88P019N015P046nsss(0)='1'  OR cVar2S3S88P058P063nsss(0)='1'  )then
          oVar1S782(0) <='1';
          else
          oVar1S782(0) <='0';
          end if;
        if(cVar2S4S88P058N063P064nsss(0)='1'  OR cVar2S5S88N058P054P019nsss(0)='1'  OR cVar2S6S88P003P015nsss(0)='1'  OR cVar2S7S88P003P015P059nsss(0)='1'  )then
          oVar1S783(0) <='1';
          else
          oVar1S783(0) <='0';
          end if;
        if(cVar2S8S88P003P058P019nsss(0)='1'  OR cVar2S9S88P035P069nsss(0)='1'  OR cVar2S10S88P035P069P037nsss(0)='1'  OR cVar2S11S88N035P019P060nsss(0)='1'  )then
          oVar1S784(0) <='1';
          else
          oVar1S784(0) <='0';
          end if;
        if(cVar2S12S88N035N019P058nsss(0)='1'  OR cVar2S13S88P002nsss(0)='1'  OR cVar2S14S88N002P042nsss(0)='1'  OR cVar2S15S88N002N042P017nsss(0)='1'  )then
          oVar1S785(0) <='1';
          else
          oVar1S785(0) <='0';
          end if;
        if(cVar2S16S88P044nsss(0)='1'  OR cVar2S17S88N044P004P064nsss(0)='1'  OR cVar2S18S88P048P033nsss(0)='1'  OR cVar2S19S88P048N033P018nsss(0)='1'  )then
          oVar1S786(0) <='1';
          else
          oVar1S786(0) <='0';
          end if;
        if(cVar2S20S88P048N031P009nsss(0)='1'  OR cVar2S21S88P017P009nsss(0)='1'  OR cVar2S22S88P027nsss(0)='1'  OR cVar2S23S88P011P028P000nsss(0)='1'  )then
          oVar1S787(0) <='1';
          else
          oVar1S787(0) <='0';
          end if;
        if(cVar2S24S88P042nsss(0)='1'  OR cVar2S25S88N042P015P009nsss(0)='1'  OR cVar2S26S88N042N015P017nsss(0)='1'  OR cVar2S27S88P012P017P064nsss(0)='1'  )then
          oVar1S788(0) <='1';
          else
          oVar1S788(0) <='0';
          end if;
        if(cVar2S28S88P012N017P004nsss(0)='1'  OR cVar2S29S88P012P041P059nsss(0)='1'  OR cVar2S30S88P036nsss(0)='1'  OR cVar2S31S88N036P018P011nsss(0)='1'  )then
          oVar1S789(0) <='1';
          else
          oVar1S789(0) <='0';
          end if;
        if(cVar2S32S88P032P061nsss(0)='1'  )then
          oVar1S790(0) <='1';
          else
          oVar1S790(0) <='0';
          end if;
        if(cVar2S0S89P034nsss(0)='1'  OR cVar2S1S89N034P026nsss(0)='1'  OR cVar2S2S89N034P026P018nsss(0)='1'  OR cVar2S3S89P036nsss(0)='1'  )then
          oVar1S791(0) <='1';
          else
          oVar1S791(0) <='0';
          end if;
        if(cVar2S4S89N036P020P009nsss(0)='1'  OR cVar2S5S89N036N020P038nsss(0)='1'  OR cVar2S6S89P064nsss(0)='1'  OR cVar2S7S89N064P066nsss(0)='1'  )then
          oVar1S792(0) <='1';
          else
          oVar1S792(0) <='0';
          end if;
        if(cVar2S8S89N064N066P056nsss(0)='1'  OR cVar2S9S89P064P041nsss(0)='1'  OR cVar2S10S89P064P052nsss(0)='1'  OR cVar2S11S89P046nsss(0)='1'  )then
          oVar1S793(0) <='1';
          else
          oVar1S793(0) <='0';
          end if;
        if(cVar2S12S89N046P033nsss(0)='1'  OR cVar2S13S89N046N033P018nsss(0)='1'  OR cVar2S14S89P029nsss(0)='1'  OR cVar2S15S89N029P046nsss(0)='1'  )then
          oVar1S794(0) <='1';
          else
          oVar1S794(0) <='0';
          end if;
        if(cVar2S16S89N029P046P037nsss(0)='1'  OR cVar2S17S89P023P006nsss(0)='1'  OR cVar2S18S89P023N006P036nsss(0)='1'  OR cVar2S19S89P048P046P004nsss(0)='1'  )then
          oVar1S795(0) <='1';
          else
          oVar1S795(0) <='0';
          end if;
        if(cVar2S20S89P048P062P040nsss(0)='1'  OR cVar2S21S89P027P032nsss(0)='1'  OR cVar2S22S89P027N032P062nsss(0)='1'  OR cVar2S23S89P027P051nsss(0)='1'  )then
          oVar1S796(0) <='1';
          else
          oVar1S796(0) <='0';
          end if;
        if(cVar2S24S89P027N051P048nsss(0)='1'  OR cVar2S25S89P010P019P018nsss(0)='1'  OR cVar2S26S89P036P056nsss(0)='1'  OR cVar2S27S89P036N056P031nsss(0)='1'  )then
          oVar1S797(0) <='1';
          else
          oVar1S797(0) <='0';
          end if;
        if(cVar2S28S89N036P016P019nsss(0)='1'  OR cVar2S29S89N036N016P030nsss(0)='1'  OR cVar2S30S89P036nsss(0)='1'  OR cVar2S31S89N036P018P019nsss(0)='1'  )then
          oVar1S798(0) <='1';
          else
          oVar1S798(0) <='0';
          end if;
        if(cVar2S32S89P060nsss(0)='1'  )then
          oVar1S799(0) <='1';
          else
          oVar1S799(0) <='0';
          end if;
        if(cVar2S0S90P036nsss(0)='1'  OR cVar2S1S90N036P035nsss(0)='1'  OR cVar2S2S90N036N035P015nsss(0)='1'  OR cVar2S3S90P000P034nsss(0)='1'  )then
          oVar1S800(0) <='1';
          else
          oVar1S800(0) <='0';
          end if;
        if(cVar2S4S90P000N034P068nsss(0)='1'  OR cVar2S5S90N000P004nsss(0)='1'  OR cVar2S6S90P023P027nsss(0)='1'  OR cVar2S7S90P023N027P068nsss(0)='1'  )then
          oVar1S801(0) <='1';
          else
          oVar1S801(0) <='0';
          end if;
        if(cVar2S8S90P023nsss(0)='1'  OR cVar2S9S90P069P060P032nsss(0)='1'  OR cVar2S10S90P069N060P037nsss(0)='1'  OR cVar2S11S90P066P019nsss(0)='1'  )then
          oVar1S802(0) <='1';
          else
          oVar1S802(0) <='0';
          end if;
        if(cVar2S12S90P066P019P016nsss(0)='1'  OR cVar2S13S90N066P016P012nsss(0)='1'  OR cVar1S14S90P017P014P047P024nsss(0)='1'  OR cVar2S15S90P046nsss(0)='1'  )then
          oVar1S803(0) <='1';
          else
          oVar1S803(0) <='0';
          end if;
        if(cVar2S16S90P040nsss(0)='1'  OR cVar2S17S90N040P002P044nsss(0)='1'  OR cVar2S18S90N040P002P014nsss(0)='1'  OR cVar2S19S90P066nsss(0)='1'  )then
          oVar1S804(0) <='1';
          else
          oVar1S804(0) <='0';
          end if;
        if(cVar2S20S90P039P066P040nsss(0)='1'  OR cVar2S21S90N039P020P043nsss(0)='1'  OR cVar2S22S90P051P055P018nsss(0)='1'  OR cVar2S23S90N051P042nsss(0)='1'  )then
          oVar1S805(0) <='1';
          else
          oVar1S805(0) <='0';
          end if;
        if(cVar2S24S90P032nsss(0)='1'  OR cVar2S25S90N032P008P015nsss(0)='1'  OR cVar2S26S90P062P066P018nsss(0)='1'  OR cVar2S27S90N062P065P037nsss(0)='1'  )then
          oVar1S806(0) <='1';
          else
          oVar1S806(0) <='0';
          end if;
        if(cVar2S28S90P015P034P065nsss(0)='1'  OR cVar2S29S90N015N057P054nsss(0)='1'  )then
          oVar1S807(0) <='1';
          else
          oVar1S807(0) <='0';
          end if;
        if(cVar2S0S91P025P046nsss(0)='1'  OR cVar2S1S91N025P035nsss(0)='1'  OR cVar2S2S91N025P035P016nsss(0)='1'  OR cVar2S3S91P006P027nsss(0)='1'  )then
          oVar1S808(0) <='1';
          else
          oVar1S808(0) <='0';
          end if;
        if(cVar2S4S91P006N027P047nsss(0)='1'  OR cVar2S5S91N006psss(0)='1'  OR cVar2S6S91P000P020P008nsss(0)='1'  OR cVar2S7S91P015P019nsss(0)='1'  )then
          oVar1S809(0) <='1';
          else
          oVar1S809(0) <='0';
          end if;
        if(cVar2S8S91N015P009P003nsss(0)='1'  OR cVar2S9S91P058nsss(0)='1'  OR cVar2S10S91P058P066P061nsss(0)='1'  OR cVar2S11S91P058N066P018nsss(0)='1'  )then
          oVar1S810(0) <='1';
          else
          oVar1S810(0) <='0';
          end if;
        if(cVar2S12S91P060P069P013nsss(0)='1'  OR cVar2S13S91P060P069P014nsss(0)='1'  OR cVar2S14S91N060P008P037nsss(0)='1'  OR cVar2S15S91N060N008P009nsss(0)='1'  )then
          oVar1S811(0) <='1';
          else
          oVar1S811(0) <='0';
          end if;
        if(cVar2S16S91P062P066P037nsss(0)='1'  OR cVar2S17S91N062P014P018nsss(0)='1'  OR cVar2S18S91P015P034P069nsss(0)='1'  OR cVar2S19S91N015N057P054nsss(0)='1'  )then
          oVar1S812(0) <='1';
          else
          oVar1S812(0) <='0';
          end if;
        if(cVar2S20S91P050nsss(0)='1'  OR cVar2S21S91P015nsss(0)='1'  OR cVar2S22S91P002P038P061nsss(0)='1'  OR cVar2S23S91P002P038P004nsss(0)='1'  )then
          oVar1S813(0) <='1';
          else
          oVar1S813(0) <='0';
          end if;
        if(cVar2S24S91P002P013P036nsss(0)='1'  OR cVar2S25S91P002N013P038nsss(0)='1'  OR cVar2S26S91P004nsss(0)='1'  OR cVar2S27S91N004P019P035nsss(0)='1'  )then
          oVar1S814(0) <='1';
          else
          oVar1S814(0) <='0';
          end if;
        if(cVar1S28S91P017N044P023P065nsss(0)='1'  OR cVar2S29S91P010P022P016nsss(0)='1'  )then
          oVar1S815(0) <='1';
          else
          oVar1S815(0) <='0';
          end if;
        if(cVar2S0S92P002P041nsss(0)='1'  OR cVar2S1S92P002P041P008nsss(0)='1'  OR cVar2S2S92P002P040nsss(0)='1'  OR cVar2S3S92P002N040P064nsss(0)='1'  )then
          oVar1S816(0) <='1';
          else
          oVar1S816(0) <='0';
          end if;
        if(cVar2S4S92P058P066nsss(0)='1'  OR cVar2S5S92P058P066P036nsss(0)='1'  OR cVar2S6S92N058P002P016nsss(0)='1'  OR cVar2S7S92N058N002P052nsss(0)='1'  )then
          oVar1S817(0) <='1';
          else
          oVar1S817(0) <='0';
          end if;
        if(cVar2S8S92P019nsss(0)='1'  OR cVar2S9S92P019P016nsss(0)='1'  OR cVar2S10S92P034P018nsss(0)='1'  OR cVar2S11S92P057nsss(0)='1'  )then
          oVar1S818(0) <='1';
          else
          oVar1S818(0) <='0';
          end if;
        if(cVar2S12S92N057P018nsss(0)='1'  OR cVar2S13S92P019nsss(0)='1'  OR cVar2S14S92P061P058P034nsss(0)='1'  OR cVar2S15S92P061P058P014nsss(0)='1'  )then
          oVar1S819(0) <='1';
          else
          oVar1S819(0) <='0';
          end if;
        if(cVar2S16S92N061P062P019nsss(0)='1'  OR cVar2S17S92N061N062P056nsss(0)='1'  OR cVar2S18S92P061nsss(0)='1'  OR cVar1S19S92N017P006P027P048nsss(0)='1'  )then
          oVar1S820(0) <='1';
          else
          oVar1S820(0) <='0';
          end if;
        if(cVar2S20S92P052nsss(0)='1'  OR cVar2S21S92N052P011nsss(0)='1'  OR cVar2S22S92P063nsss(0)='1'  OR cVar2S23S92P063P037P065nsss(0)='1'  )then
          oVar1S821(0) <='1';
          else
          oVar1S821(0) <='0';
          end if;
        if(cVar2S24S92P054P010P047nsss(0)='1'  OR cVar2S25S92P054P010P043nsss(0)='1'  OR cVar2S26S92P061P013nsss(0)='1'  OR cVar2S27S92P061N013P011nsss(0)='1'  )then
          oVar1S822(0) <='1';
          else
          oVar1S822(0) <='0';
          end if;
        if(cVar2S28S92N061P032nsss(0)='1'  OR cVar2S29S92P053nsss(0)='1'  OR cVar2S30S92N053P013P018nsss(0)='1'  OR cVar2S31S92P021P036P061nsss(0)='1'  )then
          oVar1S823(0) <='1';
          else
          oVar1S823(0) <='0';
          end if;
        if(cVar2S32S92P021N036P061nsss(0)='1'  OR cVar2S33S92P021P012P036nsss(0)='1'  OR cVar2S34S92P041P005nsss(0)='1'  OR cVar2S35S92P041N005P069nsss(0)='1'  )then
          oVar1S824(0) <='1';
          else
          oVar1S824(0) <='0';
          end if;
        if(cVar2S0S93P006P013nsss(0)='1'  OR cVar2S1S93P006N013P068nsss(0)='1'  OR cVar2S2S93N006P054P013nsss(0)='1'  OR cVar2S3S93N006P054P013nsss(0)='1'  )then
          oVar1S826(0) <='1';
          else
          oVar1S826(0) <='0';
          end if;
        if(cVar2S4S93P054P050nsss(0)='1'  OR cVar2S5S93N054P050nsss(0)='1'  OR cVar2S6S93N054N050P028nsss(0)='1'  OR cVar2S7S93P037P051P012nsss(0)='1'  )then
          oVar1S827(0) <='1';
          else
          oVar1S827(0) <='0';
          end if;
        if(cVar2S8S93P037N051P043nsss(0)='1'  OR cVar2S9S93N037P068P061nsss(0)='1'  OR cVar2S10S93N037P068P005nsss(0)='1'  OR cVar2S11S93P013P037P019nsss(0)='1'  )then
          oVar1S828(0) <='1';
          else
          oVar1S828(0) <='0';
          end if;
        if(cVar1S12S93P017P030P061P013nsss(0)='1'  OR cVar2S13S93P016P055nsss(0)='1'  OR cVar2S14S93P016N055P037nsss(0)='1'  OR cVar2S15S93P031P048nsss(0)='1'  )then
          oVar1S829(0) <='1';
          else
          oVar1S829(0) <='0';
          end if;
        if(cVar2S16S93P031P035P069nsss(0)='1'  OR cVar2S17S93P012P014nsss(0)='1'  OR cVar2S18S93P057P031nsss(0)='1'  OR cVar2S19S93P057N031P030nsss(0)='1'  )then
          oVar1S830(0) <='1';
          else
          oVar1S830(0) <='0';
          end if;
        if(cVar2S20S93N057P033P031nsss(0)='1'  OR cVar2S21S93N057N033P032nsss(0)='1'  OR cVar2S22S93P052nsss(0)='1'  OR cVar2S23S93N052P027nsss(0)='1'  )then
          oVar1S831(0) <='1';
          else
          oVar1S831(0) <='0';
          end if;
        if(cVar2S24S93P026P050nsss(0)='1'  OR cVar2S25S93P026N050P045nsss(0)='1'  OR cVar2S26S93P008nsss(0)='1'  OR cVar2S27S93N008P005nsss(0)='1'  )then
          oVar1S832(0) <='1';
          else
          oVar1S832(0) <='0';
          end if;
        if(cVar2S28S93N008N005P007nsss(0)='1'  OR cVar2S29S93P008P035P064nsss(0)='1'  OR cVar2S30S93P008P067P018nsss(0)='1'  OR cVar2S31S93P068P022P015nsss(0)='1'  )then
          oVar1S833(0) <='1';
          else
          oVar1S833(0) <='0';
          end if;
        if(cVar2S32S93P068P022P018nsss(0)='1'  OR cVar2S33S93P040nsss(0)='1'  OR cVar2S34S93N040P037P036nsss(0)='1'  OR cVar2S35S93N040N037P035nsss(0)='1'  )then
          oVar1S834(0) <='1';
          else
          oVar1S834(0) <='0';
          end if;
        if(cVar2S0S94P043P061nsss(0)='1'  OR cVar2S1S94P043N061P010nsss(0)='1'  OR cVar2S2S94P015P068nsss(0)='1'  OR cVar2S3S94P015N068P017nsss(0)='1'  )then
          oVar1S836(0) <='1';
          else
          oVar1S836(0) <='0';
          end if;
        if(cVar2S4S94P065P030nsss(0)='1'  OR cVar2S5S94P065P012nsss(0)='1'  OR cVar2S6S94P037P057P019nsss(0)='1'  OR cVar2S7S94P037N057P066nsss(0)='1'  )then
          oVar1S837(0) <='1';
          else
          oVar1S837(0) <='0';
          end if;
        if(cVar2S8S94N037P053nsss(0)='1'  OR cVar2S9S94P066nsss(0)='1'  OR cVar2S10S94N066P036nsss(0)='1'  OR cVar2S11S94P015P014P018nsss(0)='1'  )then
          oVar1S838(0) <='1';
          else
          oVar1S838(0) <='0';
          end if;
        if(cVar2S12S94P015P014P018nsss(0)='1'  OR cVar2S13S94P015P011nsss(0)='1'  OR cVar2S14S94P014nsss(0)='1'  OR cVar2S15S94P014P058nsss(0)='1'  )then
          oVar1S839(0) <='1';
          else
          oVar1S839(0) <='0';
          end if;
        if(cVar2S16S94N014P067P036nsss(0)='1'  OR cVar2S17S94P008P066nsss(0)='1'  OR cVar2S18S94N008P048P026nsss(0)='1'  OR cVar2S19S94N008P048P050nsss(0)='1'  )then
          oVar1S840(0) <='1';
          else
          oVar1S840(0) <='0';
          end if;
        if(cVar2S20S94P058P066nsss(0)='1'  OR cVar2S21S94P058N066P037nsss(0)='1'  OR cVar2S22S94P058P061P060nsss(0)='1'  OR cVar2S23S94P069nsss(0)='1'  )then
          oVar1S841(0) <='1';
          else
          oVar1S841(0) <='0';
          end if;
        if(cVar2S24S94N069P018nsss(0)='1'  OR cVar2S25S94N069P018P011nsss(0)='1'  OR cVar2S26S94P022P016P042nsss(0)='1'  OR cVar2S27S94P031nsss(0)='1'  )then
          oVar1S842(0) <='1';
          else
          oVar1S842(0) <='0';
          end if;
        if(cVar2S28S94P031P054P018nsss(0)='1'  OR cVar2S29S94P031N054P058nsss(0)='1'  OR cVar2S30S94P034P058nsss(0)='1'  OR cVar2S31S94N034P004P069nsss(0)='1'  )then
          oVar1S843(0) <='1';
          else
          oVar1S843(0) <='0';
          end if;
        if(cVar2S32S94N034N004P005nsss(0)='1'  OR cVar2S33S94P061P000nsss(0)='1'  OR cVar2S34S94P061N000P043nsss(0)='1'  OR cVar2S35S94P061P067P060nsss(0)='1'  )then
          oVar1S844(0) <='1';
          else
          oVar1S844(0) <='0';
          end if;
        if(cVar2S36S94P000P037P011nsss(0)='1'  OR cVar2S37S94P000P033P039nsss(0)='1'  )then
          oVar1S845(0) <='1';
          else
          oVar1S845(0) <='0';
          end if;
        if(cVar2S0S95P025P046nsss(0)='1'  OR cVar2S1S95P025N046P066nsss(0)='1'  OR cVar2S2S95N025P051P053nsss(0)='1'  OR cVar2S3S95N025N051P028nsss(0)='1'  )then
          oVar1S846(0) <='1';
          else
          oVar1S846(0) <='0';
          end if;
        if(cVar2S4S95P057nsss(0)='1'  OR cVar2S5S95N057P019P061nsss(0)='1'  OR cVar2S6S95P002nsss(0)='1'  OR cVar2S7S95N002P033P015nsss(0)='1'  )then
          oVar1S847(0) <='1';
          else
          oVar1S847(0) <='0';
          end if;
        if(cVar2S8S95N002N033P009nsss(0)='1'  OR cVar2S9S95P000P037P019nsss(0)='1'  OR cVar2S10S95P000N037P016nsss(0)='1'  OR cVar2S11S95N000P052P029nsss(0)='1'  )then
          oVar1S848(0) <='1';
          else
          oVar1S848(0) <='0';
          end if;
        if(cVar2S12S95N000N052P045nsss(0)='1'  OR cVar1S13S95P013P032P061P067nsss(0)='1'  OR cVar2S14S95P015P033nsss(0)='1'  OR cVar2S15S95P015N033P014nsss(0)='1'  )then
          oVar1S849(0) <='1';
          else
          oVar1S849(0) <='0';
          end if;
        if(cVar2S16S95P015P011nsss(0)='1'  OR cVar2S17S95P015N011P037nsss(0)='1'  OR cVar2S18S95P015nsss(0)='1'  OR cVar2S19S95P014P058nsss(0)='1'  )then
          oVar1S850(0) <='1';
          else
          oVar1S850(0) <='0';
          end if;
        if(cVar2S20S95P014N058P011nsss(0)='1'  OR cVar2S21S95P022nsss(0)='1'  OR cVar2S22S95N022P020nsss(0)='1'  OR cVar2S23S95P066P040P063nsss(0)='1'  )then
          oVar1S851(0) <='1';
          else
          oVar1S851(0) <='0';
          end if;
        if(cVar2S24S95P066P040P039nsss(0)='1'  OR cVar2S25S95P066P014P068nsss(0)='1'  OR cVar2S26S95P012P010nsss(0)='1'  OR cVar2S27S95N012P023P026nsss(0)='1'  )then
          oVar1S852(0) <='1';
          else
          oVar1S852(0) <='0';
          end if;
        if(cVar2S28S95P033P026nsss(0)='1'  OR cVar2S29S95P033N026P032nsss(0)='1'  OR cVar2S30S95P027P018nsss(0)='1'  OR cVar2S31S95P027P018P014nsss(0)='1'  )then
          oVar1S853(0) <='1';
          else
          oVar1S853(0) <='0';
          end if;
        if(cVar2S32S95N027P002nsss(0)='1'  OR cVar2S33S95N027P002P009nsss(0)='1'  OR cVar2S34S95P000P063nsss(0)='1'  OR cVar2S35S95P049nsss(0)='1'  )then
          oVar1S854(0) <='1';
          else
          oVar1S854(0) <='0';
          end if;
        if(cVar2S36S95N049P010nsss(0)='1'  OR cVar2S37S95N049N010P009nsss(0)='1'  OR cVar2S38S95P001P016nsss(0)='1'  OR cVar2S39S95P001P016P036nsss(0)='1'  )then
          oVar1S855(0) <='1';
          else
          oVar1S855(0) <='0';
          end if;
        if(cVar2S40S95N001P028P055nsss(0)='1'  )then
          oVar1S856(0) <='1';
          else
          oVar1S856(0) <='0';
          end if;
        if(cVar2S0S96P014nsss(0)='1'  OR cVar2S1S96N014P060P056nsss(0)='1'  OR cVar2S2S96N014P060P068nsss(0)='1'  OR cVar2S3S96P022P015nsss(0)='1'  )then
          oVar1S857(0) <='1';
          else
          oVar1S857(0) <='0';
          end if;
        if(cVar2S4S96P022N015P016nsss(0)='1'  OR cVar2S5S96N022P049P015nsss(0)='1'  OR cVar2S6S96N022N049P029nsss(0)='1'  OR cVar2S7S96P018P061nsss(0)='1'  )then
          oVar1S858(0) <='1';
          else
          oVar1S858(0) <='0';
          end if;
        if(cVar2S8S96P018N061P014nsss(0)='1'  OR cVar2S9S96N018P030nsss(0)='1'  OR cVar2S10S96N018N030P033nsss(0)='1'  OR cVar2S11S96P035P004nsss(0)='1'  )then
          oVar1S859(0) <='1';
          else
          oVar1S859(0) <='0';
          end if;
        if(cVar2S12S96P035P017P064nsss(0)='1'  OR cVar2S13S96P062P017nsss(0)='1'  OR cVar2S14S96P062N017P014nsss(0)='1'  OR cVar2S15S96P062P063P014nsss(0)='1'  )then
          oVar1S860(0) <='1';
          else
          oVar1S860(0) <='0';
          end if;
        if(cVar2S16S96P007P031P060nsss(0)='1'  OR cVar2S17S96P007P047nsss(0)='1'  OR cVar2S18S96P007N047P050nsss(0)='1'  OR cVar1S19S96P019P003P057P015nsss(0)='1'  )then
          oVar1S861(0) <='1';
          else
          oVar1S861(0) <='0';
          end if;
        if(cVar2S20S96P018nsss(0)='1'  OR cVar2S21S96P059nsss(0)='1'  OR cVar2S22S96N059P032nsss(0)='1'  OR cVar2S23S96P067P014P069nsss(0)='1'  )then
          oVar1S862(0) <='1';
          else
          oVar1S862(0) <='0';
          end if;
        if(cVar2S24S96P067N014P017nsss(0)='1'  OR cVar2S25S96N067P009P017nsss(0)='1'  OR cVar2S26S96P050P013P014nsss(0)='1'  OR cVar2S27S96P050N013P010nsss(0)='1'  )then
          oVar1S863(0) <='1';
          else
          oVar1S863(0) <='0';
          end if;
        if(cVar2S28S96P010P048P018nsss(0)='1'  OR cVar2S29S96P010N048P066nsss(0)='1'  OR cVar2S30S96N010P047P002nsss(0)='1'  OR cVar2S31S96N010P047P024nsss(0)='1'  )then
          oVar1S864(0) <='1';
          else
          oVar1S864(0) <='0';
          end if;
        if(cVar2S32S96P036P054P007nsss(0)='1'  OR cVar2S33S96P036P054P017nsss(0)='1'  OR cVar2S34S96P036P011nsss(0)='1'  OR cVar2S35S96P065nsss(0)='1'  )then
          oVar1S865(0) <='1';
          else
          oVar1S865(0) <='0';
          end if;
        if(cVar2S36S96N065P030P015nsss(0)='1'  )then
          oVar1S866(0) <='1';
          else
          oVar1S866(0) <='0';
          end if;
        if(cVar2S0S97P008nsss(0)='1'  OR cVar2S1S97P008P011nsss(0)='1'  OR cVar2S2S97P013P035nsss(0)='1'  OR cVar2S3S97P013P035P014nsss(0)='1'  )then
          oVar1S867(0) <='1';
          else
          oVar1S867(0) <='0';
          end if;
        if(cVar2S4S97N013psss(0)='1'  OR cVar2S5S97P055P058P020nsss(0)='1'  OR cVar2S6S97P055N058psss(0)='1'  OR cVar2S7S97P055P063nsss(0)='1'  )then
          oVar1S868(0) <='1';
          else
          oVar1S868(0) <='0';
          end if;
        if(cVar2S8S97P021nsss(0)='1'  OR cVar1S9S97P019P057P003P015nsss(0)='1'  OR cVar2S10S97P013nsss(0)='1'  OR cVar2S11S97P013P055nsss(0)='1'  )then
          oVar1S869(0) <='1';
          else
          oVar1S869(0) <='0';
          end if;
        if(cVar2S12S97P013P062nsss(0)='1'  OR cVar2S13S97P066P036nsss(0)='1'  OR cVar2S14S97P066P013P014nsss(0)='1'  OR cVar2S15S97P066N013P063nsss(0)='1'  )then
          oVar1S870(0) <='1';
          else
          oVar1S870(0) <='0';
          end if;
        if(cVar2S16S97P028P010P033nsss(0)='1'  OR cVar2S17S97P028N010psss(0)='1'  OR cVar2S18S97P028P062nsss(0)='1'  OR cVar2S19S97P064P033P035nsss(0)='1'  )then
          oVar1S871(0) <='1';
          else
          oVar1S871(0) <='0';
          end if;
        if(cVar2S20S97P064P033P012nsss(0)='1'  OR cVar1S21S97N019P060P021P033nsss(0)='1'  OR cVar2S22S97P038P064nsss(0)='1'  OR cVar2S23S97P038N064P018nsss(0)='1'  )then
          oVar1S872(0) <='1';
          else
          oVar1S872(0) <='0';
          end if;
        if(cVar2S24S97P056P065P001nsss(0)='1'  OR cVar2S25S97P056P065P029nsss(0)='1'  OR cVar2S26S97N056P021nsss(0)='1'  OR cVar2S27S97P017P064P034nsss(0)='1'  )then
          oVar1S873(0) <='1';
          else
          oVar1S873(0) <='0';
          end if;
        if(cVar2S28S97P017P064P015nsss(0)='1'  OR cVar2S29S97P017P057nsss(0)='1'  OR cVar2S30S97P017N057P035nsss(0)='1'  OR cVar2S31S97P037P018nsss(0)='1'  )then
          oVar1S874(0) <='1';
          else
          oVar1S874(0) <='0';
          end if;
        if(cVar2S0S98P018P065nsss(0)='1'  OR cVar2S1S98P018N065P063nsss(0)='1'  OR cVar2S2S98N018P059nsss(0)='1'  OR cVar2S3S98N018N059P055nsss(0)='1'  )then
          oVar1S876(0) <='1';
          else
          oVar1S876(0) <='0';
          end if;
        if(cVar2S4S98P066P069P015nsss(0)='1'  OR cVar2S5S98P051P048nsss(0)='1'  OR cVar2S6S98N051psss(0)='1'  OR cVar2S7S98P030P055nsss(0)='1'  )then
          oVar1S877(0) <='1';
          else
          oVar1S877(0) <='0';
          end if;
        if(cVar2S8S98N030P034P017nsss(0)='1'  OR cVar2S9S98P014P037nsss(0)='1'  OR cVar2S10S98N014P054P033nsss(0)='1'  OR cVar2S11S98N014N054P032nsss(0)='1'  )then
          oVar1S878(0) <='1';
          else
          oVar1S878(0) <='0';
          end if;
        if(cVar2S12S98P033P012nsss(0)='1'  OR cVar2S13S98P033N012P066nsss(0)='1'  OR cVar1S14S98P019P060P021P033nsss(0)='1'  OR cVar2S15S98P058nsss(0)='1'  )then
          oVar1S879(0) <='1';
          else
          oVar1S879(0) <='0';
          end if;
        if(cVar2S16S98N058P006P010nsss(0)='1'  OR cVar2S17S98P014P034nsss(0)='1'  OR cVar2S18S98N014P003P037nsss(0)='1'  OR cVar1S19S98P019P069N013P022nsss(0)='1'  )then
          oVar1S880(0) <='1';
          else
          oVar1S880(0) <='0';
          end if;
        if(cVar2S20S98P007P064nsss(0)='1'  OR cVar2S21S98P007N064P015nsss(0)='1'  OR cVar2S22S98N007P043nsss(0)='1'  OR cVar2S23S98P062nsss(0)='1'  )then
          oVar1S881(0) <='1';
          else
          oVar1S881(0) <='0';
          end if;
        if(cVar2S24S98N062P061nsss(0)='1'  OR cVar2S25S98P007P037P033nsss(0)='1'  OR cVar2S26S98P007P035nsss(0)='1'  OR cVar2S27S98P054P057P013nsss(0)='1'  )then
          oVar1S882(0) <='1';
          else
          oVar1S882(0) <='0';
          end if;
        if(cVar2S28S98P054P057P017nsss(0)='1'  OR cVar2S29S98N054P031P057nsss(0)='1'  OR cVar2S30S98P026P066P061nsss(0)='1'  )then
          oVar1S883(0) <='1';
          else
          oVar1S883(0) <='0';
          end if;
        if(cVar1S0S99P019P069P006P027nsss(0)='1'  OR cVar2S1S99P044nsss(0)='1'  OR cVar2S2S99N044P047nsss(0)='1'  OR cVar2S3S99N044N047P008nsss(0)='1'  )then
          oVar1S884(0) <='1';
          else
          oVar1S884(0) <='0';
          end if;
        if(cVar2S4S99P025P066nsss(0)='1'  OR cVar2S5S99P025N066P018nsss(0)='1'  OR cVar2S6S99N025P008nsss(0)='1'  OR cVar2S7S99P049P026nsss(0)='1'  )then
          oVar1S885(0) <='1';
          else
          oVar1S885(0) <='0';
          end if;
        if(cVar2S8S99P062P057nsss(0)='1'  OR cVar2S9S99P062N057P018nsss(0)='1'  OR cVar2S10S99N062P034P056nsss(0)='1'  OR cVar2S11S99N062P034P020nsss(0)='1'  )then
          oVar1S886(0) <='1';
          else
          oVar1S886(0) <='0';
          end if;
        if(cVar2S12S99P001P011P005nsss(0)='1'  OR cVar2S13S99P001P011P014nsss(0)='1'  OR cVar2S14S99N001P059nsss(0)='1'  OR cVar2S15S99N001N059P033nsss(0)='1'  )then
          oVar1S887(0) <='1';
          else
          oVar1S887(0) <='0';
          end if;
        if(cVar2S16S99P020P002P063nsss(0)='1'  OR cVar2S17S99P026P062P066nsss(0)='1'  OR cVar2S18S99P026N062P065nsss(0)='1'  OR cVar2S19S99P020P060nsss(0)='1'  )then
          oVar1S888(0) <='1';
          else
          oVar1S888(0) <='0';
          end if;
        if(cVar2S20S99P020P060P059nsss(0)='1'  OR cVar2S21S99P020P037nsss(0)='1'  OR cVar2S22S99P069P012P017nsss(0)='1'  OR cVar2S23S99P013nsss(0)='1'  )then
          oVar1S889(0) <='1';
          else
          oVar1S889(0) <='0';
          end if;
        if(cVar2S24S99N013P010nsss(0)='1'  OR cVar2S25S99N013N010P011nsss(0)='1'  OR cVar2S26S99P037nsss(0)='1'  OR cVar2S27S99P025P057P009nsss(0)='1'  )then
          oVar1S890(0) <='1';
          else
          oVar1S890(0) <='0';
          end if;
        if(cVar2S28S99P025N057P031nsss(0)='1'  OR cVar2S29S99P025P046nsss(0)='1'  OR cVar2S30S99P025P004P046nsss(0)='1'  OR cVar2S31S99P025N004P028nsss(0)='1'  )then
          oVar1S891(0) <='1';
          else
          oVar1S891(0) <='0';
          end if;
        if(cVar2S32S99N025P012P007nsss(0)='1'  OR cVar2S33S99P057P017P005nsss(0)='1'  OR cVar2S34S99P057P030P015nsss(0)='1'  OR cVar2S35S99P015P018nsss(0)='1'  )then
          oVar1S892(0) <='1';
          else
          oVar1S892(0) <='0';
          end if;
        if(cVar2S36S99N015P067P063nsss(0)='1'  )then
          oVar1S893(0) <='1';
          else
          oVar1S893(0) <='0';
          end if;
        if(cVar2S0S100P064P005P013nsss(0)='1'  OR cVar2S1S100P064P005P058nsss(0)='1'  OR cVar2S2S100P064P068P061nsss(0)='1'  OR cVar2S3S100P044P035nsss(0)='1'  )then
          oVar1S894(0) <='1';
          else
          oVar1S894(0) <='0';
          end if;
        if(cVar2S4S100P044N035P032nsss(0)='1'  OR cVar2S5S100N044P038P039nsss(0)='1'  OR cVar2S6S100N044N038psss(0)='1'  OR cVar2S7S100P029P037nsss(0)='1'  )then
          oVar1S895(0) <='1';
          else
          oVar1S895(0) <='0';
          end if;
        if(cVar2S8S100P029N037P034nsss(0)='1'  OR cVar2S9S100N029P034P003nsss(0)='1'  OR cVar2S10S100N029P034P068nsss(0)='1'  OR cVar2S11S100P064P060nsss(0)='1'  )then
          oVar1S896(0) <='1';
          else
          oVar1S896(0) <='0';
          end if;
        if(cVar2S12S100P064P060P014nsss(0)='1'  OR cVar2S13S100P064P037P069nsss(0)='1'  OR cVar2S14S100P061P017nsss(0)='1'  OR cVar2S15S100P061P017P015nsss(0)='1'  )then
          oVar1S897(0) <='1';
          else
          oVar1S897(0) <='0';
          end if;
        if(cVar2S16S100N061P065P017nsss(0)='1'  OR cVar2S17S100N061N065P001nsss(0)='1'  OR cVar2S18S100P052P050nsss(0)='1'  OR cVar2S19S100P052P050P015nsss(0)='1'  )then
          oVar1S898(0) <='1';
          else
          oVar1S898(0) <='0';
          end if;
        if(cVar2S20S100N052P055nsss(0)='1'  OR cVar2S21S100P058P001nsss(0)='1'  OR cVar2S22S100P058N001P006nsss(0)='1'  OR cVar2S23S100N058P057P015nsss(0)='1'  )then
          oVar1S899(0) <='1';
          else
          oVar1S899(0) <='0';
          end if;
        if(cVar2S24S100P062P013P015nsss(0)='1'  OR cVar2S25S100P027nsss(0)='1'  OR cVar2S26S100N027P037nsss(0)='1'  OR cVar2S27S100N027N037P057nsss(0)='1'  )then
          oVar1S900(0) <='1';
          else
          oVar1S900(0) <='0';
          end if;
        if(cVar2S28S100P017P037nsss(0)='1'  OR cVar2S29S100P012nsss(0)='1'  OR cVar2S30S100P052P029nsss(0)='1'  OR cVar2S31S100P052N029P019nsss(0)='1'  )then
          oVar1S901(0) <='1';
          else
          oVar1S901(0) <='0';
          end if;
        if(cVar2S32S100N052P029P000nsss(0)='1'  OR cVar2S33S100P023P005P011nsss(0)='1'  OR cVar2S34S100P023P005P069nsss(0)='1'  OR cVar2S35S100P023P042P069nsss(0)='1'  )then
          oVar1S902(0) <='1';
          else
          oVar1S902(0) <='0';
          end if;
        if(cVar2S36S100P012P064nsss(0)='1'  )then
          oVar1S903(0) <='1';
          else
          oVar1S903(0) <='0';
          end if;
        if(cVar2S0S101P000P069nsss(0)='1'  OR cVar2S1S101P000N069P018nsss(0)='1'  OR cVar2S2S101N000P057nsss(0)='1'  OR cVar2S3S101N000P057P058nsss(0)='1'  )then
          oVar1S904(0) <='1';
          else
          oVar1S904(0) <='0';
          end if;
        if(cVar2S4S101P027P060nsss(0)='1'  OR cVar2S5S101P027N060P067nsss(0)='1'  OR cVar1S6S101P036P005P023P004nsss(0)='1'  OR cVar2S7S101P065nsss(0)='1'  )then
          oVar1S905(0) <='1';
          else
          oVar1S905(0) <='0';
          end if;
        if(cVar2S8S101P033P003nsss(0)='1'  OR cVar2S9S101P033N003P066nsss(0)='1'  OR cVar1S10S101P036P005N069P032nsss(0)='1'  OR cVar2S11S101P058P010P017nsss(0)='1'  )then
          oVar1S906(0) <='1';
          else
          oVar1S906(0) <='0';
          end if;
        if(cVar2S12S101P015nsss(0)='1'  OR cVar2S13S101N015P017nsss(0)='1'  OR cVar2S14S101N015N017P058nsss(0)='1'  OR cVar2S15S101P029P062P026nsss(0)='1'  )then
          oVar1S907(0) <='1';
          else
          oVar1S907(0) <='0';
          end if;
        if(cVar2S16S101P029P062P016nsss(0)='1'  OR cVar2S17S101P029P054P011nsss(0)='1'  OR cVar2S18S101P062P033P066nsss(0)='1'  OR cVar2S19S101P062N033P068nsss(0)='1'  )then
          oVar1S908(0) <='1';
          else
          oVar1S908(0) <='0';
          end if;
        if(cVar2S20S101N062P043nsss(0)='1'  OR cVar2S21S101P021P006P037nsss(0)='1'  OR cVar2S22S101P021N006P057nsss(0)='1'  OR cVar2S23S101P018P064P015nsss(0)='1'  )then
          oVar1S909(0) <='1';
          else
          oVar1S909(0) <='0';
          end if;
        if(cVar2S24S101P018N064P069nsss(0)='1'  OR cVar2S25S101N018P033nsss(0)='1'  OR cVar2S26S101N018N033P011nsss(0)='1'  OR cVar2S27S101P010P016nsss(0)='1'  )then
          oVar1S910(0) <='1';
          else
          oVar1S910(0) <='0';
          end if;
        if(cVar2S28S101P058P016nsss(0)='1'  OR cVar2S29S101P058N016P031nsss(0)='1'  OR cVar2S30S101P058P061P016nsss(0)='1'  OR cVar2S31S101P044nsss(0)='1'  )then
          oVar1S911(0) <='1';
          else
          oVar1S911(0) <='0';
          end if;
        if(cVar2S0S102P059nsss(0)='1'  OR cVar2S1S102N059P065P033nsss(0)='1'  OR cVar2S2S102N059P065P054nsss(0)='1'  OR cVar2S3S102P009P068P015nsss(0)='1'  )then
          oVar1S913(0) <='1';
          else
          oVar1S913(0) <='0';
          end if;
        if(cVar2S4S102P055P056P035nsss(0)='1'  OR cVar2S5S102P055P056P010nsss(0)='1'  OR cVar2S6S102N055P013P003nsss(0)='1'  OR cVar2S7S102N055N013P045nsss(0)='1'  )then
          oVar1S914(0) <='1';
          else
          oVar1S914(0) <='0';
          end if;
        if(cVar2S8S102P011P013P055nsss(0)='1'  OR cVar2S9S102P011P013P012nsss(0)='1'  OR cVar2S10S102P011P003P017nsss(0)='1'  OR cVar2S11S102P017P063nsss(0)='1'  )then
          oVar1S915(0) <='1';
          else
          oVar1S915(0) <='0';
          end if;
        if(cVar2S12S102P017N063P069nsss(0)='1'  OR cVar2S13S102N017P069nsss(0)='1'  OR cVar2S14S102N017P069P033nsss(0)='1'  OR cVar2S15S102P030P057nsss(0)='1'  )then
          oVar1S916(0) <='1';
          else
          oVar1S916(0) <='0';
          end if;
        if(cVar2S16S102P030N057P013nsss(0)='1'  OR cVar2S17S102N030P056P015nsss(0)='1'  OR cVar2S18S102P056P012nsss(0)='1'  OR cVar2S19S102P056N012P013nsss(0)='1'  )then
          oVar1S917(0) <='1';
          else
          oVar1S917(0) <='0';
          end if;
        if(cVar2S20S102N056P044P013nsss(0)='1'  OR cVar1S21S102P036P000P069P009nsss(0)='1'  OR cVar2S22S102P062nsss(0)='1'  OR cVar2S23S102N062P018P015nsss(0)='1'  )then
          oVar1S918(0) <='1';
          else
          oVar1S918(0) <='0';
          end if;
        if(cVar2S24S102P034P032nsss(0)='1'  OR cVar2S25S102P065nsss(0)='1'  OR cVar2S26S102N065P057nsss(0)='1'  OR cVar2S27S102P008P026nsss(0)='1'  )then
          oVar1S919(0) <='1';
          else
          oVar1S919(0) <='0';
          end if;
        if(cVar2S28S102P008N026P031nsss(0)='1'  OR cVar2S29S102N008P011P009nsss(0)='1'  OR cVar2S30S102P058P018nsss(0)='1'  OR cVar2S31S102N058P031P067nsss(0)='1'  )then
          oVar1S920(0) <='1';
          else
          oVar1S920(0) <='0';
          end if;
        if(cVar2S0S103P017P012nsss(0)='1'  OR cVar2S1S103P017P019nsss(0)='1'  OR cVar2S2S103P045P038nsss(0)='1'  OR cVar2S3S103P045P038P019nsss(0)='1'  )then
          oVar1S922(0) <='1';
          else
          oVar1S922(0) <='0';
          end if;
        if(cVar2S4S103P045P016P018nsss(0)='1'  OR cVar2S5S103P069nsss(0)='1'  OR cVar1S6S103P036P001P034P037nsss(0)='1'  OR cVar1S7S103P036P001N034P033nsss(0)='1'  )then
          oVar1S923(0) <='1';
          else
          oVar1S923(0) <='0';
          end if;
        if(cVar2S8S103P068P037P067nsss(0)='1'  OR cVar2S9S103P007P050nsss(0)='1'  OR cVar2S10S103P007N050P052nsss(0)='1'  OR cVar2S11S103P007P018P068nsss(0)='1'  )then
          oVar1S924(0) <='1';
          else
          oVar1S924(0) <='0';
          end if;
        if(cVar2S12S103P007N018P062nsss(0)='1'  OR cVar2S13S103P052P019nsss(0)='1'  OR cVar2S14S103N052P063P015nsss(0)='1'  OR cVar1S15S103N036P011P040P038nsss(0)='1'  )then
          oVar1S925(0) <='1';
          else
          oVar1S925(0) <='0';
          end if;
        if(cVar2S16S103P010nsss(0)='1'  OR cVar2S17S103P012P013nsss(0)='1'  OR cVar2S18S103P012P013P017nsss(0)='1'  OR cVar2S19S103N012P017nsss(0)='1'  )then
          oVar1S926(0) <='1';
          else
          oVar1S926(0) <='0';
          end if;
        if(cVar2S20S103N012N017P013nsss(0)='1'  OR cVar2S21S103P010P018P017nsss(0)='1'  OR cVar2S22S103P010P018P033nsss(0)='1'  OR cVar2S23S103P067P032nsss(0)='1'  )then
          oVar1S927(0) <='1';
          else
          oVar1S927(0) <='0';
          end if;
        if(cVar2S24S103P067P032P035nsss(0)='1'  OR cVar2S25S103P067P059nsss(0)='1'  OR cVar2S26S103P067N059P048nsss(0)='1'  OR cVar2S27S103P031P007P049nsss(0)='1'  )then
          oVar1S928(0) <='1';
          else
          oVar1S928(0) <='0';
          end if;
        if(cVar2S28S103P031N007P001nsss(0)='1'  OR cVar2S29S103P031P010P067nsss(0)='1'  )then
          oVar1S929(0) <='1';
          else
          oVar1S929(0) <='0';
          end if;
        if(cVar2S0S104P009nsss(0)='1'  OR cVar2S1S104N009P050nsss(0)='1'  OR cVar2S2S104P013nsss(0)='1'  OR cVar2S3S104N013P034nsss(0)='1'  )then
          oVar1S930(0) <='1';
          else
          oVar1S930(0) <='0';
          end if;
        if(cVar2S4S104N013N034P059nsss(0)='1'  OR cVar2S5S104P057P031P027nsss(0)='1'  OR cVar2S6S104P049P026P013nsss(0)='1'  OR cVar2S7S104P049P026P050nsss(0)='1'  )then
          oVar1S931(0) <='1';
          else
          oVar1S931(0) <='0';
          end if;
        if(cVar2S8S104P049P007P046nsss(0)='1'  OR cVar2S9S104P049N007P005nsss(0)='1'  OR cVar2S10S104P047nsss(0)='1'  OR cVar2S11S104N047P050nsss(0)='1'  )then
          oVar1S932(0) <='1';
          else
          oVar1S932(0) <='0';
          end if;
        if(cVar2S12S104P057P018nsss(0)='1'  OR cVar2S13S104P057P018P012nsss(0)='1'  OR cVar2S14S104P057P019P013nsss(0)='1'  OR cVar1S15S104P036P043P022nsss(0)='1'  )then
          oVar1S933(0) <='1';
          else
          oVar1S933(0) <='0';
          end if;
        if(cVar1S16S104P036P043N022P024nsss(0)='1'  OR cVar2S17S104P062nsss(0)='1'  OR cVar2S18S104N062P016P069nsss(0)='1'  OR cVar2S19S104P005P003P049nsss(0)='1'  )then
          oVar1S934(0) <='1';
          else
          oVar1S934(0) <='0';
          end if;
        if(cVar2S20S104P005P031P069nsss(0)='1'  OR cVar2S21S104P040P019nsss(0)='1'  OR cVar2S22S104P037nsss(0)='1'  OR cVar2S23S104P066P012P067nsss(0)='1'  )then
          oVar1S935(0) <='1';
          else
          oVar1S935(0) <='0';
          end if;
        if(cVar2S0S105P033nsss(0)='1'  OR cVar2S1S105P055nsss(0)='1'  OR cVar2S2S105P055P031nsss(0)='1'  OR cVar2S3S105P014nsss(0)='1'  )then
          oVar1S937(0) <='1';
          else
          oVar1S937(0) <='0';
          end if;
        if(cVar2S4S105P031nsss(0)='1'  OR cVar2S5S105N031P032P068nsss(0)='1'  OR cVar2S6S105N031N032P062nsss(0)='1'  OR cVar2S7S105P028P018nsss(0)='1'  )then
          oVar1S938(0) <='1';
          else
          oVar1S938(0) <='0';
          end if;
        if(cVar2S8S105P028P018P019nsss(0)='1'  OR cVar2S9S105N028P026P053nsss(0)='1'  OR cVar2S10S105N028N026P029nsss(0)='1'  OR cVar2S11S105P028P057nsss(0)='1'  )then
          oVar1S939(0) <='1';
          else
          oVar1S939(0) <='0';
          end if;
        if(cVar2S12S105P028N057P025nsss(0)='1'  OR cVar2S13S105P028P030P016nsss(0)='1'  OR cVar2S14S105P018nsss(0)='1'  OR cVar2S15S105P014P058nsss(0)='1'  )then
          oVar1S940(0) <='1';
          else
          oVar1S940(0) <='0';
          end if;
        if(cVar2S16S105P051P038nsss(0)='1'  OR cVar2S17S105P051P008nsss(0)='1'  OR cVar2S18S105P003P017nsss(0)='1'  OR cVar2S19S105P003N017P051nsss(0)='1'  )then
          oVar1S941(0) <='1';
          else
          oVar1S941(0) <='0';
          end if;
        if(cVar2S20S105P003P005nsss(0)='1'  OR cVar2S21S105P003N005P034nsss(0)='1'  OR cVar2S22S105P004P034nsss(0)='1'  OR cVar2S23S105P067nsss(0)='1'  )then
          oVar1S942(0) <='1';
          else
          oVar1S942(0) <='0';
          end if;
        if(cVar2S24S105N067P035nsss(0)='1'  OR cVar2S25S105P050P029nsss(0)='1'  OR cVar2S26S105N050P022nsss(0)='1'  OR cVar2S27S105P021P042nsss(0)='1'  )then
          oVar1S943(0) <='1';
          else
          oVar1S943(0) <='0';
          end if;
        if(cVar2S28S105P031P029P018nsss(0)='1'  OR cVar2S29S105P031P054P017nsss(0)='1'  OR cVar2S30S105P031N054P058nsss(0)='1'  )then
          oVar1S944(0) <='1';
          else
          oVar1S944(0) <='0';
          end if;
        if(cVar2S0S106P008P037P026nsss(0)='1'  OR cVar2S1S106P008N037P053nsss(0)='1'  OR cVar2S2S106N008P019P015nsss(0)='1'  OR cVar2S3S106N008N019P006nsss(0)='1'  )then
          oVar1S945(0) <='1';
          else
          oVar1S945(0) <='0';
          end if;
        if(cVar2S4S106P024nsss(0)='1'  OR cVar2S5S106N024P026P063nsss(0)='1'  OR cVar2S6S106P010P017P016nsss(0)='1'  OR cVar2S7S106P010P017P066nsss(0)='1'  )then
          oVar1S946(0) <='1';
          else
          oVar1S946(0) <='0';
          end if;
        if(cVar2S8S106P051P050nsss(0)='1'  OR cVar2S9S106N051P053nsss(0)='1'  OR cVar2S10S106P023P006nsss(0)='1'  OR cVar2S11S106P023N006P018nsss(0)='1'  )then
          oVar1S947(0) <='1';
          else
          oVar1S947(0) <='0';
          end if;
        if(cVar2S12S106N023P042nsss(0)='1'  OR cVar2S13S106N023P042P021nsss(0)='1'  OR cVar2S14S106P060P063P017nsss(0)='1'  OR cVar2S15S106P060P063P017nsss(0)='1'  )then
          oVar1S948(0) <='1';
          else
          oVar1S948(0) <='0';
          end if;
        if(cVar2S16S106N060P065P037nsss(0)='1'  OR cVar2S17S106N060N065P051nsss(0)='1'  OR cVar2S18S106P002P011nsss(0)='1'  OR cVar2S19S106P002N011P018nsss(0)='1'  )then
          oVar1S949(0) <='1';
          else
          oVar1S949(0) <='0';
          end if;
        if(cVar2S20S106N002P033P007nsss(0)='1'  OR cVar2S21S106N002N033P047nsss(0)='1'  OR cVar2S22S106P033P067nsss(0)='1'  OR cVar2S23S106P059P058nsss(0)='1'  )then
          oVar1S950(0) <='1';
          else
          oVar1S950(0) <='0';
          end if;
        if(cVar2S24S106P059P060nsss(0)='1'  OR cVar2S25S106P058P059P035nsss(0)='1'  OR cVar2S26S106P058N059P011nsss(0)='1'  OR cVar2S27S106P058P014P063nsss(0)='1'  )then
          oVar1S951(0) <='1';
          else
          oVar1S951(0) <='0';
          end if;
        if(cVar1S28S106P036P005P031P020nsss(0)='1'  OR cVar2S29S106P069P060nsss(0)='1'  OR cVar2S30S106N069P061nsss(0)='1'  OR cVar2S31S106N069N061P026nsss(0)='1'  )then
          oVar1S952(0) <='1';
          else
          oVar1S952(0) <='0';
          end if;
        if(cVar2S0S107P061P037P059nsss(0)='1'  OR cVar2S1S107P061P037P066nsss(0)='1'  OR cVar2S2S107P061P037nsss(0)='1'  OR cVar2S3S107P049P069nsss(0)='1'  )then
          oVar1S954(0) <='1';
          else
          oVar1S954(0) <='0';
          end if;
        if(cVar2S4S107P012P032P053nsss(0)='1'  OR cVar2S5S107P012P032P018nsss(0)='1'  OR cVar2S6S107P012P056nsss(0)='1'  OR cVar2S7S107P012N056P032nsss(0)='1'  )then
          oVar1S955(0) <='1';
          else
          oVar1S955(0) <='0';
          end if;
        if(cVar2S8S107P026nsss(0)='1'  OR cVar2S9S107N026P009P027nsss(0)='1'  OR cVar2S10S107P033P003nsss(0)='1'  OR cVar2S11S107P033N003P016nsss(0)='1'  )then
          oVar1S956(0) <='1';
          else
          oVar1S956(0) <='0';
          end if;
        if(cVar2S12S107P032nsss(0)='1'  OR cVar2S13S107N032P058P010nsss(0)='1'  OR cVar2S14S107P010P013nsss(0)='1'  OR cVar2S15S107P010P013P032nsss(0)='1'  )then
          oVar1S957(0) <='1';
          else
          oVar1S957(0) <='0';
          end if;
        if(cVar2S16S107P030P063nsss(0)='1'  OR cVar2S17S107N030P017nsss(0)='1'  OR cVar2S18S107N030P017P005nsss(0)='1'  OR cVar2S19S107P003P062nsss(0)='1'  )then
          oVar1S958(0) <='1';
          else
          oVar1S958(0) <='0';
          end if;
        if(cVar2S20S107N003P017nsss(0)='1'  OR cVar2S21S107P035P055nsss(0)='1'  OR cVar2S22S107P035N055P063nsss(0)='1'  OR cVar2S23S107N035P009nsss(0)='1'  )then
          oVar1S959(0) <='1';
          else
          oVar1S959(0) <='0';
          end if;
        if(cVar2S24S107N035N009P014nsss(0)='1'  OR cVar2S25S107P066P058nsss(0)='1'  OR cVar2S26S107N066P024nsss(0)='1'  OR cVar2S27S107N066N024P015nsss(0)='1'  )then
          oVar1S960(0) <='1';
          else
          oVar1S960(0) <='0';
          end if;
        if(cVar2S28S107P053P030nsss(0)='1'  OR cVar2S29S107P053N030P010nsss(0)='1'  OR cVar2S30S107P023P006P018nsss(0)='1'  OR cVar2S31S107P023N006P042nsss(0)='1'  )then
          oVar1S961(0) <='1';
          else
          oVar1S961(0) <='0';
          end if;
        if(cVar2S32S107N023P059P030nsss(0)='1'  OR cVar2S33S107P026P057P011nsss(0)='1'  )then
          oVar1S962(0) <='1';
          else
          oVar1S962(0) <='0';
          end if;
        if(cVar2S0S108P030P057nsss(0)='1'  OR cVar2S1S108P030P057P061nsss(0)='1'  OR cVar2S2S108P030P029P057nsss(0)='1'  OR cVar2S3S108P029P008nsss(0)='1'  )then
          oVar1S963(0) <='1';
          else
          oVar1S963(0) <='0';
          end if;
        if(cVar2S4S108P029N008P010nsss(0)='1'  OR cVar2S5S108N029P061nsss(0)='1'  OR cVar2S6S108N029N061P030nsss(0)='1'  OR cVar2S7S108P054P015P017nsss(0)='1'  )then
          oVar1S964(0) <='1';
          else
          oVar1S964(0) <='0';
          end if;
        if(cVar2S8S108P054N015P066nsss(0)='1'  OR cVar2S9S108N054P057P030nsss(0)='1'  OR cVar2S10S108P068nsss(0)='1'  OR cVar2S11S108P056P033nsss(0)='1'  )then
          oVar1S965(0) <='1';
          else
          oVar1S965(0) <='0';
          end if;
        if(cVar2S12S108P056P033P019nsss(0)='1'  OR cVar2S13S108P056P010P018nsss(0)='1'  OR cVar2S14S108P061P055nsss(0)='1'  OR cVar2S15S108N061P017nsss(0)='1'  )then
          oVar1S966(0) <='1';
          else
          oVar1S966(0) <='0';
          end if;
        if(cVar2S16S108P060nsss(0)='1'  OR cVar2S17S108P060P059P033nsss(0)='1'  OR cVar2S18S108P060P004P056nsss(0)='1'  OR cVar2S19S108N060P068P018nsss(0)='1'  )then
          oVar1S967(0) <='1';
          else
          oVar1S967(0) <='0';
          end if;
        if(cVar2S20S108P061nsss(0)='1'  OR cVar2S21S108N061P014P005nsss(0)='1'  OR cVar2S22S108N061P014P013nsss(0)='1'  OR cVar2S23S108P069P034nsss(0)='1'  )then
          oVar1S968(0) <='1';
          else
          oVar1S968(0) <='0';
          end if;
        if(cVar2S24S108P069N034P019nsss(0)='1'  OR cVar2S25S108N069P063P014nsss(0)='1'  OR cVar2S26S108P016nsss(0)='1'  OR cVar2S27S108N016P015P022nsss(0)='1'  )then
          oVar1S969(0) <='1';
          else
          oVar1S969(0) <='0';
          end if;
        if(cVar2S28S108P043P008nsss(0)='1'  OR cVar2S29S108P043N008P025nsss(0)='1'  OR cVar2S30S108P065nsss(0)='1'  OR cVar2S31S108N065P018nsss(0)='1'  )then
          oVar1S970(0) <='1';
          else
          oVar1S970(0) <='0';
          end if;
        if(cVar2S32S108N065N018P011nsss(0)='1'  OR cVar2S33S108P057nsss(0)='1'  OR cVar2S34S108N057P013P066nsss(0)='1'  OR cVar2S35S108P030nsss(0)='1'  )then
          oVar1S971(0) <='1';
          else
          oVar1S971(0) <='0';
          end if;
        if(cVar2S36S108N030P051P006nsss(0)='1'  OR cVar2S37S108P017P009nsss(0)='1'  OR cVar2S38S108P017N009P008nsss(0)='1'  OR cVar2S39S108N017P015P011nsss(0)='1'  )then
          oVar1S972(0) <='1';
          else
          oVar1S972(0) <='0';
          end if;
        if(cVar2S0S109P057P014nsss(0)='1'  OR cVar2S1S109P057N014P018nsss(0)='1'  OR cVar2S2S109N057P048nsss(0)='1'  OR cVar2S3S109N057P048P025nsss(0)='1'  )then
          oVar1S974(0) <='1';
          else
          oVar1S974(0) <='0';
          end if;
        if(cVar2S4S109P052P067P035nsss(0)='1'  OR cVar2S5S109P031P013nsss(0)='1'  OR cVar2S6S109N031P029nsss(0)='1'  OR cVar2S7S109N031N029P015nsss(0)='1'  )then
          oVar1S975(0) <='1';
          else
          oVar1S975(0) <='0';
          end if;
        if(cVar2S8S109P047nsss(0)='1'  OR cVar2S9S109P009P063nsss(0)='1'  OR cVar2S10S109P009N063P067nsss(0)='1'  OR cVar2S11S109N009P036P037nsss(0)='1'  )then
          oVar1S976(0) <='1';
          else
          oVar1S976(0) <='0';
          end if;
        if(cVar1S12S109P064P068P051P017nsss(0)='1'  OR cVar2S13S109P013P058nsss(0)='1'  OR cVar2S14S109P013N058P018nsss(0)='1'  OR cVar2S15S109N013P052P016nsss(0)='1'  )then
          oVar1S977(0) <='1';
          else
          oVar1S977(0) <='0';
          end if;
        if(cVar2S16S109N013N052P030nsss(0)='1'  OR cVar2S17S109P008P011nsss(0)='1'  OR cVar2S18S109P008P011P056nsss(0)='1'  OR cVar2S19S109N008P009nsss(0)='1'  )then
          oVar1S978(0) <='1';
          else
          oVar1S978(0) <='0';
          end if;
        if(cVar2S20S109P003nsss(0)='1'  OR cVar2S21S109N003P007nsss(0)='1'  OR cVar2S22S109N003N007P045nsss(0)='1'  OR cVar2S23S109P042P004nsss(0)='1'  )then
          oVar1S979(0) <='1';
          else
          oVar1S979(0) <='0';
          end if;
        if(cVar2S24S109P042N004P006nsss(0)='1'  OR cVar2S25S109N042P006P052nsss(0)='1'  OR cVar2S26S109P047P024P026nsss(0)='1'  OR cVar2S27S109P047N024P026nsss(0)='1'  )then
          oVar1S980(0) <='1';
          else
          oVar1S980(0) <='0';
          end if;
        if(cVar2S28S109N047P024P005nsss(0)='1'  OR cVar2S29S109P047P006nsss(0)='1'  )then
          oVar1S981(0) <='1';
          else
          oVar1S981(0) <='0';
          end if;
        if(cVar2S0S110P050P042nsss(0)='1'  OR cVar2S1S110P050P058nsss(0)='1'  OR cVar2S2S110P031nsss(0)='1'  OR cVar1S3S110P064P056P052P009nsss(0)='1'  )then
          oVar1S982(0) <='1';
          else
          oVar1S982(0) <='0';
          end if;
        if(cVar2S4S110P015nsss(0)='1'  OR cVar2S5S110N015P029P050nsss(0)='1'  OR cVar2S6S110P016P065nsss(0)='1'  OR cVar2S7S110P016N065P068nsss(0)='1'  )then
          oVar1S983(0) <='1';
          else
          oVar1S983(0) <='0';
          end if;
        if(cVar2S8S110N016P063P034nsss(0)='1'  OR cVar2S9S110N016P063P034nsss(0)='1'  OR cVar2S10S110P024P045nsss(0)='1'  OR cVar2S11S110N024P027nsss(0)='1'  )then
          oVar1S984(0) <='1';
          else
          oVar1S984(0) <='0';
          end if;
        if(cVar2S12S110N024N027P033nsss(0)='1'  OR cVar2S13S110P036nsss(0)='1'  OR cVar2S14S110N036P016nsss(0)='1'  OR cVar2S15S110N036P016P019nsss(0)='1'  )then
          oVar1S985(0) <='1';
          else
          oVar1S985(0) <='0';
          end if;
        if(cVar2S16S110P051P019nsss(0)='1'  OR cVar2S17S110P051N019P069nsss(0)='1'  OR cVar2S18S110N051P046P010nsss(0)='1'  OR cVar2S19S110P019P028P010nsss(0)='1'  )then
          oVar1S986(0) <='1';
          else
          oVar1S986(0) <='0';
          end if;
        if(cVar2S20S110P019N028psss(0)='1'  OR cVar2S21S110P019P068P037nsss(0)='1'  OR cVar2S22S110P019N068P063nsss(0)='1'  OR cVar2S23S110P009P016nsss(0)='1'  )then
          oVar1S987(0) <='1';
          else
          oVar1S987(0) <='0';
          end if;
        if(cVar2S24S110P023nsss(0)='1'  OR cVar2S25S110P036P015P016nsss(0)='1'  OR cVar2S26S110P034nsss(0)='1'  OR cVar2S27S110N034P048P000nsss(0)='1'  )then
          oVar1S988(0) <='1';
          else
          oVar1S988(0) <='0';
          end if;
        if(cVar2S0S111P015P045nsss(0)='1'  OR cVar2S1S111N015P058nsss(0)='1'  OR cVar2S2S111N015P058P032nsss(0)='1'  OR cVar2S3S111P065nsss(0)='1'  )then
          oVar1S990(0) <='1';
          else
          oVar1S990(0) <='0';
          end if;
        if(cVar2S4S111N065P011P015nsss(0)='1'  OR cVar1S5S111P064P033P041P003nsss(0)='1'  OR cVar2S6S111P034P003nsss(0)='1'  OR cVar2S7S111N034P003P019nsss(0)='1'  )then
          oVar1S991(0) <='1';
          else
          oVar1S991(0) <='0';
          end if;
        if(cVar2S8S111N034N003P014nsss(0)='1'  OR cVar2S9S111P020P057nsss(0)='1'  OR cVar2S10S111P020N057P000nsss(0)='1'  OR cVar2S11S111P020P015P010nsss(0)='1'  )then
          oVar1S992(0) <='1';
          else
          oVar1S992(0) <='0';
          end if;
        if(cVar2S12S111P020P015P012nsss(0)='1'  OR cVar2S13S111P006P068nsss(0)='1'  OR cVar2S14S111N006P001P069nsss(0)='1'  OR cVar2S15S111P011nsss(0)='1'  )then
          oVar1S993(0) <='1';
          else
          oVar1S993(0) <='0';
          end if;
        if(cVar2S16S111P065P018P068nsss(0)='1'  OR cVar2S17S111P065N018P015nsss(0)='1'  OR cVar2S18S111P049P067nsss(0)='1'  OR cVar2S19S111P049N067P017nsss(0)='1'  )then
          oVar1S994(0) <='1';
          else
          oVar1S994(0) <='0';
          end if;
        if(cVar2S20S111N049P017P068nsss(0)='1'  OR cVar2S21S111N049N017P003nsss(0)='1'  OR cVar2S22S111P004P017nsss(0)='1'  OR cVar2S23S111P004N017P002nsss(0)='1'  )then
          oVar1S995(0) <='1';
          else
          oVar1S995(0) <='0';
          end if;
        if(cVar2S24S111N004P008nsss(0)='1'  OR cVar2S25S111P042P053nsss(0)='1'  OR cVar2S26S111P061P014P012nsss(0)='1'  OR cVar2S27S111P061P052nsss(0)='1'  )then
          oVar1S996(0) <='1';
          else
          oVar1S996(0) <='0';
          end if;
        if(cVar2S0S112P009P033P056nsss(0)='1'  OR cVar2S1S112P009P033P061nsss(0)='1'  OR cVar2S2S112P009P065P013nsss(0)='1'  OR cVar2S3S112P009N065P032nsss(0)='1'  )then
          oVar1S998(0) <='1';
          else
          oVar1S998(0) <='0';
          end if;
        if(cVar2S4S112P012P009nsss(0)='1'  OR cVar2S5S112P012N009P017nsss(0)='1'  OR cVar2S6S112N012P069nsss(0)='1'  OR cVar2S7S112N012P069P035nsss(0)='1'  )then
          oVar1S999(0) <='1';
          else
          oVar1S999(0) <='0';
          end if;
        if(cVar2S8S112P066P049nsss(0)='1'  OR cVar2S9S112P066N049P052nsss(0)='1'  OR cVar2S10S112P066P050nsss(0)='1'  OR cVar2S11S112P063nsss(0)='1'  )then
          oVar1S1000(0) <='1';
          else
          oVar1S1000(0) <='0';
          end if;
        if(cVar2S12S112N063P015P017nsss(0)='1'  OR cVar2S13S112N063N015P052nsss(0)='1'  OR cVar2S14S112P024P004nsss(0)='1'  OR cVar2S15S112P024N004P006nsss(0)='1'  )then
          oVar1S1001(0) <='1';
          else
          oVar1S1001(0) <='0';
          end if;
        if(cVar2S16S112P069P061P019nsss(0)='1'  OR cVar2S17S112P061P063nsss(0)='1'  OR cVar2S18S112P061N063P056nsss(0)='1'  OR cVar2S19S112P061P019P015nsss(0)='1'  )then
          oVar1S1002(0) <='1';
          else
          oVar1S1002(0) <='0';
          end if;
        if(cVar2S20S112P067P051nsss(0)='1'  OR cVar2S21S112P067N051P063nsss(0)='1'  OR cVar2S22S112P024nsss(0)='1'  OR cVar2S23S112N024P035P009nsss(0)='1'  )then
          oVar1S1003(0) <='1';
          else
          oVar1S1003(0) <='0';
          end if;
        if(cVar2S24S112N024N035P056nsss(0)='1'  OR cVar2S25S112P037nsss(0)='1'  OR cVar2S26S112N037P063P012nsss(0)='1'  OR cVar2S27S112P013P061P060nsss(0)='1'  )then
          oVar1S1004(0) <='1';
          else
          oVar1S1004(0) <='0';
          end if;
        if(cVar2S28S112P013P003nsss(0)='1'  OR cVar2S29S112P057P011P038nsss(0)='1'  OR cVar2S30S112P057P011P050nsss(0)='1'  OR cVar2S31S112P057P059P035nsss(0)='1'  )then
          oVar1S1005(0) <='1';
          else
          oVar1S1005(0) <='0';
          end if;
        if(cVar2S32S112P057N059P003nsss(0)='1'  OR cVar2S33S112P001P066nsss(0)='1'  OR cVar2S34S112P001P066P037nsss(0)='1'  OR cVar2S35S112N001P065P060nsss(0)='1'  )then
          oVar1S1006(0) <='1';
          else
          oVar1S1006(0) <='0';
          end if;
        if(cVar2S36S112N001N065P015nsss(0)='1'  OR cVar2S37S112P055P011nsss(0)='1'  )then
          oVar1S1007(0) <='1';
          else
          oVar1S1007(0) <='0';
          end if;
        if(cVar2S0S113P057P055nsss(0)='1'  OR cVar2S1S113P057P055P058nsss(0)='1'  OR cVar2S2S113P057P012nsss(0)='1'  OR cVar2S3S113P057N012P003nsss(0)='1'  )then
          oVar1S1008(0) <='1';
          else
          oVar1S1008(0) <='0';
          end if;
        if(cVar2S4S113P055P029nsss(0)='1'  OR cVar2S5S113P055N029P006nsss(0)='1'  OR cVar2S6S113N055P008P007nsss(0)='1'  OR cVar2S7S113N055N008P006nsss(0)='1'  )then
          oVar1S1009(0) <='1';
          else
          oVar1S1009(0) <='0';
          end if;
        if(cVar2S8S113P052P016nsss(0)='1'  OR cVar2S9S113P052P016P064nsss(0)='1'  OR cVar2S10S113P057P013nsss(0)='1'  OR cVar2S11S113P057N013P009nsss(0)='1'  )then
          oVar1S1010(0) <='1';
          else
          oVar1S1010(0) <='0';
          end if;
        if(cVar2S12S113P057P031P013nsss(0)='1'  OR cVar2S13S113P030P056nsss(0)='1'  OR cVar2S14S113P030N056P016nsss(0)='1'  OR cVar2S15S113N030P062P016nsss(0)='1'  )then
          oVar1S1011(0) <='1';
          else
          oVar1S1011(0) <='0';
          end if;
        if(cVar2S16S113N030P062P068nsss(0)='1'  OR cVar2S17S113P012nsss(0)='1'  OR cVar2S18S113N012P010nsss(0)='1'  OR cVar2S19S113N012N010P068nsss(0)='1'  )then
          oVar1S1012(0) <='1';
          else
          oVar1S1012(0) <='0';
          end if;
        if(cVar2S20S113P064P032nsss(0)='1'  OR cVar2S21S113P064N032P013nsss(0)='1'  OR cVar2S22S113N064P034P058nsss(0)='1'  OR cVar2S23S113N064N034P068nsss(0)='1'  )then
          oVar1S1013(0) <='1';
          else
          oVar1S1013(0) <='0';
          end if;
        if(cVar2S24S113P016P052P008nsss(0)='1'  OR cVar2S25S113P016N052P025nsss(0)='1'  OR cVar2S26S113P016P035P068nsss(0)='1'  OR cVar2S27S113P016N035P007nsss(0)='1'  )then
          oVar1S1014(0) <='1';
          else
          oVar1S1014(0) <='0';
          end if;
        if(cVar2S28S113P012nsss(0)='1'  OR cVar2S29S113P037P032P019nsss(0)='1'  OR cVar2S30S113P037N032P029nsss(0)='1'  OR cVar2S31S113N037P033P019nsss(0)='1'  )then
          oVar1S1015(0) <='1';
          else
          oVar1S1015(0) <='0';
          end if;
        if(cVar2S32S113N037N033P030nsss(0)='1'  OR cVar1S33S113P014P018P022P037nsss(0)='1'  OR cVar2S34S113P066P017nsss(0)='1'  OR cVar2S35S113P034P061P023nsss(0)='1'  )then
          oVar1S1016(0) <='1';
          else
          oVar1S1016(0) <='0';
          end if;
        if(cVar2S36S113P034P061P016nsss(0)='1'  OR cVar2S37S113P034P016P063nsss(0)='1'  OR cVar2S38S113P034N016P063nsss(0)='1'  OR cVar2S39S113P064P007P008nsss(0)='1'  )then
          oVar1S1017(0) <='1';
          else
          oVar1S1017(0) <='0';
          end if;
        if(cVar2S40S113P064P007P055nsss(0)='1'  OR cVar2S41S113P064P068P019nsss(0)='1'  OR cVar2S42S113P064N068P024nsss(0)='1'  OR cVar2S43S113P030P008P012nsss(0)='1'  )then
          oVar1S1018(0) <='1';
          else
          oVar1S1018(0) <='0';
          end if;
        if(cVar2S44S113P030P012nsss(0)='1'  )then
          oVar1S1019(0) <='1';
          else
          oVar1S1019(0) <='0';
          end if;
        if(cVar2S0S114P033nsss(0)='1'  OR cVar2S1S114P049P009nsss(0)='1'  OR cVar2S2S114P049N009P035nsss(0)='1'  OR cVar2S3S114N049P060nsss(0)='1'  )then
          oVar1S1020(0) <='1';
          else
          oVar1S1020(0) <='0';
          end if;
        if(cVar2S4S114N049P060P033nsss(0)='1'  OR cVar2S5S114P013P003nsss(0)='1'  OR cVar2S6S114P013N003P067nsss(0)='1'  OR cVar2S7S114P013P036nsss(0)='1'  )then
          oVar1S1021(0) <='1';
          else
          oVar1S1021(0) <='0';
          end if;
        if(cVar2S8S114P033P059P008nsss(0)='1'  OR cVar2S9S114N033P028P035nsss(0)='1'  OR cVar2S10S114P007P059P019nsss(0)='1'  OR cVar2S11S114P007N059P065nsss(0)='1'  )then
          oVar1S1022(0) <='1';
          else
          oVar1S1022(0) <='0';
          end if;
        if(cVar2S12S114N007P035nsss(0)='1'  OR cVar2S13S114N007N035P062nsss(0)='1'  OR cVar2S14S114P029nsss(0)='1'  OR cVar2S15S114N029P036nsss(0)='1'  )then
          oVar1S1023(0) <='1';
          else
          oVar1S1023(0) <='0';
          end if;
        if(cVar2S16S114P013P028nsss(0)='1'  OR cVar2S17S114P013N028P012nsss(0)='1'  OR cVar2S18S114P013P016P014nsss(0)='1'  OR cVar2S19S114P021P011nsss(0)='1'  )then
          oVar1S1024(0) <='1';
          else
          oVar1S1024(0) <='0';
          end if;
        if(cVar2S20S114P021P011P012nsss(0)='1'  OR cVar2S21S114P021P010P037nsss(0)='1'  OR cVar2S22S114P033P032P036nsss(0)='1'  OR cVar2S23S114P033N032P034nsss(0)='1'  )then
          oVar1S1025(0) <='1';
          else
          oVar1S1025(0) <='0';
          end if;
        if(cVar2S24S114P033P032P007nsss(0)='1'  OR cVar2S25S114P033P032P059nsss(0)='1'  OR cVar2S26S114P034P040P010nsss(0)='1'  OR cVar2S27S114P034P017P016nsss(0)='1'  )then
          oVar1S1026(0) <='1';
          else
          oVar1S1026(0) <='0';
          end if;
        if(cVar2S28S114P034N017P033nsss(0)='1'  OR cVar2S29S114P056P012nsss(0)='1'  OR cVar2S30S114P056N012P037nsss(0)='1'  OR cVar2S31S114P056P012P057nsss(0)='1'  )then
          oVar1S1027(0) <='1';
          else
          oVar1S1027(0) <='0';
          end if;
        if(cVar2S32S114P013P060P059nsss(0)='1'  OR cVar2S33S114N013P016P037nsss(0)='1'  OR cVar2S34S114N013P016P068nsss(0)='1'  OR cVar2S35S114P007nsss(0)='1'  )then
          oVar1S1028(0) <='1';
          else
          oVar1S1028(0) <='0';
          end if;
        if(cVar2S36S114P007P062P015nsss(0)='1'  OR cVar2S37S114P017P015P063nsss(0)='1'  OR cVar2S38S114P017P044nsss(0)='1'  )then
          oVar1S1029(0) <='1';
          else
          oVar1S1029(0) <='0';
          end if;
        if(cVar2S0S115P028P019nsss(0)='1'  OR cVar2S1S115P028N019P068nsss(0)='1'  OR cVar2S2S115N028P037nsss(0)='1'  OR cVar2S3S115N028N037P016nsss(0)='1'  )then
          oVar1S1030(0) <='1';
          else
          oVar1S1030(0) <='0';
          end if;
        if(cVar2S4S115P016P037P059nsss(0)='1'  OR cVar2S5S115P016P037P062nsss(0)='1'  OR cVar2S6S115N016P060nsss(0)='1'  OR cVar2S7S115P011P013P036nsss(0)='1'  )then
          oVar1S1031(0) <='1';
          else
          oVar1S1031(0) <='0';
          end if;
        if(cVar2S8S115P011N013P054nsss(0)='1'  OR cVar2S9S115P011P066nsss(0)='1'  OR cVar2S10S115P011P066P025nsss(0)='1'  OR cVar2S11S115P019P036P015nsss(0)='1'  )then
          oVar1S1032(0) <='1';
          else
          oVar1S1032(0) <='0';
          end if;
        if(cVar2S12S115P019N036P010nsss(0)='1'  OR cVar2S13S115N019P062P066nsss(0)='1'  OR cVar2S14S115P036P030nsss(0)='1'  OR cVar2S15S115P036N030P012nsss(0)='1'  )then
          oVar1S1033(0) <='1';
          else
          oVar1S1033(0) <='0';
          end if;
        if(cVar2S16S115P036P053P019nsss(0)='1'  OR cVar2S17S115P032P069nsss(0)='1'  OR cVar2S18S115P032N069P035nsss(0)='1'  OR cVar2S19S115N032P001nsss(0)='1'  )then
          oVar1S1034(0) <='1';
          else
          oVar1S1034(0) <='0';
          end if;
        if(cVar2S20S115P006nsss(0)='1'  OR cVar2S21S115N006P016P008nsss(0)='1'  OR cVar2S22S115N006N016P011nsss(0)='1'  OR cVar2S23S115P045nsss(0)='1'  )then
          oVar1S1035(0) <='1';
          else
          oVar1S1035(0) <='0';
          end if;
        if(cVar2S24S115N045P002P015nsss(0)='1'  OR cVar2S25S115N045N002P051nsss(0)='1'  OR cVar2S26S115P007P047nsss(0)='1'  OR cVar2S27S115P007N047P021nsss(0)='1'  )then
          oVar1S1036(0) <='1';
          else
          oVar1S1036(0) <='0';
          end if;
        if(cVar2S28S115P007P059P013nsss(0)='1'  OR cVar2S29S115P061nsss(0)='1'  OR cVar2S30S115N061P037P035nsss(0)='1'  OR cVar2S31S115P005nsss(0)='1'  )then
          oVar1S1037(0) <='1';
          else
          oVar1S1037(0) <='0';
          end if;
        if(cVar2S32S115N005P009nsss(0)='1'  OR cVar2S33S115P066nsss(0)='1'  OR cVar2S34S115N066P067nsss(0)='1'  OR cVar2S35S115P059P065nsss(0)='1'  )then
          oVar1S1038(0) <='1';
          else
          oVar1S1038(0) <='0';
          end if;
        if(cVar2S36S115N059P028nsss(0)='1'  OR cVar2S37S115N059N028P032nsss(0)='1'  OR cVar2S38S115P033P009nsss(0)='1'  OR cVar2S39S115P033N009P060nsss(0)='1'  )then
          oVar1S1039(0) <='1';
          else
          oVar1S1039(0) <='0';
          end if;
        if(cVar2S40S115N033P028P067nsss(0)='1'  OR cVar2S41S115P058P032P060nsss(0)='1'  OR cVar2S42S115P058N032P031nsss(0)='1'  )then
          oVar1S1040(0) <='1';
          else
          oVar1S1040(0) <='0';
          end if;
        if(cVar2S0S116P026nsss(0)='1'  OR cVar2S1S116N026P006nsss(0)='1'  OR cVar2S2S116N026N006P058nsss(0)='1'  OR cVar2S3S116P046nsss(0)='1'  )then
          oVar1S1041(0) <='1';
          else
          oVar1S1041(0) <='0';
          end if;
        if(cVar2S4S116N046P069P010nsss(0)='1'  OR cVar2S5S116N046P069psss(0)='1'  OR cVar2S6S116P048P028nsss(0)='1'  OR cVar2S7S116P048N028P061nsss(0)='1'  )then
          oVar1S1042(0) <='1';
          else
          oVar1S1042(0) <='0';
          end if;
        if(cVar2S8S116P048P006P017nsss(0)='1'  OR cVar2S9S116P048N006P026nsss(0)='1'  OR cVar2S10S116P012nsss(0)='1'  OR cVar2S11S116N012P016nsss(0)='1'  )then
          oVar1S1043(0) <='1';
          else
          oVar1S1043(0) <='0';
          end if;
        if(cVar2S12S116P035P036nsss(0)='1'  OR cVar2S13S116P015P036P069nsss(0)='1'  OR cVar2S14S116P015N036P037nsss(0)='1'  OR cVar2S15S116P015P065P064nsss(0)='1'  )then
          oVar1S1044(0) <='1';
          else
          oVar1S1044(0) <='0';
          end if;
        if(cVar2S16S116P015N065P017nsss(0)='1'  OR cVar2S17S116P002P067P059nsss(0)='1'  OR cVar2S18S116P002N067P013nsss(0)='1'  OR cVar2S19S116P002N015P019nsss(0)='1'  )then
          oVar1S1045(0) <='1';
          else
          oVar1S1045(0) <='0';
          end if;
        if(cVar2S20S116P017P037P016nsss(0)='1'  OR cVar2S21S116P017P037P015nsss(0)='1'  OR cVar2S22S116P017P016nsss(0)='1'  OR cVar2S23S116P017P016P037nsss(0)='1'  )then
          oVar1S1046(0) <='1';
          else
          oVar1S1046(0) <='0';
          end if;
        if(cVar2S24S116P012P015nsss(0)='1'  OR cVar2S25S116N012P017P068nsss(0)='1'  OR cVar2S26S116N012N017P015nsss(0)='1'  OR cVar2S27S116P045P047nsss(0)='1'  )then
          oVar1S1047(0) <='1';
          else
          oVar1S1047(0) <='0';
          end if;
        if(cVar2S28S116P045N047P019nsss(0)='1'  OR cVar2S29S116N045P043P041nsss(0)='1'  OR cVar2S30S116P060P036nsss(0)='1'  OR cVar2S31S116N060P034P067nsss(0)='1'  )then
          oVar1S1048(0) <='1';
          else
          oVar1S1048(0) <='0';
          end if;
        if(cVar2S32S116P010P034P054nsss(0)='1'  OR cVar2S33S116P010N034P065nsss(0)='1'  OR cVar2S34S116P010P013P068nsss(0)='1'  OR cVar2S35S116P005P047P030nsss(0)='1'  )then
          oVar1S1049(0) <='1';
          else
          oVar1S1049(0) <='0';
          end if;
        if(cVar2S36S116P058P008nsss(0)='1'  OR cVar2S37S116P058N008P020nsss(0)='1'  OR cVar2S38S116N058P008P037nsss(0)='1'  OR cVar2S39S116N058P008P028nsss(0)='1'  )then
          oVar1S1050(0) <='1';
          else
          oVar1S1050(0) <='0';
          end if;
        if(cVar2S40S116P033P036P041nsss(0)='1'  OR cVar2S41S116P033N036P039nsss(0)='1'  )then
          oVar1S1051(0) <='1';
          else
          oVar1S1051(0) <='0';
          end if;
        if(cVar2S0S117P016nsss(0)='1'  OR cVar2S1S117N016P033nsss(0)='1'  OR cVar2S2S117P035P064nsss(0)='1'  OR cVar2S3S117N035P013P019nsss(0)='1'  )then
          oVar1S1052(0) <='1';
          else
          oVar1S1052(0) <='0';
          end if;
        if(cVar2S4S117P065P028nsss(0)='1'  OR cVar2S5S117N065P019P017nsss(0)='1'  OR cVar2S6S117P058nsss(0)='1'  OR cVar2S7S117P018P051P049nsss(0)='1'  )then
          oVar1S1053(0) <='1';
          else
          oVar1S1053(0) <='0';
          end if;
        if(cVar2S8S117N018P049P048nsss(0)='1'  OR cVar2S9S117N018N049P053nsss(0)='1'  OR cVar2S10S117P031P007P009nsss(0)='1'  OR cVar2S11S117P031P007P019nsss(0)='1'  )then
          oVar1S1054(0) <='1';
          else
          oVar1S1054(0) <='0';
          end if;
        if(cVar2S12S117N031P035nsss(0)='1'  OR cVar2S13S117N031N035P043nsss(0)='1'  OR cVar2S14S117P035P062nsss(0)='1'  OR cVar2S15S117P035P037P016nsss(0)='1'  )then
          oVar1S1055(0) <='1';
          else
          oVar1S1055(0) <='0';
          end if;
        if(cVar2S16S117P027nsss(0)='1'  OR cVar2S17S117P010P002P013nsss(0)='1'  OR cVar2S18S117P010P002P037nsss(0)='1'  OR cVar2S19S117P010P054P011nsss(0)='1'  )then
          oVar1S1056(0) <='1';
          else
          oVar1S1056(0) <='0';
          end if;
        if(cVar2S20S117P010N054P050nsss(0)='1'  OR cVar2S21S117P024P019nsss(0)='1'  OR cVar2S22S117N024P010nsss(0)='1'  OR cVar2S23S117P019nsss(0)='1'  )then
          oVar1S1057(0) <='1';
          else
          oVar1S1057(0) <='0';
          end if;
        if(cVar2S24S117P019P049nsss(0)='1'  OR cVar2S25S117P069P016nsss(0)='1'  OR cVar2S26S117N069P048nsss(0)='1'  OR cVar1S27S117P066P018P049P051nsss(0)='1'  )then
          oVar1S1058(0) <='1';
          else
          oVar1S1058(0) <='0';
          end if;
        if(cVar2S28S117P068P009P017nsss(0)='1'  OR cVar2S29S117P068P009P037nsss(0)='1'  OR cVar2S30S117P016P069nsss(0)='1'  OR cVar2S31S117P016N069P011nsss(0)='1'  )then
          oVar1S1059(0) <='1';
          else
          oVar1S1059(0) <='0';
          end if;
        if(cVar2S32S117P016P059P015nsss(0)='1'  OR cVar2S33S117P016P026P036nsss(0)='1'  OR cVar2S34S117N016P034P046nsss(0)='1'  OR cVar2S35S117N016P034P019nsss(0)='1'  )then
          oVar1S1060(0) <='1';
          else
          oVar1S1060(0) <='0';
          end if;
        if(cVar2S0S118P064P063nsss(0)='1'  OR cVar2S1S118P006P061P042nsss(0)='1'  OR cVar2S2S118P006P061P060nsss(0)='1'  OR cVar2S3S118P006P017P015nsss(0)='1'  )then
          oVar1S1062(0) <='1';
          else
          oVar1S1062(0) <='0';
          end if;
        if(cVar2S4S118P016P017nsss(0)='1'  OR cVar2S5S118P011nsss(0)='1'  OR cVar2S6S118N011P013nsss(0)='1'  OR cVar2S7S118P068P036nsss(0)='1'  )then
          oVar1S1063(0) <='1';
          else
          oVar1S1063(0) <='0';
          end if;
        if(cVar2S8S118P068P036P042nsss(0)='1'  OR cVar2S9S118P068P018P017nsss(0)='1'  OR cVar2S10S118P068N018P055nsss(0)='1'  OR cVar2S11S118P066P034nsss(0)='1'  )then
          oVar1S1064(0) <='1';
          else
          oVar1S1064(0) <='0';
          end if;
        if(cVar2S12S118P066P034P012nsss(0)='1'  OR cVar2S13S118N066P030P018nsss(0)='1'  OR cVar2S14S118P048P029nsss(0)='1'  OR cVar2S15S118P048N029P011nsss(0)='1'  )then
          oVar1S1065(0) <='1';
          else
          oVar1S1065(0) <='0';
          end if;
        if(cVar2S16S118P048P025nsss(0)='1'  OR cVar2S17S118P048P066P037nsss(0)='1'  OR cVar2S18S118P048P066P026nsss(0)='1'  OR cVar2S19S118N048P045nsss(0)='1'  )then
          oVar1S1066(0) <='1';
          else
          oVar1S1066(0) <='0';
          end if;
        if(cVar2S20S118N048N045P062nsss(0)='1'  OR cVar2S21S118P063nsss(0)='1'  OR cVar2S22S118N063P019nsss(0)='1'  OR cVar2S23S118P006P065nsss(0)='1'  )then
          oVar1S1067(0) <='1';
          else
          oVar1S1067(0) <='0';
          end if;
        if(cVar2S24S118P006P028nsss(0)='1'  OR cVar2S25S118P006N028P056nsss(0)='1'  OR cVar2S26S118P008P033P036nsss(0)='1'  OR cVar2S27S118P008N033P005nsss(0)='1'  )then
          oVar1S1068(0) <='1';
          else
          oVar1S1068(0) <='0';
          end if;
        if(cVar2S28S118P008P060P036nsss(0)='1'  OR cVar1S29S118P035N046P022P065nsss(0)='1'  OR cVar2S30S118P013nsss(0)='1'  OR cVar2S31S118N013P006nsss(0)='1'  )then
          oVar1S1069(0) <='1';
          else
          oVar1S1069(0) <='0';
          end if;
        if(cVar2S0S119P001P026nsss(0)='1'  OR cVar2S1S119P001P026P067nsss(0)='1'  OR cVar2S2S119P052P061nsss(0)='1'  OR cVar2S3S119P036P018nsss(0)='1'  )then
          oVar1S1071(0) <='1';
          else
          oVar1S1071(0) <='0';
          end if;
        if(cVar2S4S119N036P050P019nsss(0)='1'  OR cVar2S5S119N036N050P011nsss(0)='1'  OR cVar2S6S119P034P019P030nsss(0)='1'  OR cVar2S7S119N034P069P066nsss(0)='1'  )then
          oVar1S1072(0) <='1';
          else
          oVar1S1072(0) <='0';
          end if;
        if(cVar2S8S119N034N069P050nsss(0)='1'  OR cVar2S9S119P036P068P008nsss(0)='1'  OR cVar2S10S119P036N068P066nsss(0)='1'  OR cVar2S11S119P036P053P022nsss(0)='1'  )then
          oVar1S1073(0) <='1';
          else
          oVar1S1073(0) <='0';
          end if;
        if(cVar2S12S119P024P047nsss(0)='1'  OR cVar2S13S119P024N047P017nsss(0)='1'  OR cVar2S14S119N024P052nsss(0)='1'  OR cVar2S15S119N024N052P013nsss(0)='1'  )then
          oVar1S1074(0) <='1';
          else
          oVar1S1074(0) <='0';
          end if;
        if(cVar2S16S119P057P053nsss(0)='1'  OR cVar2S17S119N057P009P069nsss(0)='1'  OR cVar2S18S119P060P066nsss(0)='1'  OR cVar2S19S119P060P066P053nsss(0)='1'  )then
          oVar1S1075(0) <='1';
          else
          oVar1S1075(0) <='0';
          end if;
        if(cVar2S20S119P060P057P017nsss(0)='1'  OR cVar2S21S119P059P018P019nsss(0)='1'  OR cVar2S22S119P059P037nsss(0)='1'  OR cVar2S23S119P035P034P013nsss(0)='1'  )then
          oVar1S1076(0) <='1';
          else
          oVar1S1076(0) <='0';
          end if;
        if(cVar2S24S119P035P034P017nsss(0)='1'  OR cVar2S25S119P035P009P066nsss(0)='1'  OR cVar2S26S119P063P067P035nsss(0)='1'  OR cVar2S27S119P063P067P018nsss(0)='1'  )then
          oVar1S1077(0) <='1';
          else
          oVar1S1077(0) <='0';
          end if;
        if(cVar2S28S119P063P069P019nsss(0)='1'  OR cVar2S29S119P063N069P004nsss(0)='1'  OR cVar2S30S119P063P036nsss(0)='1'  OR cVar2S31S119P063N036P034nsss(0)='1'  )then
          oVar1S1078(0) <='1';
          else
          oVar1S1078(0) <='0';
          end if;
        if(cVar2S32S119P066P019nsss(0)='1'  OR cVar1S33S119P065P008N011P056nsss(0)='1'  OR cVar2S34S119P019P015P067nsss(0)='1'  OR cVar2S35S119N019P058nsss(0)='1'  )then
          oVar1S1079(0) <='1';
          else
          oVar1S1079(0) <='0';
          end if;
        if(cVar2S0S120P017P019nsss(0)='1'  OR cVar2S1S120P017P019P013nsss(0)='1'  OR cVar2S2S120P017P060nsss(0)='1'  OR cVar2S3S120P017N060P034nsss(0)='1'  )then
          oVar1S1081(0) <='1';
          else
          oVar1S1081(0) <='0';
          end if;
        if(cVar2S4S120P068P056nsss(0)='1'  OR cVar2S5S120P068P036P061nsss(0)='1'  OR cVar2S6S120P018P069P036nsss(0)='1'  OR cVar2S7S120P018N069psss(0)='1'  )then
          oVar1S1082(0) <='1';
          else
          oVar1S1082(0) <='0';
          end if;
        if(cVar2S8S120P018P017nsss(0)='1'  OR cVar2S9S120P018P017P035nsss(0)='1'  OR cVar2S10S120P052nsss(0)='1'  OR cVar2S11S120N052P031nsss(0)='1'  )then
          oVar1S1083(0) <='1';
          else
          oVar1S1083(0) <='0';
          end if;
        if(cVar2S12S120N052P031P013nsss(0)='1'  OR cVar2S13S120P016P068nsss(0)='1'  OR cVar2S14S120P016N068P018nsss(0)='1'  OR cVar2S15S120P016P014nsss(0)='1'  )then
          oVar1S1084(0) <='1';
          else
          oVar1S1084(0) <='0';
          end if;
        if(cVar2S16S120P014P017nsss(0)='1'  OR cVar2S17S120P018P016nsss(0)='1'  OR cVar2S18S120P027nsss(0)='1'  OR cVar2S19S120N027P010P032nsss(0)='1'  )then
          oVar1S1085(0) <='1';
          else
          oVar1S1085(0) <='0';
          end if;
        if(cVar2S20S120N027P010P056nsss(0)='1'  OR cVar2S21S120P056P003P029nsss(0)='1'  OR cVar2S22S120N056P012nsss(0)='1'  OR cVar2S23S120N056P012P060nsss(0)='1'  )then
          oVar1S1086(0) <='1';
          else
          oVar1S1086(0) <='0';
          end if;
        if(cVar2S24S120P048nsss(0)='1'  OR cVar2S25S120N048P068P018nsss(0)='1'  OR cVar2S26S120P024P032nsss(0)='1'  OR cVar2S27S120P061P019nsss(0)='1'  )then
          oVar1S1087(0) <='1';
          else
          oVar1S1087(0) <='0';
          end if;
        if(cVar2S28S120P061N019P067nsss(0)='1'  OR cVar2S29S120N061P059P025nsss(0)='1'  OR cVar2S30S120N061P059P064nsss(0)='1'  OR cVar2S31S120P017P019nsss(0)='1'  )then
          oVar1S1088(0) <='1';
          else
          oVar1S1088(0) <='0';
          end if;
        if(cVar2S32S120N017P027nsss(0)='1'  OR cVar2S33S120P017P063P057nsss(0)='1'  OR cVar2S34S120P017P061P055nsss(0)='1'  OR cVar2S35S120P017N061P029nsss(0)='1'  )then
          oVar1S1089(0) <='1';
          else
          oVar1S1089(0) <='0';
          end if;
        if(cVar2S36S120P035P007nsss(0)='1'  OR cVar2S37S120N035P063P011nsss(0)='1'  )then
          oVar1S1090(0) <='1';
          else
          oVar1S1090(0) <='0';
          end if;
        if(cVar2S0S121P056nsss(0)='1'  OR cVar2S1S121N056P008nsss(0)='1'  OR cVar2S2S121N056N008P019nsss(0)='1'  OR cVar2S3S121P056P048P046nsss(0)='1'  )then
          oVar1S1091(0) <='1';
          else
          oVar1S1091(0) <='0';
          end if;
        if(cVar2S4S121P056P015nsss(0)='1'  OR cVar2S5S121P014nsss(0)='1'  OR cVar2S6S121P015P062P050nsss(0)='1'  OR cVar2S7S121P004P025nsss(0)='1'  )then
          oVar1S1092(0) <='1';
          else
          oVar1S1092(0) <='0';
          end if;
        if(cVar2S8S121P004N025P015nsss(0)='1'  OR cVar2S9S121N004P027nsss(0)='1'  OR cVar2S10S121P051P009P055nsss(0)='1'  OR cVar2S11S121P051N009P005nsss(0)='1'  )then
          oVar1S1093(0) <='1';
          else
          oVar1S1093(0) <='0';
          end if;
        if(cVar2S12S121N051P027P008nsss(0)='1'  OR cVar2S13S121P067nsss(0)='1'  OR cVar2S14S121N067P016nsss(0)='1'  OR cVar2S15S121N067N016P048nsss(0)='1'  )then
          oVar1S1094(0) <='1';
          else
          oVar1S1094(0) <='0';
          end if;
        if(cVar2S16S121P048P046P018nsss(0)='1'  OR cVar2S17S121N048P067P037nsss(0)='1'  OR cVar2S18S121N048N067P059nsss(0)='1'  OR cVar2S19S121P015nsss(0)='1'  )then
          oVar1S1095(0) <='1';
          else
          oVar1S1095(0) <='0';
          end if;
        if(cVar2S20S121P066P016nsss(0)='1'  OR cVar2S21S121P066P016P032nsss(0)='1'  OR cVar2S22S121P066P013P012nsss(0)='1'  OR cVar2S23S121P066N013P014nsss(0)='1'  )then
          oVar1S1096(0) <='1';
          else
          oVar1S1096(0) <='0';
          end if;
        if(cVar2S24S121P067P019nsss(0)='1'  OR cVar2S25S121P060P032nsss(0)='1'  OR cVar2S26S121P060N032P007nsss(0)='1'  OR cVar2S27S121N060P032P045nsss(0)='1'  )then
          oVar1S1097(0) <='1';
          else
          oVar1S1097(0) <='0';
          end if;
        if(cVar2S28S121P039nsss(0)='1'  OR cVar2S29S121P062nsss(0)='1'  OR cVar2S30S121N062P018P034nsss(0)='1'  OR cVar2S31S121P063P011nsss(0)='1'  )then
          oVar1S1098(0) <='1';
          else
          oVar1S1098(0) <='0';
          end if;
        if(cVar2S32S121P063N011P053nsss(0)='1'  )then
          oVar1S1099(0) <='1';
          else
          oVar1S1099(0) <='0';
          end if;
        if(cVar1S0S122P052P009P056nsss(0)='1'  OR cVar2S1S122P037nsss(0)='1'  OR cVar2S2S122P050nsss(0)='1'  OR cVar2S3S122N050P019nsss(0)='1'  )then
          oVar1S1100(0) <='1';
          else
          oVar1S1100(0) <='0';
          end if;
        if(cVar2S4S122P061P048P021nsss(0)='1'  OR cVar2S5S122P061P048P017nsss(0)='1'  OR cVar2S6S122P061P059nsss(0)='1'  OR cVar2S7S122P048nsss(0)='1'  )then
          oVar1S1101(0) <='1';
          else
          oVar1S1101(0) <='0';
          end if;
        if(cVar1S8S122P052N009P056P015nsss(0)='1'  OR cVar2S9S122P012nsss(0)='1'  OR cVar2S10S122P004P025nsss(0)='1'  OR cVar2S11S122P004N025P016nsss(0)='1'  )then
          oVar1S1102(0) <='1';
          else
          oVar1S1102(0) <='0';
          end if;
        if(cVar2S12S122N004P027P025nsss(0)='1'  OR cVar2S13S122N004N027P035nsss(0)='1'  OR cVar2S14S122P016nsss(0)='1'  OR cVar1S15S122N052P046P050P006nsss(0)='1'  )then
          oVar1S1103(0) <='1';
          else
          oVar1S1103(0) <='0';
          end if;
        if(cVar2S16S122P041P036P019nsss(0)='1'  OR cVar2S17S122P041N036P035nsss(0)='1'  OR cVar2S18S122P041P005nsss(0)='1'  OR cVar2S19S122P011P036P062nsss(0)='1'  )then
          oVar1S1104(0) <='1';
          else
          oVar1S1104(0) <='0';
          end if;
        if(cVar2S20S122N011P056nsss(0)='1'  OR cVar2S21S122P001P018P059nsss(0)='1'  OR cVar2S22S122P001N018P003nsss(0)='1'  OR cVar2S23S122P007P029P022nsss(0)='1'  )then
          oVar1S1105(0) <='1';
          else
          oVar1S1105(0) <='0';
          end if;
        if(cVar2S0S123P044P015P066nsss(0)='1'  OR cVar2S1S123P044P015P018nsss(0)='1'  OR cVar2S2S123N044P058P007nsss(0)='1'  OR cVar2S3S123N044N058psss(0)='1'  )then
          oVar1S1107(0) <='1';
          else
          oVar1S1107(0) <='0';
          end if;
        if(cVar2S4S123P004nsss(0)='1'  OR cVar2S5S123N004P003nsss(0)='1'  OR cVar2S6S123P065P063nsss(0)='1'  OR cVar2S7S123P065P069P035nsss(0)='1'  )then
          oVar1S1108(0) <='1';
          else
          oVar1S1108(0) <='0';
          end if;
        if(cVar2S8S123P065P069P057nsss(0)='1'  OR cVar2S9S123P030nsss(0)='1'  OR cVar2S10S123N030P015P069nsss(0)='1'  OR cVar2S11S123N030N015P033nsss(0)='1'  )then
          oVar1S1109(0) <='1';
          else
          oVar1S1109(0) <='0';
          end if;
        if(cVar2S12S123P013P032nsss(0)='1'  OR cVar2S13S123P013P011P031nsss(0)='1'  OR cVar2S14S123P013N011P054nsss(0)='1'  OR cVar2S15S123P005nsss(0)='1'  )then
          oVar1S1110(0) <='1';
          else
          oVar1S1110(0) <='0';
          end if;
        if(cVar2S16S123P005P012nsss(0)='1'  OR cVar2S17S123P043nsss(0)='1'  OR cVar2S18S123P064P004P014nsss(0)='1'  OR cVar2S19S123P064N004P007nsss(0)='1'  )then
          oVar1S1111(0) <='1';
          else
          oVar1S1111(0) <='0';
          end if;
        if(cVar2S20S123P064P067nsss(0)='1'  OR cVar2S21S123P064P067P016nsss(0)='1'  OR cVar2S22S123P018P058P067nsss(0)='1'  OR cVar2S23S123P018P058P033nsss(0)='1'  )then
          oVar1S1112(0) <='1';
          else
          oVar1S1112(0) <='0';
          end if;
        if(cVar2S24S123P018P058P015nsss(0)='1'  OR cVar2S25S123P018N058P012nsss(0)='1'  OR cVar2S26S123P011P069nsss(0)='1'  OR cVar2S27S123P011N069P066nsss(0)='1'  )then
          oVar1S1113(0) <='1';
          else
          oVar1S1113(0) <='0';
          end if;
        if(cVar2S28S123N011P056nsss(0)='1'  OR cVar2S29S123N011N056P027nsss(0)='1'  OR cVar2S30S123P062P018nsss(0)='1'  OR cVar2S31S123P015P034nsss(0)='1'  )then
          oVar1S1114(0) <='1';
          else
          oVar1S1114(0) <='0';
          end if;
        if(cVar2S32S123P015N034P066nsss(0)='1'  OR cVar2S33S123P015P014nsss(0)='1'  OR cVar2S34S123P000nsss(0)='1'  OR cVar2S35S123N000P061nsss(0)='1'  )then
          oVar1S1115(0) <='1';
          else
          oVar1S1115(0) <='0';
          end if;
        if(cVar2S36S123N000P061P011nsss(0)='1'  OR cVar2S37S123P010P028nsss(0)='1'  OR cVar2S38S123P010N028P055nsss(0)='1'  OR cVar2S39S123N010P042P016nsss(0)='1'  )then
          oVar1S1116(0) <='1';
          else
          oVar1S1116(0) <='0';
          end if;
        if(cVar2S40S123N010P042P019nsss(0)='1'  OR cVar2S41S123P014P034P035nsss(0)='1'  OR cVar2S42S123P014N034P025nsss(0)='1'  OR cVar2S43S123N014P028nsss(0)='1'  )then
          oVar1S1117(0) <='1';
          else
          oVar1S1117(0) <='0';
          end if;
        if(cVar2S0S124P040P012P023nsss(0)='1'  OR cVar2S1S124P040P012P057nsss(0)='1'  OR cVar2S2S124P040P017nsss(0)='1'  OR cVar2S3S124P042P069P016nsss(0)='1'  )then
          oVar1S1119(0) <='1';
          else
          oVar1S1119(0) <='0';
          end if;
        if(cVar2S4S124N042P023nsss(0)='1'  OR cVar2S5S124P003P066P015nsss(0)='1'  OR cVar2S6S124P003N066P019nsss(0)='1'  OR cVar2S7S124P017P037nsss(0)='1'  )then
          oVar1S1120(0) <='1';
          else
          oVar1S1120(0) <='0';
          end if;
        if(cVar2S8S124P017P037P034nsss(0)='1'  OR cVar2S9S124N017P033P060nsss(0)='1'  OR cVar2S10S124N017N033P060nsss(0)='1'  OR cVar2S11S124P015P019nsss(0)='1'  )then
          oVar1S1121(0) <='1';
          else
          oVar1S1121(0) <='0';
          end if;
        if(cVar2S12S124N015P018P068nsss(0)='1'  OR cVar2S13S124N015P018P014nsss(0)='1'  OR cVar2S14S124P067P017nsss(0)='1'  OR cVar1S15S124N036P017P034P043nsss(0)='1'  )then
          oVar1S1122(0) <='1';
          else
          oVar1S1122(0) <='0';
          end if;
        if(cVar2S16S124P009P058nsss(0)='1'  OR cVar2S17S124P009N058P066nsss(0)='1'  OR cVar2S18S124N009P020P018nsss(0)='1'  OR cVar2S19S124N009N020P029nsss(0)='1'  )then
          oVar1S1123(0) <='1';
          else
          oVar1S1123(0) <='0';
          end if;
        if(cVar2S20S124P010P039nsss(0)='1'  OR cVar2S21S124N010P046P058nsss(0)='1'  OR cVar2S22S124P040nsss(0)='1'  OR cVar2S23S124N040P037P016nsss(0)='1'  )then
          oVar1S1124(0) <='1';
          else
          oVar1S1124(0) <='0';
          end if;
        if(cVar2S24S124P052P005P041nsss(0)='1'  OR cVar2S25S124P052P059P014nsss(0)='1'  OR cVar2S26S124P012P014nsss(0)='1'  OR cVar2S27S124P012P014P054nsss(0)='1'  )then
          oVar1S1125(0) <='1';
          else
          oVar1S1125(0) <='0';
          end if;
        if(cVar2S28S124P040P025nsss(0)='1'  OR cVar2S29S124P040N025P008nsss(0)='1'  OR cVar2S30S124P025P023P034nsss(0)='1'  OR cVar2S31S124P025P047P007nsss(0)='1'  )then
          oVar1S1126(0) <='1';
          else
          oVar1S1126(0) <='0';
          end if;
        if(cVar2S0S125P067P069P068nsss(0)='1'  OR cVar2S1S125P067N069psss(0)='1'  OR cVar2S2S125P067P037nsss(0)='1'  OR cVar2S3S125P036P014nsss(0)='1'  )then
          oVar1S1128(0) <='1';
          else
          oVar1S1128(0) <='0';
          end if;
        if(cVar2S4S125P036N014P018nsss(0)='1'  OR cVar2S5S125P063nsss(0)='1'  OR cVar2S6S125P035P037nsss(0)='1'  OR cVar2S7S125P035N037P052nsss(0)='1'  )then
          oVar1S1129(0) <='1';
          else
          oVar1S1129(0) <='0';
          end if;
        if(cVar2S8S125N035P069nsss(0)='1'  OR cVar2S9S125P052P013P028nsss(0)='1'  OR cVar2S10S125P052N013psss(0)='1'  OR cVar2S11S125P052P050P014nsss(0)='1'  )then
          oVar1S1130(0) <='1';
          else
          oVar1S1130(0) <='0';
          end if;
        if(cVar2S12S125P030P031P012nsss(0)='1'  OR cVar2S13S125N030P004nsss(0)='1'  OR cVar2S14S125N030N004P033nsss(0)='1'  OR cVar2S15S125P067P066nsss(0)='1'  )then
          oVar1S1131(0) <='1';
          else
          oVar1S1131(0) <='0';
          end if;
        if(cVar2S16S125P067P066P016nsss(0)='1'  OR cVar2S17S125N067P065P016nsss(0)='1'  OR cVar2S18S125N067N065P031nsss(0)='1'  OR cVar2S19S125P016P024P068nsss(0)='1'  )then
          oVar1S1132(0) <='1';
          else
          oVar1S1132(0) <='0';
          end if;
        if(cVar2S20S125P016P024P068nsss(0)='1'  OR cVar2S21S125N016P007P033nsss(0)='1'  OR cVar2S22S125P019nsss(0)='1'  OR cVar2S23S125N019P014nsss(0)='1'  )then
          oVar1S1133(0) <='1';
          else
          oVar1S1133(0) <='0';
          end if;
        if(cVar2S24S125P014nsss(0)='1'  OR cVar2S25S125P011P009P030nsss(0)='1'  OR cVar2S26S125P011P019nsss(0)='1'  OR cVar2S27S125P056P015nsss(0)='1'  )then
          oVar1S1134(0) <='1';
          else
          oVar1S1134(0) <='0';
          end if;
        if(cVar2S28S125P056P014nsss(0)='1'  OR cVar2S29S125P017P059nsss(0)='1'  OR cVar2S30S125P017N059P018nsss(0)='1'  OR cVar2S31S125N017P003P063nsss(0)='1'  )then
          oVar1S1135(0) <='1';
          else
          oVar1S1135(0) <='0';
          end if;
        if(cVar2S32S125P008P033P014nsss(0)='1'  OR cVar2S33S125P008N033P011nsss(0)='1'  OR cVar2S34S125P054P013nsss(0)='1'  OR cVar2S35S125N054P057nsss(0)='1'  )then
          oVar1S1136(0) <='1';
          else
          oVar1S1136(0) <='0';
          end if;
        if(cVar2S36S125P056P015nsss(0)='1'  )then
          oVar1S1137(0) <='1';
          else
          oVar1S1137(0) <='0';
          end if;
        if(cVar1S0S126P069P018P026P064nsss(0)='1'  OR cVar2S1S126P019nsss(0)='1'  OR cVar2S2S126N019P012P017nsss(0)='1'  OR cVar2S3S126P008nsss(0)='1'  )then
          oVar1S1138(0) <='1';
          else
          oVar1S1138(0) <='0';
          end if;
        if(cVar2S4S126P067P064nsss(0)='1'  OR cVar2S5S126P067N064P060nsss(0)='1'  OR cVar2S6S126P067P045nsss(0)='1'  OR cVar2S7S126P067N045P014nsss(0)='1'  )then
          oVar1S1139(0) <='1';
          else
          oVar1S1139(0) <='0';
          end if;
        if(cVar2S8S126P062P019nsss(0)='1'  OR cVar2S9S126P062P019P017nsss(0)='1'  OR cVar2S10S126P062P063P014nsss(0)='1'  OR cVar2S11S126P064P063nsss(0)='1'  )then
          oVar1S1140(0) <='1';
          else
          oVar1S1140(0) <='0';
          end if;
        if(cVar2S12S126N064P019P013nsss(0)='1'  OR cVar1S13S126P069P018P068P040nsss(0)='1'  OR cVar2S14S126P063P019nsss(0)='1'  OR cVar2S15S126P063N019P065nsss(0)='1'  )then
          oVar1S1141(0) <='1';
          else
          oVar1S1141(0) <='0';
          end if;
        if(cVar2S16S126N063P033P012nsss(0)='1'  OR cVar2S17S126P014P015nsss(0)='1'  OR cVar2S18S126P014P015P012nsss(0)='1'  OR cVar2S19S126P014P013P047nsss(0)='1'  )then
          oVar1S1142(0) <='1';
          else
          oVar1S1142(0) <='0';
          end if;
        if(cVar2S20S126P045P002nsss(0)='1'  OR cVar2S21S126P043P022nsss(0)='1'  OR cVar2S22S126P043N022P023nsss(0)='1'  OR cVar2S23S126N043P022P031nsss(0)='1'  )then
          oVar1S1143(0) <='1';
          else
          oVar1S1143(0) <='0';
          end if;
        if(cVar2S24S126P068P065P060nsss(0)='1'  OR cVar2S25S126P068P058P062nsss(0)='1'  OR cVar2S26S126P068N058P032nsss(0)='1'  OR cVar2S27S126P062P068P016nsss(0)='1'  )then
          oVar1S1144(0) <='1';
          else
          oVar1S1144(0) <='0';
          end if;
        if(cVar2S28S126P062N068P065nsss(0)='1'  OR cVar2S29S126N062P015P016nsss(0)='1'  OR cVar2S30S126N062N015P006nsss(0)='1'  OR cVar2S31S126P047P007P053nsss(0)='1'  )then
          oVar1S1145(0) <='1';
          else
          oVar1S1145(0) <='0';
          end if;
        if(cVar2S32S126P047P019P024nsss(0)='1'  OR cVar2S33S126P024P019nsss(0)='1'  OR cVar2S34S126P024P019P049nsss(0)='1'  OR cVar2S35S126N024P035P015nsss(0)='1'  )then
          oVar1S1146(0) <='1';
          else
          oVar1S1146(0) <='0';
          end if;
        if(cVar2S36S126N024N035P048nsss(0)='1'  )then
          oVar1S1147(0) <='1';
          else
          oVar1S1147(0) <='0';
          end if;
        if(cVar2S0S127P000nsss(0)='1'  OR cVar2S1S127P000P044P052nsss(0)='1'  OR cVar2S2S127P067P025nsss(0)='1'  OR cVar2S3S127P067P025P010nsss(0)='1'  )then
          oVar1S1148(0) <='1';
          else
          oVar1S1148(0) <='0';
          end if;
        if(cVar2S4S127P067P066P019nsss(0)='1'  OR cVar2S5S127P067N066P026nsss(0)='1'  OR cVar2S6S127P036P051P028nsss(0)='1'  OR cVar2S7S127P036N051P010nsss(0)='1'  )then
          oVar1S1149(0) <='1';
          else
          oVar1S1149(0) <='0';
          end if;
        if(cVar2S8S127P036P030P014nsss(0)='1'  OR cVar2S9S127P026nsss(0)='1'  OR cVar2S10S127N026P067P066nsss(0)='1'  OR cVar2S11S127P007P000P068nsss(0)='1'  )then
          oVar1S1150(0) <='1';
          else
          oVar1S1150(0) <='0';
          end if;
        if(cVar2S12S127P007N000psss(0)='1'  OR cVar2S13S127P007P011nsss(0)='1'  OR cVar2S14S127P005P051nsss(0)='1'  OR cVar2S15S127P008P060nsss(0)='1'  )then
          oVar1S1151(0) <='1';
          else
          oVar1S1151(0) <='0';
          end if;
        if(cVar2S16S127P008N060P014nsss(0)='1'  OR cVar2S17S127N008P052nsss(0)='1'  OR cVar2S18S127N008N052P010nsss(0)='1'  OR cVar2S19S127P053P017P066nsss(0)='1'  )then
          oVar1S1152(0) <='1';
          else
          oVar1S1152(0) <='0';
          end if;
        if(cVar2S20S127P053N017P007nsss(0)='1'  OR cVar2S21S127P053P010nsss(0)='1'  OR cVar2S22S127P015P013nsss(0)='1'  OR cVar2S23S127P015P063P011nsss(0)='1'  )then
          oVar1S1153(0) <='1';
          else
          oVar1S1153(0) <='0';
          end if;
        if(cVar2S24S127P015N063P013nsss(0)='1'  OR cVar2S25S127P063P067P034nsss(0)='1'  OR cVar2S26S127P063P067P017nsss(0)='1'  OR cVar2S27S127P063P019P017nsss(0)='1'  )then
          oVar1S1154(0) <='1';
          else
          oVar1S1154(0) <='0';
          end if;
        if(cVar2S28S127P063N019P017nsss(0)='1'  OR cVar1S29S127P064P018P054P065nsss(0)='1'  OR cVar2S30S127P052nsss(0)='1'  OR cVar2S31S127N052P019P016nsss(0)='1'  )then
          oVar1S1155(0) <='1';
          else
          oVar1S1155(0) <='0';
          end if;
        if(cVar2S32S127P003P015P037nsss(0)='1'  OR cVar2S33S127P003N015P014nsss(0)='1'  OR cVar2S34S127N003P043P004nsss(0)='1'  OR cVar2S35S127P049nsss(0)='1'  )then
          oVar1S1156(0) <='1';
          else
          oVar1S1156(0) <='0';
          end if;
        if(cVar1S36S127P064N018P050P027nsss(0)='1'  OR cVar2S37S127P035P037nsss(0)='1'  OR cVar2S38S127N035P069nsss(0)='1'  )then
          oVar1S1157(0) <='1';
          else
          oVar1S1157(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV4 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar1S0(0)='1'  OR oVar1S1(0)='1'  OR oVar1S2(0)='1'  OR oVar1S3(0)='1'  )then
          oVar2S0(0) <='1';
          else
          oVar2S0(0) <='0';
          end if;
        if(oVar1S4(0)='1'  OR oVar1S5(0)='1'  OR oVar1S6(0)='1'  OR oVar1S7(0)='1'  )then
          oVar2S1(0) <='1';
          else
          oVar2S1(0) <='0';
          end if;
        if(oVar1S8(0)='1'  OR oVar1S9(0)='1'  )then
          oVar2S2(0) <='1';
          else
          oVar2S2(0) <='0';
          end if;
        if(oVar1S10(0)='1'  OR oVar1S11(0)='1'  OR oVar1S12(0)='1'  OR oVar1S13(0)='1'  )then
          oVar2S3(0) <='1';
          else
          oVar2S3(0) <='0';
          end if;
        if(oVar1S14(0)='1'  OR oVar1S15(0)='1'  OR oVar1S16(0)='1'  OR oVar1S17(0)='1'  )then
          oVar2S4(0) <='1';
          else
          oVar2S4(0) <='0';
          end if;
        if(oVar1S19(0)='1'  OR oVar1S20(0)='1'  OR oVar1S21(0)='1'  OR oVar1S22(0)='1'  )then
          oVar2S6(0) <='1';
          else
          oVar2S6(0) <='0';
          end if;
        if(oVar1S23(0)='1'  OR oVar1S24(0)='1'  OR oVar1S25(0)='1'  OR oVar1S26(0)='1'  )then
          oVar2S7(0) <='1';
          else
          oVar2S7(0) <='0';
          end if;
        if(oVar1S27(0)='1'  OR oVar1S28(0)='1'  OR oVar1S29(0)='1'  )then
          oVar2S8(0) <='1';
          else
          oVar2S8(0) <='0';
          end if;
        if(oVar1S30(0)='1'  OR oVar1S31(0)='1'  OR oVar1S32(0)='1'  OR oVar1S33(0)='1'  )then
          oVar2S9(0) <='1';
          else
          oVar2S9(0) <='0';
          end if;
        if(oVar1S34(0)='1'  OR oVar1S35(0)='1'  OR oVar1S36(0)='1'  )then
          oVar2S10(0) <='1';
          else
          oVar2S10(0) <='0';
          end if;
        if(oVar1S38(0)='1'  OR oVar1S39(0)='1'  OR oVar1S40(0)='1'  OR oVar1S41(0)='1'  )then
          oVar2S12(0) <='1';
          else
          oVar2S12(0) <='0';
          end if;
        if(oVar1S42(0)='1'  OR oVar1S43(0)='1'  OR oVar1S44(0)='1'  OR oVar1S45(0)='1'  )then
          oVar2S13(0) <='1';
          else
          oVar2S13(0) <='0';
          end if;
        if(oVar1S46(0)='1'  OR oVar1S47(0)='1'  OR oVar1S48(0)='1'  OR oVar1S49(0)='1'  )then
          oVar2S15(0) <='1';
          else
          oVar2S15(0) <='0';
          end if;
        if(oVar1S50(0)='1'  OR oVar1S51(0)='1'  OR oVar1S52(0)='1'  OR oVar1S53(0)='1'  )then
          oVar2S16(0) <='1';
          else
          oVar2S16(0) <='0';
          end if;
        if(oVar1S54(0)='1'  )then
          oVar2S17(0) <='1';
          else
          oVar2S17(0) <='0';
          end if;
        if(oVar1S55(0)='1'  OR oVar1S56(0)='1'  OR oVar1S57(0)='1'  OR oVar1S58(0)='1'  )then
          oVar2S18(0) <='1';
          else
          oVar2S18(0) <='0';
          end if;
        if(oVar1S59(0)='1'  OR oVar1S60(0)='1'  OR oVar1S61(0)='1'  )then
          oVar2S19(0) <='1';
          else
          oVar2S19(0) <='0';
          end if;
        if(oVar1S62(0)='1'  OR oVar1S63(0)='1'  OR oVar1S64(0)='1'  OR oVar1S65(0)='1'  )then
          oVar2S20(0) <='1';
          else
          oVar2S20(0) <='0';
          end if;
        if(oVar1S66(0)='1'  OR oVar1S67(0)='1'  OR oVar1S68(0)='1'  OR oVar1S69(0)='1'  )then
          oVar2S21(0) <='1';
          else
          oVar2S21(0) <='0';
          end if;
        if(oVar1S70(0)='1'  OR oVar1S71(0)='1'  OR oVar1S72(0)='1'  OR oVar1S73(0)='1'  )then
          oVar2S23(0) <='1';
          else
          oVar2S23(0) <='0';
          end if;
        if(oVar1S74(0)='1'  OR oVar1S75(0)='1'  OR oVar1S76(0)='1'  )then
          oVar2S24(0) <='1';
          else
          oVar2S24(0) <='0';
          end if;
        if(oVar1S77(0)='1'  OR oVar1S78(0)='1'  OR oVar1S79(0)='1'  OR oVar1S80(0)='1'  )then
          oVar2S25(0) <='1';
          else
          oVar2S25(0) <='0';
          end if;
        if(oVar1S81(0)='1'  OR oVar1S82(0)='1'  OR oVar1S83(0)='1'  OR oVar1S84(0)='1'  )then
          oVar2S26(0) <='1';
          else
          oVar2S26(0) <='0';
          end if;
        if(oVar1S85(0)='1'  )then
          oVar2S27(0) <='1';
          else
          oVar2S27(0) <='0';
          end if;
        if(oVar1S87(0)='1'  OR oVar1S88(0)='1'  OR oVar1S89(0)='1'  OR oVar1S90(0)='1'  )then
          oVar2S28(0) <='1';
          else
          oVar2S28(0) <='0';
          end if;
        if(oVar1S91(0)='1'  OR oVar1S92(0)='1'  OR oVar1S93(0)='1'  OR oVar1S94(0)='1'  )then
          oVar2S29(0) <='1';
          else
          oVar2S29(0) <='0';
          end if;
        if(oVar1S95(0)='1'  )then
          oVar2S30(0) <='1';
          else
          oVar2S30(0) <='0';
          end if;
        if(oVar1S97(0)='1'  OR oVar1S98(0)='1'  OR oVar1S99(0)='1'  OR oVar1S100(0)='1'  )then
          oVar2S31(0) <='1';
          else
          oVar2S31(0) <='0';
          end if;
        if(oVar1S101(0)='1'  OR oVar1S102(0)='1'  )then
          oVar2S32(0) <='1';
          else
          oVar2S32(0) <='0';
          end if;
        if(oVar1S104(0)='1'  OR oVar1S105(0)='1'  OR oVar1S106(0)='1'  OR oVar1S107(0)='1'  )then
          oVar2S33(0) <='1';
          else
          oVar2S33(0) <='0';
          end if;
        if(oVar1S108(0)='1'  OR oVar1S109(0)='1'  OR oVar1S110(0)='1'  OR oVar1S111(0)='1'  )then
          oVar2S34(0) <='1';
          else
          oVar2S34(0) <='0';
          end if;
        if(oVar1S112(0)='1'  OR oVar1S113(0)='1'  )then
          oVar2S35(0) <='1';
          else
          oVar2S35(0) <='0';
          end if;
        if(oVar1S114(0)='1'  OR oVar1S115(0)='1'  OR oVar1S116(0)='1'  OR oVar1S117(0)='1'  )then
          oVar2S36(0) <='1';
          else
          oVar2S36(0) <='0';
          end if;
        if(oVar1S118(0)='1'  OR oVar1S119(0)='1'  OR oVar1S120(0)='1'  OR oVar1S121(0)='1'  )then
          oVar2S37(0) <='1';
          else
          oVar2S37(0) <='0';
          end if;
        if(oVar1S122(0)='1'  OR oVar1S123(0)='1'  )then
          oVar2S38(0) <='1';
          else
          oVar2S38(0) <='0';
          end if;
        if(oVar1S124(0)='1'  OR oVar1S125(0)='1'  OR oVar1S126(0)='1'  OR oVar1S127(0)='1'  )then
          oVar2S39(0) <='1';
          else
          oVar2S39(0) <='0';
          end if;
        if(oVar1S128(0)='1'  OR oVar1S129(0)='1'  OR oVar1S130(0)='1'  OR oVar1S131(0)='1'  )then
          oVar2S40(0) <='1';
          else
          oVar2S40(0) <='0';
          end if;
        if(oVar1S132(0)='1'  )then
          oVar2S41(0) <='1';
          else
          oVar2S41(0) <='0';
          end if;
        if(oVar1S133(0)='1'  OR oVar1S134(0)='1'  OR oVar1S135(0)='1'  OR oVar1S136(0)='1'  )then
          oVar2S42(0) <='1';
          else
          oVar2S42(0) <='0';
          end if;
        if(oVar1S137(0)='1'  OR oVar1S138(0)='1'  OR oVar1S139(0)='1'  OR oVar1S140(0)='1'  )then
          oVar2S43(0) <='1';
          else
          oVar2S43(0) <='0';
          end if;
        if(oVar1S141(0)='1'  OR oVar1S142(0)='1'  OR oVar1S143(0)='1'  OR oVar1S144(0)='1'  )then
          oVar2S45(0) <='1';
          else
          oVar2S45(0) <='0';
          end if;
        if(oVar1S145(0)='1'  OR oVar1S146(0)='1'  OR oVar1S147(0)='1'  OR oVar1S148(0)='1'  )then
          oVar2S46(0) <='1';
          else
          oVar2S46(0) <='0';
          end if;
        if(oVar1S150(0)='1'  OR oVar1S151(0)='1'  OR oVar1S152(0)='1'  OR oVar1S153(0)='1'  )then
          oVar2S48(0) <='1';
          else
          oVar2S48(0) <='0';
          end if;
        if(oVar1S154(0)='1'  OR oVar1S155(0)='1'  OR oVar1S156(0)='1'  OR oVar1S157(0)='1'  )then
          oVar2S49(0) <='1';
          else
          oVar2S49(0) <='0';
          end if;
        if(oVar1S158(0)='1'  )then
          oVar2S50(0) <='1';
          else
          oVar2S50(0) <='0';
          end if;
        if(oVar1S159(0)='1'  OR oVar1S160(0)='1'  OR oVar1S161(0)='1'  OR oVar1S162(0)='1'  )then
          oVar2S51(0) <='1';
          else
          oVar2S51(0) <='0';
          end if;
        if(oVar1S163(0)='1'  OR oVar1S164(0)='1'  OR oVar1S165(0)='1'  OR oVar1S166(0)='1'  )then
          oVar2S52(0) <='1';
          else
          oVar2S52(0) <='0';
          end if;
        if(oVar1S167(0)='1'  )then
          oVar2S53(0) <='1';
          else
          oVar2S53(0) <='0';
          end if;
        if(oVar1S168(0)='1'  OR oVar1S169(0)='1'  OR oVar1S170(0)='1'  OR oVar1S171(0)='1'  )then
          oVar2S54(0) <='1';
          else
          oVar2S54(0) <='0';
          end if;
        if(oVar1S172(0)='1'  OR oVar1S173(0)='1'  OR oVar1S174(0)='1'  OR oVar1S175(0)='1'  )then
          oVar2S55(0) <='1';
          else
          oVar2S55(0) <='0';
          end if;
        if(oVar1S176(0)='1'  OR oVar1S177(0)='1'  )then
          oVar2S56(0) <='1';
          else
          oVar2S56(0) <='0';
          end if;
        if(oVar1S178(0)='1'  OR oVar1S179(0)='1'  OR oVar1S180(0)='1'  OR oVar1S181(0)='1'  )then
          oVar2S57(0) <='1';
          else
          oVar2S57(0) <='0';
          end if;
        if(oVar1S182(0)='1'  OR oVar1S183(0)='1'  OR oVar1S184(0)='1'  OR oVar1S185(0)='1'  )then
          oVar2S58(0) <='1';
          else
          oVar2S58(0) <='0';
          end if;
        if(oVar1S186(0)='1'  )then
          oVar2S59(0) <='1';
          else
          oVar2S59(0) <='0';
          end if;
        if(oVar1S187(0)='1'  OR oVar1S188(0)='1'  OR oVar1S189(0)='1'  OR oVar1S190(0)='1'  )then
          oVar2S60(0) <='1';
          else
          oVar2S60(0) <='0';
          end if;
        if(oVar1S191(0)='1'  OR oVar1S192(0)='1'  OR oVar1S193(0)='1'  OR oVar1S194(0)='1'  )then
          oVar2S61(0) <='1';
          else
          oVar2S61(0) <='0';
          end if;
        if(oVar1S195(0)='1'  )then
          oVar2S62(0) <='1';
          else
          oVar2S62(0) <='0';
          end if;
        if(oVar1S196(0)='1'  OR oVar1S197(0)='1'  OR oVar1S198(0)='1'  OR oVar1S199(0)='1'  )then
          oVar2S63(0) <='1';
          else
          oVar2S63(0) <='0';
          end if;
        if(oVar1S200(0)='1'  OR oVar1S201(0)='1'  OR oVar1S202(0)='1'  OR oVar1S203(0)='1'  )then
          oVar2S64(0) <='1';
          else
          oVar2S64(0) <='0';
          end if;
        if(oVar1S204(0)='1'  OR oVar1S205(0)='1'  OR oVar1S206(0)='1'  OR oVar1S207(0)='1'  )then
          oVar2S66(0) <='1';
          else
          oVar2S66(0) <='0';
          end if;
        if(oVar1S208(0)='1'  OR oVar1S209(0)='1'  )then
          oVar2S67(0) <='1';
          else
          oVar2S67(0) <='0';
          end if;
        if(oVar1S210(0)='1'  OR oVar1S211(0)='1'  OR oVar1S212(0)='1'  OR oVar1S213(0)='1'  )then
          oVar2S68(0) <='1';
          else
          oVar2S68(0) <='0';
          end if;
        if(oVar1S214(0)='1'  OR oVar1S215(0)='1'  OR oVar1S216(0)='1'  OR oVar1S217(0)='1'  )then
          oVar2S69(0) <='1';
          else
          oVar2S69(0) <='0';
          end if;
        if(oVar1S218(0)='1'  OR oVar1S219(0)='1'  OR oVar1S220(0)='1'  OR oVar1S221(0)='1'  )then
          oVar2S71(0) <='1';
          else
          oVar2S71(0) <='0';
          end if;
        if(oVar1S222(0)='1'  OR oVar1S223(0)='1'  OR oVar1S224(0)='1'  OR oVar1S225(0)='1'  )then
          oVar2S72(0) <='1';
          else
          oVar2S72(0) <='0';
          end if;
        if(oVar1S226(0)='1'  OR oVar1S227(0)='1'  OR oVar1S228(0)='1'  OR oVar1S229(0)='1'  )then
          oVar2S74(0) <='1';
          else
          oVar2S74(0) <='0';
          end if;
        if(oVar1S230(0)='1'  OR oVar1S231(0)='1'  OR oVar1S232(0)='1'  OR oVar1S233(0)='1'  )then
          oVar2S75(0) <='1';
          else
          oVar2S75(0) <='0';
          end if;
        if(oVar1S234(0)='1'  OR oVar1S235(0)='1'  OR oVar1S236(0)='1'  )then
          oVar2S76(0) <='1';
          else
          oVar2S76(0) <='0';
          end if;
        if(oVar1S237(0)='1'  OR oVar1S238(0)='1'  OR oVar1S239(0)='1'  OR oVar1S240(0)='1'  )then
          oVar2S77(0) <='1';
          else
          oVar2S77(0) <='0';
          end if;
        if(oVar1S241(0)='1'  OR oVar1S242(0)='1'  )then
          oVar2S78(0) <='1';
          else
          oVar2S78(0) <='0';
          end if;
        if(oVar1S244(0)='1'  OR oVar1S245(0)='1'  OR oVar1S246(0)='1'  OR oVar1S247(0)='1'  )then
          oVar2S79(0) <='1';
          else
          oVar2S79(0) <='0';
          end if;
        if(oVar1S248(0)='1'  OR oVar1S249(0)='1'  OR oVar1S250(0)='1'  )then
          oVar2S80(0) <='1';
          else
          oVar2S80(0) <='0';
          end if;
        if(oVar1S251(0)='1'  OR oVar1S252(0)='1'  OR oVar1S253(0)='1'  OR oVar1S254(0)='1'  )then
          oVar2S81(0) <='1';
          else
          oVar2S81(0) <='0';
          end if;
        if(oVar1S255(0)='1'  OR oVar1S256(0)='1'  )then
          oVar2S82(0) <='1';
          else
          oVar2S82(0) <='0';
          end if;
        if(oVar1S257(0)='1'  OR oVar1S258(0)='1'  OR oVar1S259(0)='1'  OR oVar1S260(0)='1'  )then
          oVar2S83(0) <='1';
          else
          oVar2S83(0) <='0';
          end if;
        if(oVar1S261(0)='1'  OR oVar1S262(0)='1'  OR oVar1S263(0)='1'  OR oVar1S264(0)='1'  )then
          oVar2S84(0) <='1';
          else
          oVar2S84(0) <='0';
          end if;
        if(oVar1S265(0)='1'  OR oVar1S266(0)='1'  )then
          oVar2S85(0) <='1';
          else
          oVar2S85(0) <='0';
          end if;
        if(oVar1S267(0)='1'  OR oVar1S268(0)='1'  OR oVar1S269(0)='1'  OR oVar1S270(0)='1'  )then
          oVar2S86(0) <='1';
          else
          oVar2S86(0) <='0';
          end if;
        if(oVar1S271(0)='1'  OR oVar1S272(0)='1'  OR oVar1S273(0)='1'  OR oVar1S274(0)='1'  )then
          oVar2S87(0) <='1';
          else
          oVar2S87(0) <='0';
          end if;
        if(oVar1S275(0)='1'  OR oVar1S276(0)='1'  OR oVar1S277(0)='1'  )then
          oVar2S88(0) <='1';
          else
          oVar2S88(0) <='0';
          end if;
        if(oVar1S279(0)='1'  OR oVar1S280(0)='1'  OR oVar1S281(0)='1'  OR oVar1S282(0)='1'  )then
          oVar2S90(0) <='1';
          else
          oVar2S90(0) <='0';
          end if;
        if(oVar1S283(0)='1'  OR oVar1S284(0)='1'  OR oVar1S285(0)='1'  OR oVar1S286(0)='1'  )then
          oVar2S91(0) <='1';
          else
          oVar2S91(0) <='0';
          end if;
        if(oVar1S287(0)='1'  )then
          oVar2S92(0) <='1';
          else
          oVar2S92(0) <='0';
          end if;
        if(oVar1S288(0)='1'  OR oVar1S289(0)='1'  OR oVar1S290(0)='1'  OR oVar1S291(0)='1'  )then
          oVar2S93(0) <='1';
          else
          oVar2S93(0) <='0';
          end if;
        if(oVar1S292(0)='1'  OR oVar1S293(0)='1'  OR oVar1S294(0)='1'  OR oVar1S295(0)='1'  )then
          oVar2S94(0) <='1';
          else
          oVar2S94(0) <='0';
          end if;
        if(oVar1S297(0)='1'  OR oVar1S298(0)='1'  OR oVar1S299(0)='1'  OR oVar1S300(0)='1'  )then
          oVar2S96(0) <='1';
          else
          oVar2S96(0) <='0';
          end if;
        if(oVar1S301(0)='1'  OR oVar1S302(0)='1'  OR oVar1S303(0)='1'  OR oVar1S304(0)='1'  )then
          oVar2S97(0) <='1';
          else
          oVar2S97(0) <='0';
          end if;
        if(oVar1S305(0)='1'  OR oVar1S306(0)='1'  OR oVar1S307(0)='1'  OR oVar1S308(0)='1'  )then
          oVar2S98(0) <='1';
          else
          oVar2S98(0) <='0';
          end if;
        if(oVar1S309(0)='1'  OR oVar1S310(0)='1'  OR oVar1S311(0)='1'  OR oVar1S312(0)='1'  )then
          oVar2S100(0) <='1';
          else
          oVar2S100(0) <='0';
          end if;
        if(oVar1S313(0)='1'  OR oVar1S314(0)='1'  OR oVar1S315(0)='1'  )then
          oVar2S101(0) <='1';
          else
          oVar2S101(0) <='0';
          end if;
        if(oVar1S317(0)='1'  OR oVar1S318(0)='1'  OR oVar1S319(0)='1'  OR oVar1S320(0)='1'  )then
          oVar2S103(0) <='1';
          else
          oVar2S103(0) <='0';
          end if;
        if(oVar1S321(0)='1'  OR oVar1S322(0)='1'  OR oVar1S323(0)='1'  OR oVar1S324(0)='1'  )then
          oVar2S104(0) <='1';
          else
          oVar2S104(0) <='0';
          end if;
        if(oVar1S325(0)='1'  )then
          oVar2S105(0) <='1';
          else
          oVar2S105(0) <='0';
          end if;
        if(oVar1S326(0)='1'  OR oVar1S327(0)='1'  OR oVar1S328(0)='1'  OR oVar1S329(0)='1'  )then
          oVar2S106(0) <='1';
          else
          oVar2S106(0) <='0';
          end if;
        if(oVar1S330(0)='1'  OR oVar1S331(0)='1'  OR oVar1S332(0)='1'  OR oVar1S333(0)='1'  )then
          oVar2S107(0) <='1';
          else
          oVar2S107(0) <='0';
          end if;
        if(oVar1S334(0)='1'  )then
          oVar2S108(0) <='1';
          else
          oVar2S108(0) <='0';
          end if;
        if(oVar1S335(0)='1'  OR oVar1S336(0)='1'  OR oVar1S337(0)='1'  OR oVar1S338(0)='1'  )then
          oVar2S109(0) <='1';
          else
          oVar2S109(0) <='0';
          end if;
        if(oVar1S339(0)='1'  OR oVar1S340(0)='1'  OR oVar1S341(0)='1'  OR oVar1S342(0)='1'  )then
          oVar2S110(0) <='1';
          else
          oVar2S110(0) <='0';
          end if;
        if(oVar1S343(0)='1'  OR oVar1S344(0)='1'  )then
          oVar2S111(0) <='1';
          else
          oVar2S111(0) <='0';
          end if;
        if(oVar1S345(0)='1'  OR oVar1S346(0)='1'  OR oVar1S347(0)='1'  OR oVar1S348(0)='1'  )then
          oVar2S112(0) <='1';
          else
          oVar2S112(0) <='0';
          end if;
        if(oVar1S349(0)='1'  OR oVar1S350(0)='1'  OR oVar1S351(0)='1'  OR oVar1S352(0)='1'  )then
          oVar2S113(0) <='1';
          else
          oVar2S113(0) <='0';
          end if;
        if(oVar1S353(0)='1'  OR oVar1S354(0)='1'  OR oVar1S355(0)='1'  )then
          oVar2S114(0) <='1';
          else
          oVar2S114(0) <='0';
          end if;
        if(oVar1S356(0)='1'  OR oVar1S357(0)='1'  OR oVar1S358(0)='1'  OR oVar1S359(0)='1'  )then
          oVar2S115(0) <='1';
          else
          oVar2S115(0) <='0';
          end if;
        if(oVar1S360(0)='1'  OR oVar1S361(0)='1'  OR oVar1S362(0)='1'  OR oVar1S363(0)='1'  )then
          oVar2S116(0) <='1';
          else
          oVar2S116(0) <='0';
          end if;
        if(oVar1S364(0)='1'  OR oVar1S365(0)='1'  )then
          oVar2S117(0) <='1';
          else
          oVar2S117(0) <='0';
          end if;
        if(oVar1S366(0)='1'  OR oVar1S367(0)='1'  OR oVar1S368(0)='1'  OR oVar1S369(0)='1'  )then
          oVar2S118(0) <='1';
          else
          oVar2S118(0) <='0';
          end if;
        if(oVar1S370(0)='1'  OR oVar1S371(0)='1'  OR oVar1S372(0)='1'  OR oVar1S373(0)='1'  )then
          oVar2S119(0) <='1';
          else
          oVar2S119(0) <='0';
          end if;
        if(oVar1S374(0)='1'  OR oVar1S375(0)='1'  OR oVar1S376(0)='1'  OR oVar1S377(0)='1'  )then
          oVar2S121(0) <='1';
          else
          oVar2S121(0) <='0';
          end if;
        if(oVar1S378(0)='1'  OR oVar1S379(0)='1'  OR oVar1S380(0)='1'  OR oVar1S381(0)='1'  )then
          oVar2S122(0) <='1';
          else
          oVar2S122(0) <='0';
          end if;
        if(oVar1S382(0)='1'  OR oVar1S383(0)='1'  )then
          oVar2S123(0) <='1';
          else
          oVar2S123(0) <='0';
          end if;
        if(oVar1S384(0)='1'  OR oVar1S385(0)='1'  OR oVar1S386(0)='1'  OR oVar1S387(0)='1'  )then
          oVar2S124(0) <='1';
          else
          oVar2S124(0) <='0';
          end if;
        if(oVar1S388(0)='1'  OR oVar1S389(0)='1'  OR oVar1S390(0)='1'  OR oVar1S391(0)='1'  )then
          oVar2S125(0) <='1';
          else
          oVar2S125(0) <='0';
          end if;
        if(oVar1S392(0)='1'  )then
          oVar2S126(0) <='1';
          else
          oVar2S126(0) <='0';
          end if;
        if(oVar1S393(0)='1'  OR oVar1S394(0)='1'  OR oVar1S395(0)='1'  OR oVar1S396(0)='1'  )then
          oVar2S127(0) <='1';
          else
          oVar2S127(0) <='0';
          end if;
        if(oVar1S397(0)='1'  OR oVar1S398(0)='1'  OR oVar1S399(0)='1'  )then
          oVar2S128(0) <='1';
          else
          oVar2S128(0) <='0';
          end if;
        if(oVar1S400(0)='1'  OR oVar1S401(0)='1'  OR oVar1S402(0)='1'  OR oVar1S403(0)='1'  )then
          oVar2S129(0) <='1';
          else
          oVar2S129(0) <='0';
          end if;
        if(oVar1S404(0)='1'  OR oVar1S405(0)='1'  OR oVar1S406(0)='1'  OR oVar1S407(0)='1'  )then
          oVar2S130(0) <='1';
          else
          oVar2S130(0) <='0';
          end if;
        if(oVar1S408(0)='1'  OR oVar1S409(0)='1'  OR oVar1S410(0)='1'  OR oVar1S411(0)='1'  )then
          oVar2S132(0) <='1';
          else
          oVar2S132(0) <='0';
          end if;
        if(oVar1S412(0)='1'  OR oVar1S413(0)='1'  OR oVar1S414(0)='1'  OR oVar1S415(0)='1'  )then
          oVar2S133(0) <='1';
          else
          oVar2S133(0) <='0';
          end if;
        if(oVar1S416(0)='1'  )then
          oVar2S134(0) <='1';
          else
          oVar2S134(0) <='0';
          end if;
        if(oVar1S417(0)='1'  OR oVar1S418(0)='1'  OR oVar1S419(0)='1'  OR oVar1S420(0)='1'  )then
          oVar2S135(0) <='1';
          else
          oVar2S135(0) <='0';
          end if;
        if(oVar1S421(0)='1'  OR oVar1S422(0)='1'  OR oVar1S423(0)='1'  OR oVar1S424(0)='1'  )then
          oVar2S136(0) <='1';
          else
          oVar2S136(0) <='0';
          end if;
        if(oVar1S425(0)='1'  )then
          oVar2S137(0) <='1';
          else
          oVar2S137(0) <='0';
          end if;
        if(oVar1S426(0)='1'  OR oVar1S427(0)='1'  OR oVar1S428(0)='1'  OR oVar1S429(0)='1'  )then
          oVar2S138(0) <='1';
          else
          oVar2S138(0) <='0';
          end if;
        if(oVar1S430(0)='1'  OR oVar1S431(0)='1'  OR oVar1S432(0)='1'  )then
          oVar2S139(0) <='1';
          else
          oVar2S139(0) <='0';
          end if;
        if(oVar1S434(0)='1'  OR oVar1S435(0)='1'  OR oVar1S436(0)='1'  OR oVar1S437(0)='1'  )then
          oVar2S141(0) <='1';
          else
          oVar2S141(0) <='0';
          end if;
        if(oVar1S438(0)='1'  OR oVar1S439(0)='1'  OR oVar1S440(0)='1'  OR oVar1S441(0)='1'  )then
          oVar2S142(0) <='1';
          else
          oVar2S142(0) <='0';
          end if;
        if(oVar1S442(0)='1'  OR oVar1S443(0)='1'  OR oVar1S444(0)='1'  OR oVar1S445(0)='1'  )then
          oVar2S144(0) <='1';
          else
          oVar2S144(0) <='0';
          end if;
        if(oVar1S446(0)='1'  OR oVar1S447(0)='1'  OR oVar1S448(0)='1'  OR oVar1S449(0)='1'  )then
          oVar2S145(0) <='1';
          else
          oVar2S145(0) <='0';
          end if;
        if(oVar1S450(0)='1'  )then
          oVar2S146(0) <='1';
          else
          oVar2S146(0) <='0';
          end if;
        if(oVar1S451(0)='1'  OR oVar1S452(0)='1'  OR oVar1S453(0)='1'  OR oVar1S454(0)='1'  )then
          oVar2S147(0) <='1';
          else
          oVar2S147(0) <='0';
          end if;
        if(oVar1S455(0)='1'  OR oVar1S456(0)='1'  OR oVar1S457(0)='1'  OR oVar1S458(0)='1'  )then
          oVar2S148(0) <='1';
          else
          oVar2S148(0) <='0';
          end if;
        if(oVar1S460(0)='1'  OR oVar1S461(0)='1'  OR oVar1S462(0)='1'  OR oVar1S463(0)='1'  )then
          oVar2S150(0) <='1';
          else
          oVar2S150(0) <='0';
          end if;
        if(oVar1S464(0)='1'  OR oVar1S465(0)='1'  OR oVar1S466(0)='1'  )then
          oVar2S151(0) <='1';
          else
          oVar2S151(0) <='0';
          end if;
        if(oVar1S468(0)='1'  OR oVar1S469(0)='1'  OR oVar1S470(0)='1'  OR oVar1S471(0)='1'  )then
          oVar2S153(0) <='1';
          else
          oVar2S153(0) <='0';
          end if;
        if(oVar1S472(0)='1'  OR oVar1S473(0)='1'  OR oVar1S474(0)='1'  OR oVar1S475(0)='1'  )then
          oVar2S154(0) <='1';
          else
          oVar2S154(0) <='0';
          end if;
        if(oVar1S476(0)='1'  OR oVar1S477(0)='1'  )then
          oVar2S155(0) <='1';
          else
          oVar2S155(0) <='0';
          end if;
        if(oVar1S478(0)='1'  OR oVar1S479(0)='1'  OR oVar1S480(0)='1'  OR oVar1S481(0)='1'  )then
          oVar2S156(0) <='1';
          else
          oVar2S156(0) <='0';
          end if;
        if(oVar1S482(0)='1'  OR oVar1S483(0)='1'  OR oVar1S484(0)='1'  OR oVar1S485(0)='1'  )then
          oVar2S157(0) <='1';
          else
          oVar2S157(0) <='0';
          end if;
        if(oVar1S486(0)='1'  )then
          oVar2S158(0) <='1';
          else
          oVar2S158(0) <='0';
          end if;
        if(oVar1S488(0)='1'  OR oVar1S489(0)='1'  OR oVar1S490(0)='1'  OR oVar1S491(0)='1'  )then
          oVar2S159(0) <='1';
          else
          oVar2S159(0) <='0';
          end if;
        if(oVar1S492(0)='1'  OR oVar1S493(0)='1'  OR oVar1S494(0)='1'  OR oVar1S495(0)='1'  )then
          oVar2S160(0) <='1';
          else
          oVar2S160(0) <='0';
          end if;
        if(oVar1S497(0)='1'  OR oVar1S498(0)='1'  OR oVar1S499(0)='1'  OR oVar1S500(0)='1'  )then
          oVar2S162(0) <='1';
          else
          oVar2S162(0) <='0';
          end if;
        if(oVar1S501(0)='1'  OR oVar1S502(0)='1'  OR oVar1S503(0)='1'  OR oVar1S504(0)='1'  )then
          oVar2S163(0) <='1';
          else
          oVar2S163(0) <='0';
          end if;
        if(oVar1S505(0)='1'  OR oVar1S506(0)='1'  OR oVar1S507(0)='1'  OR oVar1S508(0)='1'  )then
          oVar2S165(0) <='1';
          else
          oVar2S165(0) <='0';
          end if;
        if(oVar1S509(0)='1'  OR oVar1S510(0)='1'  OR oVar1S511(0)='1'  OR oVar1S512(0)='1'  )then
          oVar2S166(0) <='1';
          else
          oVar2S166(0) <='0';
          end if;
        if(oVar1S513(0)='1'  OR oVar1S514(0)='1'  OR oVar1S515(0)='1'  OR oVar1S516(0)='1'  )then
          oVar2S168(0) <='1';
          else
          oVar2S168(0) <='0';
          end if;
        if(oVar1S517(0)='1'  OR oVar1S518(0)='1'  OR oVar1S519(0)='1'  OR oVar1S520(0)='1'  )then
          oVar2S169(0) <='1';
          else
          oVar2S169(0) <='0';
          end if;
        if(oVar1S521(0)='1'  OR oVar1S522(0)='1'  )then
          oVar2S170(0) <='1';
          else
          oVar2S170(0) <='0';
          end if;
        if(oVar1S523(0)='1'  OR oVar1S524(0)='1'  OR oVar1S525(0)='1'  OR oVar1S526(0)='1'  )then
          oVar2S171(0) <='1';
          else
          oVar2S171(0) <='0';
          end if;
        if(oVar1S527(0)='1'  OR oVar1S528(0)='1'  OR oVar1S529(0)='1'  )then
          oVar2S172(0) <='1';
          else
          oVar2S172(0) <='0';
          end if;
        if(oVar1S530(0)='1'  OR oVar1S531(0)='1'  OR oVar1S532(0)='1'  OR oVar1S533(0)='1'  )then
          oVar2S173(0) <='1';
          else
          oVar2S173(0) <='0';
          end if;
        if(oVar1S534(0)='1'  OR oVar1S535(0)='1'  OR oVar1S536(0)='1'  OR oVar1S537(0)='1'  )then
          oVar2S174(0) <='1';
          else
          oVar2S174(0) <='0';
          end if;
        if(oVar1S538(0)='1'  OR oVar1S539(0)='1'  )then
          oVar2S175(0) <='1';
          else
          oVar2S175(0) <='0';
          end if;
        if(oVar1S540(0)='1'  OR oVar1S541(0)='1'  OR oVar1S542(0)='1'  OR oVar1S543(0)='1'  )then
          oVar2S176(0) <='1';
          else
          oVar2S176(0) <='0';
          end if;
        if(oVar1S544(0)='1'  OR oVar1S545(0)='1'  OR oVar1S546(0)='1'  OR oVar1S547(0)='1'  )then
          oVar2S177(0) <='1';
          else
          oVar2S177(0) <='0';
          end if;
        if(oVar1S548(0)='1'  )then
          oVar2S178(0) <='1';
          else
          oVar2S178(0) <='0';
          end if;
        if(oVar1S549(0)='1'  OR oVar1S550(0)='1'  OR oVar1S551(0)='1'  OR oVar1S552(0)='1'  )then
          oVar2S179(0) <='1';
          else
          oVar2S179(0) <='0';
          end if;
        if(oVar1S553(0)='1'  OR oVar1S554(0)='1'  OR oVar1S555(0)='1'  OR oVar1S556(0)='1'  )then
          oVar2S180(0) <='1';
          else
          oVar2S180(0) <='0';
          end if;
        if(oVar1S557(0)='1'  OR oVar1S558(0)='1'  )then
          oVar2S181(0) <='1';
          else
          oVar2S181(0) <='0';
          end if;
        if(oVar1S559(0)='1'  OR oVar1S560(0)='1'  OR oVar1S561(0)='1'  OR oVar1S562(0)='1'  )then
          oVar2S182(0) <='1';
          else
          oVar2S182(0) <='0';
          end if;
        if(oVar1S563(0)='1'  OR oVar1S564(0)='1'  OR oVar1S565(0)='1'  OR oVar1S566(0)='1'  )then
          oVar2S183(0) <='1';
          else
          oVar2S183(0) <='0';
          end if;
        if(oVar1S568(0)='1'  OR oVar1S569(0)='1'  OR oVar1S570(0)='1'  OR oVar1S571(0)='1'  )then
          oVar2S185(0) <='1';
          else
          oVar2S185(0) <='0';
          end if;
        if(oVar1S572(0)='1'  OR oVar1S573(0)='1'  )then
          oVar2S186(0) <='1';
          else
          oVar2S186(0) <='0';
          end if;
        if(oVar1S574(0)='1'  OR oVar1S575(0)='1'  OR oVar1S576(0)='1'  OR oVar1S577(0)='1'  )then
          oVar2S187(0) <='1';
          else
          oVar2S187(0) <='0';
          end if;
        if(oVar1S578(0)='1'  OR oVar1S579(0)='1'  OR oVar1S580(0)='1'  )then
          oVar2S188(0) <='1';
          else
          oVar2S188(0) <='0';
          end if;
        if(oVar1S582(0)='1'  OR oVar1S583(0)='1'  OR oVar1S584(0)='1'  OR oVar1S585(0)='1'  )then
          oVar2S190(0) <='1';
          else
          oVar2S190(0) <='0';
          end if;
        if(oVar1S586(0)='1'  OR oVar1S587(0)='1'  OR oVar1S588(0)='1'  OR oVar1S589(0)='1'  )then
          oVar2S191(0) <='1';
          else
          oVar2S191(0) <='0';
          end if;
        if(oVar1S590(0)='1'  )then
          oVar2S192(0) <='1';
          else
          oVar2S192(0) <='0';
          end if;
        if(oVar1S591(0)='1'  OR oVar1S592(0)='1'  OR oVar1S593(0)='1'  OR oVar1S594(0)='1'  )then
          oVar2S193(0) <='1';
          else
          oVar2S193(0) <='0';
          end if;
        if(oVar1S595(0)='1'  OR oVar1S596(0)='1'  OR oVar1S597(0)='1'  OR oVar1S598(0)='1'  )then
          oVar2S194(0) <='1';
          else
          oVar2S194(0) <='0';
          end if;
        if(oVar1S600(0)='1'  OR oVar1S601(0)='1'  OR oVar1S602(0)='1'  OR oVar1S603(0)='1'  )then
          oVar2S196(0) <='1';
          else
          oVar2S196(0) <='0';
          end if;
        if(oVar1S604(0)='1'  OR oVar1S605(0)='1'  OR oVar1S606(0)='1'  OR oVar1S607(0)='1'  )then
          oVar2S197(0) <='1';
          else
          oVar2S197(0) <='0';
          end if;
        if(oVar1S608(0)='1'  )then
          oVar2S198(0) <='1';
          else
          oVar2S198(0) <='0';
          end if;
        if(oVar1S609(0)='1'  OR oVar1S610(0)='1'  OR oVar1S611(0)='1'  OR oVar1S612(0)='1'  )then
          oVar2S199(0) <='1';
          else
          oVar2S199(0) <='0';
          end if;
        if(oVar1S613(0)='1'  OR oVar1S614(0)='1'  OR oVar1S615(0)='1'  OR oVar1S616(0)='1'  )then
          oVar2S200(0) <='1';
          else
          oVar2S200(0) <='0';
          end if;
        if(oVar1S617(0)='1'  OR oVar1S618(0)='1'  OR oVar1S619(0)='1'  )then
          oVar2S201(0) <='1';
          else
          oVar2S201(0) <='0';
          end if;
        if(oVar1S621(0)='1'  OR oVar1S622(0)='1'  OR oVar1S623(0)='1'  OR oVar1S624(0)='1'  )then
          oVar2S203(0) <='1';
          else
          oVar2S203(0) <='0';
          end if;
        if(oVar1S625(0)='1'  OR oVar1S626(0)='1'  OR oVar1S627(0)='1'  )then
          oVar2S204(0) <='1';
          else
          oVar2S204(0) <='0';
          end if;
        if(oVar1S629(0)='1'  OR oVar1S630(0)='1'  OR oVar1S631(0)='1'  OR oVar1S632(0)='1'  )then
          oVar2S206(0) <='1';
          else
          oVar2S206(0) <='0';
          end if;
        if(oVar1S633(0)='1'  OR oVar1S634(0)='1'  OR oVar1S635(0)='1'  OR oVar1S636(0)='1'  )then
          oVar2S207(0) <='1';
          else
          oVar2S207(0) <='0';
          end if;
        if(oVar1S637(0)='1'  )then
          oVar2S208(0) <='1';
          else
          oVar2S208(0) <='0';
          end if;
        if(oVar1S638(0)='1'  OR oVar1S639(0)='1'  OR oVar1S640(0)='1'  OR oVar1S641(0)='1'  )then
          oVar2S209(0) <='1';
          else
          oVar2S209(0) <='0';
          end if;
        if(oVar1S642(0)='1'  OR oVar1S643(0)='1'  OR oVar1S644(0)='1'  )then
          oVar2S210(0) <='1';
          else
          oVar2S210(0) <='0';
          end if;
        if(oVar1S646(0)='1'  OR oVar1S647(0)='1'  OR oVar1S648(0)='1'  OR oVar1S649(0)='1'  )then
          oVar2S212(0) <='1';
          else
          oVar2S212(0) <='0';
          end if;
        if(oVar1S650(0)='1'  OR oVar1S651(0)='1'  OR oVar1S652(0)='1'  OR oVar1S653(0)='1'  )then
          oVar2S213(0) <='1';
          else
          oVar2S213(0) <='0';
          end if;
        if(oVar1S654(0)='1'  OR oVar1S655(0)='1'  OR oVar1S656(0)='1'  OR oVar1S657(0)='1'  )then
          oVar2S215(0) <='1';
          else
          oVar2S215(0) <='0';
          end if;
        if(oVar1S658(0)='1'  OR oVar1S659(0)='1'  OR oVar1S660(0)='1'  )then
          oVar2S216(0) <='1';
          else
          oVar2S216(0) <='0';
          end if;
        if(oVar1S662(0)='1'  OR oVar1S663(0)='1'  OR oVar1S664(0)='1'  OR oVar1S665(0)='1'  )then
          oVar2S218(0) <='1';
          else
          oVar2S218(0) <='0';
          end if;
        if(oVar1S666(0)='1'  OR oVar1S667(0)='1'  OR oVar1S668(0)='1'  OR oVar1S669(0)='1'  )then
          oVar2S219(0) <='1';
          else
          oVar2S219(0) <='0';
          end if;
        if(oVar1S670(0)='1'  )then
          oVar2S220(0) <='1';
          else
          oVar2S220(0) <='0';
          end if;
        if(oVar1S671(0)='1'  OR oVar1S672(0)='1'  OR oVar1S673(0)='1'  OR oVar1S674(0)='1'  )then
          oVar2S221(0) <='1';
          else
          oVar2S221(0) <='0';
          end if;
        if(oVar1S675(0)='1'  OR oVar1S676(0)='1'  OR oVar1S677(0)='1'  OR oVar1S678(0)='1'  )then
          oVar2S222(0) <='1';
          else
          oVar2S222(0) <='0';
          end if;
        if(oVar1S679(0)='1'  )then
          oVar2S223(0) <='1';
          else
          oVar2S223(0) <='0';
          end if;
        if(oVar1S680(0)='1'  OR oVar1S681(0)='1'  OR oVar1S682(0)='1'  OR oVar1S683(0)='1'  )then
          oVar2S224(0) <='1';
          else
          oVar2S224(0) <='0';
          end if;
        if(oVar1S684(0)='1'  OR oVar1S685(0)='1'  OR oVar1S686(0)='1'  OR oVar1S687(0)='1'  )then
          oVar2S225(0) <='1';
          else
          oVar2S225(0) <='0';
          end if;
        if(oVar1S688(0)='1'  OR oVar1S689(0)='1'  OR oVar1S690(0)='1'  OR oVar1S691(0)='1'  )then
          oVar2S227(0) <='1';
          else
          oVar2S227(0) <='0';
          end if;
        if(oVar1S692(0)='1'  OR oVar1S693(0)='1'  OR oVar1S694(0)='1'  OR oVar1S695(0)='1'  )then
          oVar2S228(0) <='1';
          else
          oVar2S228(0) <='0';
          end if;
        if(oVar1S696(0)='1'  )then
          oVar2S229(0) <='1';
          else
          oVar2S229(0) <='0';
          end if;
        if(oVar1S697(0)='1'  OR oVar1S698(0)='1'  OR oVar1S699(0)='1'  OR oVar1S700(0)='1'  )then
          oVar2S230(0) <='1';
          else
          oVar2S230(0) <='0';
          end if;
        if(oVar1S701(0)='1'  OR oVar1S702(0)='1'  OR oVar1S703(0)='1'  OR oVar1S704(0)='1'  )then
          oVar2S231(0) <='1';
          else
          oVar2S231(0) <='0';
          end if;
        if(oVar1S705(0)='1'  OR oVar1S706(0)='1'  OR oVar1S707(0)='1'  OR oVar1S708(0)='1'  )then
          oVar2S233(0) <='1';
          else
          oVar2S233(0) <='0';
          end if;
        if(oVar1S709(0)='1'  OR oVar1S710(0)='1'  OR oVar1S711(0)='1'  OR oVar1S712(0)='1'  )then
          oVar2S234(0) <='1';
          else
          oVar2S234(0) <='0';
          end if;
        if(oVar1S713(0)='1'  OR oVar1S714(0)='1'  )then
          oVar2S235(0) <='1';
          else
          oVar2S235(0) <='0';
          end if;
        if(oVar1S715(0)='1'  OR oVar1S716(0)='1'  OR oVar1S717(0)='1'  OR oVar1S718(0)='1'  )then
          oVar2S236(0) <='1';
          else
          oVar2S236(0) <='0';
          end if;
        if(oVar1S719(0)='1'  OR oVar1S720(0)='1'  OR oVar1S721(0)='1'  OR oVar1S722(0)='1'  )then
          oVar2S237(0) <='1';
          else
          oVar2S237(0) <='0';
          end if;
        if(oVar1S723(0)='1'  OR oVar1S724(0)='1'  )then
          oVar2S238(0) <='1';
          else
          oVar2S238(0) <='0';
          end if;
        if(oVar1S725(0)='1'  OR oVar1S726(0)='1'  OR oVar1S727(0)='1'  OR oVar1S728(0)='1'  )then
          oVar2S239(0) <='1';
          else
          oVar2S239(0) <='0';
          end if;
        if(oVar1S729(0)='1'  OR oVar1S730(0)='1'  OR oVar1S731(0)='1'  )then
          oVar2S240(0) <='1';
          else
          oVar2S240(0) <='0';
          end if;
        if(oVar1S732(0)='1'  OR oVar1S733(0)='1'  OR oVar1S734(0)='1'  OR oVar1S735(0)='1'  )then
          oVar2S241(0) <='1';
          else
          oVar2S241(0) <='0';
          end if;
        if(oVar1S736(0)='1'  OR oVar1S737(0)='1'  )then
          oVar2S242(0) <='1';
          else
          oVar2S242(0) <='0';
          end if;
        if(oVar1S739(0)='1'  OR oVar1S740(0)='1'  OR oVar1S741(0)='1'  OR oVar1S742(0)='1'  )then
          oVar2S243(0) <='1';
          else
          oVar2S243(0) <='0';
          end if;
        if(oVar1S743(0)='1'  OR oVar1S744(0)='1'  OR oVar1S745(0)='1'  OR oVar1S746(0)='1'  )then
          oVar2S244(0) <='1';
          else
          oVar2S244(0) <='0';
          end if;
        if(oVar1S747(0)='1'  OR oVar1S748(0)='1'  )then
          oVar2S245(0) <='1';
          else
          oVar2S245(0) <='0';
          end if;
        if(oVar1S749(0)='1'  OR oVar1S750(0)='1'  OR oVar1S751(0)='1'  OR oVar1S752(0)='1'  )then
          oVar2S246(0) <='1';
          else
          oVar2S246(0) <='0';
          end if;
        if(oVar1S753(0)='1'  OR oVar1S754(0)='1'  OR oVar1S755(0)='1'  OR oVar1S756(0)='1'  )then
          oVar2S247(0) <='1';
          else
          oVar2S247(0) <='0';
          end if;
        if(oVar1S757(0)='1'  OR oVar1S758(0)='1'  OR oVar1S759(0)='1'  )then
          oVar2S248(0) <='1';
          else
          oVar2S248(0) <='0';
          end if;
        if(oVar1S760(0)='1'  OR oVar1S761(0)='1'  OR oVar1S762(0)='1'  OR oVar1S763(0)='1'  )then
          oVar2S249(0) <='1';
          else
          oVar2S249(0) <='0';
          end if;
        if(oVar1S764(0)='1'  OR oVar1S765(0)='1'  OR oVar1S766(0)='1'  OR oVar1S767(0)='1'  )then
          oVar2S250(0) <='1';
          else
          oVar2S250(0) <='0';
          end if;
        if(oVar1S768(0)='1'  OR oVar1S769(0)='1'  OR oVar1S770(0)='1'  )then
          oVar2S251(0) <='1';
          else
          oVar2S251(0) <='0';
          end if;
        if(oVar1S771(0)='1'  OR oVar1S772(0)='1'  OR oVar1S773(0)='1'  OR oVar1S774(0)='1'  )then
          oVar2S252(0) <='1';
          else
          oVar2S252(0) <='0';
          end if;
        if(oVar1S775(0)='1'  OR oVar1S776(0)='1'  OR oVar1S777(0)='1'  OR oVar1S778(0)='1'  )then
          oVar2S253(0) <='1';
          else
          oVar2S253(0) <='0';
          end if;
        if(oVar1S779(0)='1'  OR oVar1S780(0)='1'  )then
          oVar2S254(0) <='1';
          else
          oVar2S254(0) <='0';
          end if;
        if(oVar1S782(0)='1'  OR oVar1S783(0)='1'  OR oVar1S784(0)='1'  OR oVar1S785(0)='1'  )then
          oVar2S255(0) <='1';
          else
          oVar2S255(0) <='0';
          end if;
        if(oVar1S786(0)='1'  OR oVar1S787(0)='1'  OR oVar1S788(0)='1'  OR oVar1S789(0)='1'  )then
          oVar2S256(0) <='1';
          else
          oVar2S256(0) <='0';
          end if;
        if(oVar1S790(0)='1'  )then
          oVar2S257(0) <='1';
          else
          oVar2S257(0) <='0';
          end if;
        if(oVar1S791(0)='1'  OR oVar1S792(0)='1'  OR oVar1S793(0)='1'  OR oVar1S794(0)='1'  )then
          oVar2S258(0) <='1';
          else
          oVar2S258(0) <='0';
          end if;
        if(oVar1S795(0)='1'  OR oVar1S796(0)='1'  OR oVar1S797(0)='1'  OR oVar1S798(0)='1'  )then
          oVar2S259(0) <='1';
          else
          oVar2S259(0) <='0';
          end if;
        if(oVar1S799(0)='1'  )then
          oVar2S260(0) <='1';
          else
          oVar2S260(0) <='0';
          end if;
        if(oVar1S800(0)='1'  OR oVar1S801(0)='1'  OR oVar1S802(0)='1'  OR oVar1S803(0)='1'  )then
          oVar2S261(0) <='1';
          else
          oVar2S261(0) <='0';
          end if;
        if(oVar1S804(0)='1'  OR oVar1S805(0)='1'  OR oVar1S806(0)='1'  OR oVar1S807(0)='1'  )then
          oVar2S262(0) <='1';
          else
          oVar2S262(0) <='0';
          end if;
        if(oVar1S808(0)='1'  OR oVar1S809(0)='1'  OR oVar1S810(0)='1'  OR oVar1S811(0)='1'  )then
          oVar2S264(0) <='1';
          else
          oVar2S264(0) <='0';
          end if;
        if(oVar1S812(0)='1'  OR oVar1S813(0)='1'  OR oVar1S814(0)='1'  OR oVar1S815(0)='1'  )then
          oVar2S265(0) <='1';
          else
          oVar2S265(0) <='0';
          end if;
        if(oVar1S816(0)='1'  OR oVar1S817(0)='1'  OR oVar1S818(0)='1'  OR oVar1S819(0)='1'  )then
          oVar2S267(0) <='1';
          else
          oVar2S267(0) <='0';
          end if;
        if(oVar1S820(0)='1'  OR oVar1S821(0)='1'  OR oVar1S822(0)='1'  OR oVar1S823(0)='1'  )then
          oVar2S268(0) <='1';
          else
          oVar2S268(0) <='0';
          end if;
        if(oVar1S824(0)='1'  )then
          oVar2S269(0) <='1';
          else
          oVar2S269(0) <='0';
          end if;
        if(oVar1S826(0)='1'  OR oVar1S827(0)='1'  OR oVar1S828(0)='1'  OR oVar1S829(0)='1'  )then
          oVar2S270(0) <='1';
          else
          oVar2S270(0) <='0';
          end if;
        if(oVar1S830(0)='1'  OR oVar1S831(0)='1'  OR oVar1S832(0)='1'  OR oVar1S833(0)='1'  )then
          oVar2S271(0) <='1';
          else
          oVar2S271(0) <='0';
          end if;
        if(oVar1S834(0)='1'  )then
          oVar2S272(0) <='1';
          else
          oVar2S272(0) <='0';
          end if;
        if(oVar1S836(0)='1'  OR oVar1S837(0)='1'  OR oVar1S838(0)='1'  OR oVar1S839(0)='1'  )then
          oVar2S273(0) <='1';
          else
          oVar2S273(0) <='0';
          end if;
        if(oVar1S840(0)='1'  OR oVar1S841(0)='1'  OR oVar1S842(0)='1'  OR oVar1S843(0)='1'  )then
          oVar2S274(0) <='1';
          else
          oVar2S274(0) <='0';
          end if;
        if(oVar1S844(0)='1'  OR oVar1S845(0)='1'  )then
          oVar2S275(0) <='1';
          else
          oVar2S275(0) <='0';
          end if;
        if(oVar1S846(0)='1'  OR oVar1S847(0)='1'  OR oVar1S848(0)='1'  OR oVar1S849(0)='1'  )then
          oVar2S276(0) <='1';
          else
          oVar2S276(0) <='0';
          end if;
        if(oVar1S850(0)='1'  OR oVar1S851(0)='1'  OR oVar1S852(0)='1'  OR oVar1S853(0)='1'  )then
          oVar2S277(0) <='1';
          else
          oVar2S277(0) <='0';
          end if;
        if(oVar1S854(0)='1'  OR oVar1S855(0)='1'  OR oVar1S856(0)='1'  )then
          oVar2S278(0) <='1';
          else
          oVar2S278(0) <='0';
          end if;
        if(oVar1S857(0)='1'  OR oVar1S858(0)='1'  OR oVar1S859(0)='1'  OR oVar1S860(0)='1'  )then
          oVar2S279(0) <='1';
          else
          oVar2S279(0) <='0';
          end if;
        if(oVar1S861(0)='1'  OR oVar1S862(0)='1'  OR oVar1S863(0)='1'  OR oVar1S864(0)='1'  )then
          oVar2S280(0) <='1';
          else
          oVar2S280(0) <='0';
          end if;
        if(oVar1S865(0)='1'  OR oVar1S866(0)='1'  )then
          oVar2S281(0) <='1';
          else
          oVar2S281(0) <='0';
          end if;
        if(oVar1S867(0)='1'  OR oVar1S868(0)='1'  OR oVar1S869(0)='1'  OR oVar1S870(0)='1'  )then
          oVar2S282(0) <='1';
          else
          oVar2S282(0) <='0';
          end if;
        if(oVar1S871(0)='1'  OR oVar1S872(0)='1'  OR oVar1S873(0)='1'  OR oVar1S874(0)='1'  )then
          oVar2S283(0) <='1';
          else
          oVar2S283(0) <='0';
          end if;
        if(oVar1S876(0)='1'  OR oVar1S877(0)='1'  OR oVar1S878(0)='1'  OR oVar1S879(0)='1'  )then
          oVar2S285(0) <='1';
          else
          oVar2S285(0) <='0';
          end if;
        if(oVar1S880(0)='1'  OR oVar1S881(0)='1'  OR oVar1S882(0)='1'  OR oVar1S883(0)='1'  )then
          oVar2S286(0) <='1';
          else
          oVar2S286(0) <='0';
          end if;
        if(oVar1S884(0)='1'  OR oVar1S885(0)='1'  OR oVar1S886(0)='1'  OR oVar1S887(0)='1'  )then
          oVar2S288(0) <='1';
          else
          oVar2S288(0) <='0';
          end if;
        if(oVar1S888(0)='1'  OR oVar1S889(0)='1'  OR oVar1S890(0)='1'  OR oVar1S891(0)='1'  )then
          oVar2S289(0) <='1';
          else
          oVar2S289(0) <='0';
          end if;
        if(oVar1S892(0)='1'  OR oVar1S893(0)='1'  )then
          oVar2S290(0) <='1';
          else
          oVar2S290(0) <='0';
          end if;
        if(oVar1S894(0)='1'  OR oVar1S895(0)='1'  OR oVar1S896(0)='1'  OR oVar1S897(0)='1'  )then
          oVar2S291(0) <='1';
          else
          oVar2S291(0) <='0';
          end if;
        if(oVar1S898(0)='1'  OR oVar1S899(0)='1'  OR oVar1S900(0)='1'  OR oVar1S901(0)='1'  )then
          oVar2S292(0) <='1';
          else
          oVar2S292(0) <='0';
          end if;
        if(oVar1S902(0)='1'  OR oVar1S903(0)='1'  )then
          oVar2S293(0) <='1';
          else
          oVar2S293(0) <='0';
          end if;
        if(oVar1S904(0)='1'  OR oVar1S905(0)='1'  OR oVar1S906(0)='1'  OR oVar1S907(0)='1'  )then
          oVar2S294(0) <='1';
          else
          oVar2S294(0) <='0';
          end if;
        if(oVar1S908(0)='1'  OR oVar1S909(0)='1'  OR oVar1S910(0)='1'  OR oVar1S911(0)='1'  )then
          oVar2S295(0) <='1';
          else
          oVar2S295(0) <='0';
          end if;
        if(oVar1S913(0)='1'  OR oVar1S914(0)='1'  OR oVar1S915(0)='1'  OR oVar1S916(0)='1'  )then
          oVar2S297(0) <='1';
          else
          oVar2S297(0) <='0';
          end if;
        if(oVar1S917(0)='1'  OR oVar1S918(0)='1'  OR oVar1S919(0)='1'  OR oVar1S920(0)='1'  )then
          oVar2S298(0) <='1';
          else
          oVar2S298(0) <='0';
          end if;
        if(oVar1S922(0)='1'  OR oVar1S923(0)='1'  OR oVar1S924(0)='1'  OR oVar1S925(0)='1'  )then
          oVar2S300(0) <='1';
          else
          oVar2S300(0) <='0';
          end if;
        if(oVar1S926(0)='1'  OR oVar1S927(0)='1'  OR oVar1S928(0)='1'  OR oVar1S929(0)='1'  )then
          oVar2S301(0) <='1';
          else
          oVar2S301(0) <='0';
          end if;
        if(oVar1S930(0)='1'  OR oVar1S931(0)='1'  OR oVar1S932(0)='1'  OR oVar1S933(0)='1'  )then
          oVar2S303(0) <='1';
          else
          oVar2S303(0) <='0';
          end if;
        if(oVar1S934(0)='1'  OR oVar1S935(0)='1'  )then
          oVar2S304(0) <='1';
          else
          oVar2S304(0) <='0';
          end if;
        if(oVar1S937(0)='1'  OR oVar1S938(0)='1'  OR oVar1S939(0)='1'  OR oVar1S940(0)='1'  )then
          oVar2S305(0) <='1';
          else
          oVar2S305(0) <='0';
          end if;
        if(oVar1S941(0)='1'  OR oVar1S942(0)='1'  OR oVar1S943(0)='1'  OR oVar1S944(0)='1'  )then
          oVar2S306(0) <='1';
          else
          oVar2S306(0) <='0';
          end if;
        if(oVar1S945(0)='1'  OR oVar1S946(0)='1'  OR oVar1S947(0)='1'  OR oVar1S948(0)='1'  )then
          oVar2S308(0) <='1';
          else
          oVar2S308(0) <='0';
          end if;
        if(oVar1S949(0)='1'  OR oVar1S950(0)='1'  OR oVar1S951(0)='1'  OR oVar1S952(0)='1'  )then
          oVar2S309(0) <='1';
          else
          oVar2S309(0) <='0';
          end if;
        if(oVar1S954(0)='1'  OR oVar1S955(0)='1'  OR oVar1S956(0)='1'  OR oVar1S957(0)='1'  )then
          oVar2S311(0) <='1';
          else
          oVar2S311(0) <='0';
          end if;
        if(oVar1S958(0)='1'  OR oVar1S959(0)='1'  OR oVar1S960(0)='1'  OR oVar1S961(0)='1'  )then
          oVar2S312(0) <='1';
          else
          oVar2S312(0) <='0';
          end if;
        if(oVar1S962(0)='1'  )then
          oVar2S313(0) <='1';
          else
          oVar2S313(0) <='0';
          end if;
        if(oVar1S963(0)='1'  OR oVar1S964(0)='1'  OR oVar1S965(0)='1'  OR oVar1S966(0)='1'  )then
          oVar2S314(0) <='1';
          else
          oVar2S314(0) <='0';
          end if;
        if(oVar1S967(0)='1'  OR oVar1S968(0)='1'  OR oVar1S969(0)='1'  OR oVar1S970(0)='1'  )then
          oVar2S315(0) <='1';
          else
          oVar2S315(0) <='0';
          end if;
        if(oVar1S971(0)='1'  OR oVar1S972(0)='1'  )then
          oVar2S316(0) <='1';
          else
          oVar2S316(0) <='0';
          end if;
        if(oVar1S974(0)='1'  OR oVar1S975(0)='1'  OR oVar1S976(0)='1'  OR oVar1S977(0)='1'  )then
          oVar2S317(0) <='1';
          else
          oVar2S317(0) <='0';
          end if;
        if(oVar1S978(0)='1'  OR oVar1S979(0)='1'  OR oVar1S980(0)='1'  OR oVar1S981(0)='1'  )then
          oVar2S318(0) <='1';
          else
          oVar2S318(0) <='0';
          end if;
        if(oVar1S982(0)='1'  OR oVar1S983(0)='1'  OR oVar1S984(0)='1'  OR oVar1S985(0)='1'  )then
          oVar2S320(0) <='1';
          else
          oVar2S320(0) <='0';
          end if;
        if(oVar1S986(0)='1'  OR oVar1S987(0)='1'  OR oVar1S988(0)='1'  )then
          oVar2S321(0) <='1';
          else
          oVar2S321(0) <='0';
          end if;
        if(oVar1S990(0)='1'  OR oVar1S991(0)='1'  OR oVar1S992(0)='1'  OR oVar1S993(0)='1'  )then
          oVar2S323(0) <='1';
          else
          oVar2S323(0) <='0';
          end if;
        if(oVar1S994(0)='1'  OR oVar1S995(0)='1'  OR oVar1S996(0)='1'  )then
          oVar2S324(0) <='1';
          else
          oVar2S324(0) <='0';
          end if;
        if(oVar1S998(0)='1'  OR oVar1S999(0)='1'  OR oVar1S1000(0)='1'  OR oVar1S1001(0)='1'  )then
          oVar2S326(0) <='1';
          else
          oVar2S326(0) <='0';
          end if;
        if(oVar1S1002(0)='1'  OR oVar1S1003(0)='1'  OR oVar1S1004(0)='1'  OR oVar1S1005(0)='1'  )then
          oVar2S327(0) <='1';
          else
          oVar2S327(0) <='0';
          end if;
        if(oVar1S1006(0)='1'  OR oVar1S1007(0)='1'  )then
          oVar2S328(0) <='1';
          else
          oVar2S328(0) <='0';
          end if;
        if(oVar1S1008(0)='1'  OR oVar1S1009(0)='1'  OR oVar1S1010(0)='1'  OR oVar1S1011(0)='1'  )then
          oVar2S329(0) <='1';
          else
          oVar2S329(0) <='0';
          end if;
        if(oVar1S1012(0)='1'  OR oVar1S1013(0)='1'  OR oVar1S1014(0)='1'  OR oVar1S1015(0)='1'  )then
          oVar2S330(0) <='1';
          else
          oVar2S330(0) <='0';
          end if;
        if(oVar1S1016(0)='1'  OR oVar1S1017(0)='1'  OR oVar1S1018(0)='1'  OR oVar1S1019(0)='1'  )then
          oVar2S331(0) <='1';
          else
          oVar2S331(0) <='0';
          end if;
        if(oVar1S1020(0)='1'  OR oVar1S1021(0)='1'  OR oVar1S1022(0)='1'  OR oVar1S1023(0)='1'  )then
          oVar2S333(0) <='1';
          else
          oVar2S333(0) <='0';
          end if;
        if(oVar1S1024(0)='1'  OR oVar1S1025(0)='1'  OR oVar1S1026(0)='1'  OR oVar1S1027(0)='1'  )then
          oVar2S334(0) <='1';
          else
          oVar2S334(0) <='0';
          end if;
        if(oVar1S1028(0)='1'  OR oVar1S1029(0)='1'  )then
          oVar2S335(0) <='1';
          else
          oVar2S335(0) <='0';
          end if;
        if(oVar1S1030(0)='1'  OR oVar1S1031(0)='1'  OR oVar1S1032(0)='1'  OR oVar1S1033(0)='1'  )then
          oVar2S336(0) <='1';
          else
          oVar2S336(0) <='0';
          end if;
        if(oVar1S1034(0)='1'  OR oVar1S1035(0)='1'  OR oVar1S1036(0)='1'  OR oVar1S1037(0)='1'  )then
          oVar2S337(0) <='1';
          else
          oVar2S337(0) <='0';
          end if;
        if(oVar1S1038(0)='1'  OR oVar1S1039(0)='1'  OR oVar1S1040(0)='1'  )then
          oVar2S338(0) <='1';
          else
          oVar2S338(0) <='0';
          end if;
        if(oVar1S1041(0)='1'  OR oVar1S1042(0)='1'  OR oVar1S1043(0)='1'  OR oVar1S1044(0)='1'  )then
          oVar2S339(0) <='1';
          else
          oVar2S339(0) <='0';
          end if;
        if(oVar1S1045(0)='1'  OR oVar1S1046(0)='1'  OR oVar1S1047(0)='1'  OR oVar1S1048(0)='1'  )then
          oVar2S340(0) <='1';
          else
          oVar2S340(0) <='0';
          end if;
        if(oVar1S1049(0)='1'  OR oVar1S1050(0)='1'  OR oVar1S1051(0)='1'  )then
          oVar2S341(0) <='1';
          else
          oVar2S341(0) <='0';
          end if;
        if(oVar1S1052(0)='1'  OR oVar1S1053(0)='1'  OR oVar1S1054(0)='1'  OR oVar1S1055(0)='1'  )then
          oVar2S342(0) <='1';
          else
          oVar2S342(0) <='0';
          end if;
        if(oVar1S1056(0)='1'  OR oVar1S1057(0)='1'  OR oVar1S1058(0)='1'  OR oVar1S1059(0)='1'  )then
          oVar2S343(0) <='1';
          else
          oVar2S343(0) <='0';
          end if;
        if(oVar1S1060(0)='1'  )then
          oVar2S344(0) <='1';
          else
          oVar2S344(0) <='0';
          end if;
        if(oVar1S1062(0)='1'  OR oVar1S1063(0)='1'  OR oVar1S1064(0)='1'  OR oVar1S1065(0)='1'  )then
          oVar2S345(0) <='1';
          else
          oVar2S345(0) <='0';
          end if;
        if(oVar1S1066(0)='1'  OR oVar1S1067(0)='1'  OR oVar1S1068(0)='1'  OR oVar1S1069(0)='1'  )then
          oVar2S346(0) <='1';
          else
          oVar2S346(0) <='0';
          end if;
        if(oVar1S1071(0)='1'  OR oVar1S1072(0)='1'  OR oVar1S1073(0)='1'  OR oVar1S1074(0)='1'  )then
          oVar2S348(0) <='1';
          else
          oVar2S348(0) <='0';
          end if;
        if(oVar1S1075(0)='1'  OR oVar1S1076(0)='1'  OR oVar1S1077(0)='1'  OR oVar1S1078(0)='1'  )then
          oVar2S349(0) <='1';
          else
          oVar2S349(0) <='0';
          end if;
        if(oVar1S1079(0)='1'  )then
          oVar2S350(0) <='1';
          else
          oVar2S350(0) <='0';
          end if;
        if(oVar1S1081(0)='1'  OR oVar1S1082(0)='1'  OR oVar1S1083(0)='1'  OR oVar1S1084(0)='1'  )then
          oVar2S351(0) <='1';
          else
          oVar2S351(0) <='0';
          end if;
        if(oVar1S1085(0)='1'  OR oVar1S1086(0)='1'  OR oVar1S1087(0)='1'  OR oVar1S1088(0)='1'  )then
          oVar2S352(0) <='1';
          else
          oVar2S352(0) <='0';
          end if;
        if(oVar1S1089(0)='1'  OR oVar1S1090(0)='1'  )then
          oVar2S353(0) <='1';
          else
          oVar2S353(0) <='0';
          end if;
        if(oVar1S1091(0)='1'  OR oVar1S1092(0)='1'  OR oVar1S1093(0)='1'  OR oVar1S1094(0)='1'  )then
          oVar2S354(0) <='1';
          else
          oVar2S354(0) <='0';
          end if;
        if(oVar1S1095(0)='1'  OR oVar1S1096(0)='1'  OR oVar1S1097(0)='1'  OR oVar1S1098(0)='1'  )then
          oVar2S355(0) <='1';
          else
          oVar2S355(0) <='0';
          end if;
        if(oVar1S1099(0)='1'  )then
          oVar2S356(0) <='1';
          else
          oVar2S356(0) <='0';
          end if;
        if(oVar1S1100(0)='1'  OR oVar1S1101(0)='1'  OR oVar1S1102(0)='1'  OR oVar1S1103(0)='1'  )then
          oVar2S357(0) <='1';
          else
          oVar2S357(0) <='0';
          end if;
        if(oVar1S1104(0)='1'  OR oVar1S1105(0)='1'  )then
          oVar2S358(0) <='1';
          else
          oVar2S358(0) <='0';
          end if;
        if(oVar1S1107(0)='1'  OR oVar1S1108(0)='1'  OR oVar1S1109(0)='1'  OR oVar1S1110(0)='1'  )then
          oVar2S359(0) <='1';
          else
          oVar2S359(0) <='0';
          end if;
        if(oVar1S1111(0)='1'  OR oVar1S1112(0)='1'  OR oVar1S1113(0)='1'  OR oVar1S1114(0)='1'  )then
          oVar2S360(0) <='1';
          else
          oVar2S360(0) <='0';
          end if;
        if(oVar1S1115(0)='1'  OR oVar1S1116(0)='1'  OR oVar1S1117(0)='1'  )then
          oVar2S361(0) <='1';
          else
          oVar2S361(0) <='0';
          end if;
        if(oVar1S1119(0)='1'  OR oVar1S1120(0)='1'  OR oVar1S1121(0)='1'  OR oVar1S1122(0)='1'  )then
          oVar2S363(0) <='1';
          else
          oVar2S363(0) <='0';
          end if;
        if(oVar1S1123(0)='1'  OR oVar1S1124(0)='1'  OR oVar1S1125(0)='1'  OR oVar1S1126(0)='1'  )then
          oVar2S364(0) <='1';
          else
          oVar2S364(0) <='0';
          end if;
        if(oVar1S1128(0)='1'  OR oVar1S1129(0)='1'  OR oVar1S1130(0)='1'  OR oVar1S1131(0)='1'  )then
          oVar2S366(0) <='1';
          else
          oVar2S366(0) <='0';
          end if;
        if(oVar1S1132(0)='1'  OR oVar1S1133(0)='1'  OR oVar1S1134(0)='1'  OR oVar1S1135(0)='1'  )then
          oVar2S367(0) <='1';
          else
          oVar2S367(0) <='0';
          end if;
        if(oVar1S1136(0)='1'  OR oVar1S1137(0)='1'  )then
          oVar2S368(0) <='1';
          else
          oVar2S368(0) <='0';
          end if;
        if(oVar1S1138(0)='1'  OR oVar1S1139(0)='1'  OR oVar1S1140(0)='1'  OR oVar1S1141(0)='1'  )then
          oVar2S369(0) <='1';
          else
          oVar2S369(0) <='0';
          end if;
        if(oVar1S1142(0)='1'  OR oVar1S1143(0)='1'  OR oVar1S1144(0)='1'  OR oVar1S1145(0)='1'  )then
          oVar2S370(0) <='1';
          else
          oVar2S370(0) <='0';
          end if;
        if(oVar1S1146(0)='1'  OR oVar1S1147(0)='1'  )then
          oVar2S371(0) <='1';
          else
          oVar2S371(0) <='0';
          end if;
        if(oVar1S1148(0)='1'  OR oVar1S1149(0)='1'  OR oVar1S1150(0)='1'  OR oVar1S1151(0)='1'  )then
          oVar2S372(0) <='1';
          else
          oVar2S372(0) <='0';
          end if;
        if(oVar1S1152(0)='1'  OR oVar1S1153(0)='1'  OR oVar1S1154(0)='1'  OR oVar1S1155(0)='1'  )then
          oVar2S373(0) <='1';
          else
          oVar2S373(0) <='0';
          end if;
        if(oVar1S1156(0)='1'  OR oVar1S1157(0)='1'  )then
          oVar2S374(0) <='1';
          else
          oVar2S374(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV5 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar2S199(0)='1' OR oVar2S200(0)='1' OR oVar2S201(0)='1' )then
          ADDM4K3S8(7)<='1';
          else
          ADDM4K3S8(7)<='0';
          end if;
        if(oVar2S329(0)='1' OR oVar2S330(0)='1' OR oVar2S331(0)='1' )then
          ADDM4K3S8(6)<='1';
          else
          ADDM4K3S8(6)<='0';
          end if;
        if(oVar2S196(0)='1' OR oVar2S197(0)='1' OR oVar2S198(0)='1' )then
          ADDM4K3S8(5)<='1';
          else
          ADDM4K3S8(5)<='0';
          end if;
        if(oVar2S173(0)='1' OR oVar2S174(0)='1' OR oVar2S175(0)='1' )then
          ADDM4K3S8(4)<='1';
          else
          ADDM4K3S8(4)<='0';
          end if;
        if(oVar2S127(0)='1' OR oVar2S128(0)='1' )then
          ADDM4K3S8(3)<='1';
          else
          ADDM4K3S8(3)<='0';
          end if;
        if(oVar2S150(0)='1' OR oVar2S151(0)='1' )then
          ADDM4K3S8(2)<='1';
          else
          ADDM4K3S8(2)<='0';
          end if;
        if(oVar2S141(0)='1' OR oVar2S142(0)='1' )then
          ADDM4K3S8(1)<='1';
          else
          ADDM4K3S8(1)<='0';
          end if;
        if(oVar2S81(0)='1' OR oVar2S82(0)='1' )then
          ADDM4K3S8(0)<='1';
          else
          ADDM4K3S8(0)<='0';
          end if;
        if(oVar2S147(0)='1' OR oVar2S148(0)='1' )then
          ADDM4K3S9(7)<='1';
          else
          ADDM4K3S9(7)<='0';
          end if;
        if(oVar2S68(0)='1' OR oVar2S69(0)='1' )then
          ADDM4K3S9(6)<='1';
          else
          ADDM4K3S9(6)<='0';
          end if;
        if(oVar2S159(0)='1' OR oVar2S160(0)='1' )then
          ADDM4K3S9(5)<='1';
          else
          ADDM4K3S9(5)<='0';
          end if;
        if(oVar2S135(0)='1' OR oVar2S136(0)='1' OR oVar2S137(0)='1' )then
          ADDM4K3S9(4)<='1';
          else
          ADDM4K3S9(4)<='0';
          end if;
        if(oVar2S79(0)='1' OR oVar2S80(0)='1' )then
          ADDM4K3S9(3)<='1';
          else
          ADDM4K3S9(3)<='0';
          end if;
        if(oVar2S156(0)='1' OR oVar2S157(0)='1' OR oVar2S158(0)='1' )then
          ADDM4K3S9(2)<='1';
          else
          ADDM4K3S9(2)<='0';
          end if;
        if(oVar2S71(0)='1' OR oVar2S72(0)='1' )then
          ADDM4K3S9(1)<='1';
          else
          ADDM4K3S9(1)<='0';
          end if;
        if(oVar2S168(0)='1' OR oVar2S169(0)='1' OR oVar2S170(0)='1' )then
          ADDM4K3S9(0)<='1';
          else
          ADDM4K3S9(0)<='0';
          end if;
        if(oVar2S112(0)='1' OR oVar2S113(0)='1' OR oVar2S114(0)='1' )then
          ADDM4K3S12(7)<='1';
          else
          ADDM4K3S12(7)<='0';
          end if;
        if(oVar2S60(0)='1' OR oVar2S61(0)='1' OR oVar2S62(0)='1' )then
          ADDM4K3S12(6)<='1';
          else
          ADDM4K3S12(6)<='0';
          end if;
        if(oVar2S109(0)='1' OR oVar2S110(0)='1' OR oVar2S111(0)='1' )then
          ADDM4K3S12(5)<='1';
          else
          ADDM4K3S12(5)<='0';
          end if;
        if(oVar2S100(0)='1' OR oVar2S101(0)='1' )then
          ADDM4K3S12(4)<='1';
          else
          ADDM4K3S12(4)<='0';
          end if;
        if(oVar2S106(0)='1' OR oVar2S107(0)='1' OR oVar2S108(0)='1' )then
          ADDM4K3S12(3)<='1';
          else
          ADDM4K3S12(3)<='0';
          end if;
        if(oVar2S83(0)='1' OR oVar2S84(0)='1' OR oVar2S85(0)='1' )then
          ADDM4K3S12(2)<='1';
          else
          ADDM4K3S12(2)<='0';
          end if;
        if(oVar2S90(0)='1' OR oVar2S91(0)='1' OR oVar2S92(0)='1' )then
          ADDM4K3S12(1)<='1';
          else
          ADDM4K3S12(1)<='0';
          end if;
        if(oVar2S63(0)='1' OR oVar2S64(0)='1' )then
          ADDM4K3S12(0)<='1';
          else
          ADDM4K3S12(0)<='0';
          end if;
        if(oVar2S23(0)='1' OR oVar2S24(0)='1' )then
          ADDM4K3S13(7)<='1';
          else
          ADDM4K3S13(7)<='0';
          end if;
        if(oVar2S103(0)='1' OR oVar2S104(0)='1' OR oVar2S105(0)='1' )then
          ADDM4K3S13(6)<='1';
          else
          ADDM4K3S13(6)<='0';
          end if;
        if(oVar2S74(0)='1' OR oVar2S75(0)='1' OR oVar2S76(0)='1' )then
          ADDM4K3S13(5)<='1';
          else
          ADDM4K3S13(5)<='0';
          end if;
        if(oVar2S57(0)='1' OR oVar2S58(0)='1' OR oVar2S59(0)='1' )then
          ADDM4K3S13(4)<='1';
          else
          ADDM4K3S13(4)<='0';
          end if;
        if(oVar2S42(0)='1' OR oVar2S43(0)='1' )then
          ADDM4K3S13(3)<='1';
          else
          ADDM4K3S13(3)<='0';
          end if;
        if(oVar2S54(0)='1' OR oVar2S55(0)='1' OR oVar2S56(0)='1' )then
          ADDM4K3S13(2)<='1';
          else
          ADDM4K3S13(2)<='0';
          end if;
        if(oVar2S96(0)='1' OR oVar2S97(0)='1' OR oVar2S98(0)='1' )then
          ADDM4K3S13(1)<='1';
          else
          ADDM4K3S13(1)<='0';
          end if;
        if(oVar2S25(0)='1' OR oVar2S26(0)='1' OR oVar2S27(0)='1' )then
          ADDM4K3S13(0)<='1';
          else
          ADDM4K3S13(0)<='0';
          end if;
        if(oVar2S118(0)='1' OR oVar2S119(0)='1' )then
          ADDM4K3S10(7)<='1';
          else
          ADDM4K3S10(7)<='0';
          end if;
        if(oVar2S153(0)='1' OR oVar2S154(0)='1' OR oVar2S155(0)='1' )then
          ADDM4K3S10(6)<='1';
          else
          ADDM4K3S10(6)<='0';
          end if;
        if(oVar2S144(0)='1' OR oVar2S145(0)='1' OR oVar2S146(0)='1' )then
          ADDM4K3S10(5)<='1';
          else
          ADDM4K3S10(5)<='0';
          end if;
        if(oVar2S176(0)='1' OR oVar2S177(0)='1' OR oVar2S178(0)='1' )then
          ADDM4K3S10(4)<='1';
          else
          ADDM4K3S10(4)<='0';
          end if;
        if(oVar2S171(0)='1' OR oVar2S172(0)='1' )then
          ADDM4K3S10(3)<='1';
          else
          ADDM4K3S10(3)<='0';
          end if;
        if(oVar2S182(0)='1' OR oVar2S183(0)='1' )then
          ADDM4K3S10(2)<='1';
          else
          ADDM4K3S10(2)<='0';
          end if;
        if(oVar2S66(0)='1' OR oVar2S67(0)='1' )then
          ADDM4K3S10(1)<='1';
          else
          ADDM4K3S10(1)<='0';
          end if;
        if(oVar2S45(0)='1' OR oVar2S46(0)='1' )then
          ADDM4K3S10(0)<='1';
          else
          ADDM4K3S10(0)<='0';
          end if;
        if(oVar2S179(0)='1' OR oVar2S180(0)='1' OR oVar2S181(0)='1' )then
          ADDM4K3S11(7)<='1';
          else
          ADDM4K3S11(7)<='0';
          end if;
        if(oVar2S124(0)='1' OR oVar2S125(0)='1' OR oVar2S126(0)='1' )then
          ADDM4K3S11(6)<='1';
          else
          ADDM4K3S11(6)<='0';
          end if;
        if(oVar2S129(0)='1' OR oVar2S130(0)='1' )then
          ADDM4K3S11(5)<='1';
          else
          ADDM4K3S11(5)<='0';
          end if;
        if(oVar2S121(0)='1' OR oVar2S122(0)='1' OR oVar2S123(0)='1' )then
          ADDM4K3S11(4)<='1';
          else
          ADDM4K3S11(4)<='0';
          end if;
        if(oVar2S77(0)='1' OR oVar2S78(0)='1' )then
          ADDM4K3S11(3)<='1';
          else
          ADDM4K3S11(3)<='0';
          end if;
        if(oVar2S93(0)='1' OR oVar2S94(0)='1' )then
          ADDM4K3S11(2)<='1';
          else
          ADDM4K3S11(2)<='0';
          end if;
        if(oVar2S115(0)='1' OR oVar2S116(0)='1' OR oVar2S117(0)='1' )then
          ADDM4K3S11(1)<='1';
          else
          ADDM4K3S11(1)<='0';
          end if;
        if(oVar2S132(0)='1' OR oVar2S133(0)='1' OR oVar2S134(0)='1' )then
          ADDM4K3S11(0)<='1';
          else
          ADDM4K3S11(0)<='0';
          end if;
        if(oVar2S86(0)='1' OR oVar2S87(0)='1' OR oVar2S88(0)='1' )then
          ADDM4K3S14(7)<='1';
          else
          ADDM4K3S14(7)<='0';
          end if;
        if(oVar2S31(0)='1' OR oVar2S32(0)='1' )then
          ADDM4K3S14(6)<='1';
          else
          ADDM4K3S14(6)<='0';
          end if;
        if(oVar2S48(0)='1' OR oVar2S49(0)='1' OR oVar2S50(0)='1' )then
          ADDM4K3S14(5)<='1';
          else
          ADDM4K3S14(5)<='0';
          end if;
        if(oVar2S51(0)='1' OR oVar2S52(0)='1' OR oVar2S53(0)='1' )then
          ADDM4K3S14(4)<='1';
          else
          ADDM4K3S14(4)<='0';
          end if;
        if(oVar2S36(0)='1' OR oVar2S37(0)='1' OR oVar2S38(0)='1' )then
          ADDM4K3S14(3)<='1';
          else
          ADDM4K3S14(3)<='0';
          end if;
        if(oVar2S39(0)='1' OR oVar2S40(0)='1' OR oVar2S41(0)='1' )then
          ADDM4K3S14(2)<='1';
          else
          ADDM4K3S14(2)<='0';
          end if;
        if(oVar2S20(0)='1' OR oVar2S21(0)='1' )then
          ADDM4K3S14(1)<='1';
          else
          ADDM4K3S14(1)<='0';
          end if;
        if(oVar2S28(0)='1' OR oVar2S29(0)='1' OR oVar2S30(0)='1' )then
          ADDM4K3S14(0)<='1';
          else
          ADDM4K3S14(0)<='0';
          end if;
        if(oVar2S18(0)='1' OR oVar2S19(0)='1' )then
          ADDM4K3S15(7)<='1';
          else
          ADDM4K3S15(7)<='0';
          end if;
        if(oVar2S33(0)='1' OR oVar2S34(0)='1' OR oVar2S35(0)='1' )then
          ADDM4K3S15(6)<='1';
          else
          ADDM4K3S15(6)<='0';
          end if;
        if(oVar2S15(0)='1' OR oVar2S16(0)='1' OR oVar2S17(0)='1' )then
          ADDM4K3S15(5)<='1';
          else
          ADDM4K3S15(5)<='0';
          end if;
        if(oVar2S12(0)='1' OR oVar2S13(0)='1' )then
          ADDM4K3S15(4)<='1';
          else
          ADDM4K3S15(4)<='0';
          end if;
        if(oVar2S9(0)='1' OR oVar2S10(0)='1' )then
          ADDM4K3S15(3)<='1';
          else
          ADDM4K3S15(3)<='0';
          end if;
        if(oVar2S6(0)='1' OR oVar2S7(0)='1' OR oVar2S8(0)='1' )then
          ADDM4K3S15(2)<='1';
          else
          ADDM4K3S15(2)<='0';
          end if;
        if(oVar2S3(0)='1' OR oVar2S4(0)='1' )then
          ADDM4K3S15(1)<='1';
          else
          ADDM4K3S15(1)<='0';
          end if;
        if(oVar2S0(0)='1' OR oVar2S1(0)='1' OR oVar2S2(0)='1' )then
          ADDM4K3S15(0)<='1';
          else
          ADDM4K3S15(0)<='0';
          end if;
        if(oVar2S185(0)='1' OR oVar2S186(0)='1' )then
          ADDM4K3S2(7)<='1';
          else
          ADDM4K3S2(7)<='0';
          end if;
        if(oVar2S363(0)='1' OR oVar2S364(0)='1' )then
          ADDM4K3S2(6)<='1';
          else
          ADDM4K3S2(6)<='0';
          end if;
        if(oVar2S209(0)='1' OR oVar2S210(0)='1' )then
          ADDM4K3S2(5)<='1';
          else
          ADDM4K3S2(5)<='0';
          end if;
        if(oVar2S267(0)='1' OR oVar2S268(0)='1' OR oVar2S269(0)='1' )then
          ADDM4K3S2(4)<='1';
          else
          ADDM4K3S2(4)<='0';
          end if;
        if(oVar2S291(0)='1' OR oVar2S292(0)='1' OR oVar2S293(0)='1' )then
          ADDM4K3S2(3)<='1';
          else
          ADDM4K3S2(3)<='0';
          end if;
        if(oVar2S288(0)='1' OR oVar2S289(0)='1' OR oVar2S290(0)='1' )then
          ADDM4K3S2(2)<='1';
          else
          ADDM4K3S2(2)<='0';
          end if;
        if(oVar2S270(0)='1' OR oVar2S271(0)='1' OR oVar2S272(0)='1' )then
          ADDM4K3S2(1)<='1';
          else
          ADDM4K3S2(1)<='0';
          end if;
        if(oVar2S285(0)='1' OR oVar2S286(0)='1' )then
          ADDM4K3S2(0)<='1';
          else
          ADDM4K3S2(0)<='0';
          end if;
        if(oVar2S300(0)='1' OR oVar2S301(0)='1' )then
          ADDM4K3S3(7)<='1';
          else
          ADDM4K3S3(7)<='0';
          end if;
        if(oVar2S372(0)='1' OR oVar2S373(0)='1' OR oVar2S374(0)='1' )then
          ADDM4K3S3(6)<='1';
          else
          ADDM4K3S3(6)<='0';
          end if;
        if(oVar2S294(0)='1' OR oVar2S295(0)='1' )then
          ADDM4K3S3(5)<='1';
          else
          ADDM4K3S3(5)<='0';
          end if;
        if(oVar2S333(0)='1' OR oVar2S334(0)='1' OR oVar2S335(0)='1' )then
          ADDM4K3S3(4)<='1';
          else
          ADDM4K3S3(4)<='0';
          end if;
        if(oVar2S224(0)='1' OR oVar2S225(0)='1' )then
          ADDM4K3S3(3)<='1';
          else
          ADDM4K3S3(3)<='0';
          end if;
        if(oVar2S345(0)='1' OR oVar2S346(0)='1' )then
          ADDM4K3S3(2)<='1';
          else
          ADDM4K3S3(2)<='0';
          end if;
        if(oVar2S351(0)='1' OR oVar2S352(0)='1' OR oVar2S353(0)='1' )then
          ADDM4K3S3(1)<='1';
          else
          ADDM4K3S3(1)<='0';
          end if;
        if(oVar2S348(0)='1' OR oVar2S349(0)='1' OR oVar2S350(0)='1' )then
          ADDM4K3S3(0)<='1';
          else
          ADDM4K3S3(0)<='0';
          end if;
        if(oVar2S297(0)='1' OR oVar2S298(0)='1' )then
          ADDM4K3S4(7)<='1';
          else
          ADDM4K3S4(7)<='0';
          end if;
        if(oVar2S255(0)='1' OR oVar2S256(0)='1' OR oVar2S257(0)='1' )then
          ADDM4K3S4(6)<='1';
          else
          ADDM4K3S4(6)<='0';
          end if;
        if(oVar2S165(0)='1' OR oVar2S166(0)='1' )then
          ADDM4K3S4(5)<='1';
          else
          ADDM4K3S4(5)<='0';
          end if;
        if(oVar2S239(0)='1' OR oVar2S240(0)='1' )then
          ADDM4K3S4(4)<='1';
          else
          ADDM4K3S4(4)<='0';
          end if;
        if(oVar2S276(0)='1' OR oVar2S277(0)='1' OR oVar2S278(0)='1' )then
          ADDM4K3S4(3)<='1';
          else
          ADDM4K3S4(3)<='0';
          end if;
        if(oVar2S317(0)='1' OR oVar2S318(0)='1' )then
          ADDM4K3S4(2)<='1';
          else
          ADDM4K3S4(2)<='0';
          end if;
        if(oVar2S187(0)='1' OR oVar2S188(0)='1' )then
          ADDM4K3S4(1)<='1';
          else
          ADDM4K3S4(1)<='0';
          end if;
        if(oVar2S359(0)='1' OR oVar2S360(0)='1' OR oVar2S361(0)='1' )then
          ADDM4K3S4(0)<='1';
          else
          ADDM4K3S4(0)<='0';
          end if;
        if(oVar2S190(0)='1' OR oVar2S191(0)='1' OR oVar2S192(0)='1' )then
          ADDM4K3S5(7)<='1';
          else
          ADDM4K3S5(7)<='0';
          end if;
        if(oVar2S342(0)='1' OR oVar2S343(0)='1' OR oVar2S344(0)='1' )then
          ADDM4K3S5(6)<='1';
          else
          ADDM4K3S5(6)<='0';
          end if;
        if(oVar2S282(0)='1' OR oVar2S283(0)='1' )then
          ADDM4K3S5(5)<='1';
          else
          ADDM4K3S5(5)<='0';
          end if;
        if(oVar2S314(0)='1' OR oVar2S315(0)='1' OR oVar2S316(0)='1' )then
          ADDM4K3S5(4)<='1';
          else
          ADDM4K3S5(4)<='0';
          end if;
        if(oVar2S326(0)='1' OR oVar2S327(0)='1' OR oVar2S328(0)='1' )then
          ADDM4K3S5(3)<='1';
          else
          ADDM4K3S5(3)<='0';
          end if;
        if(oVar2S230(0)='1' OR oVar2S231(0)='1' )then
          ADDM4K3S5(2)<='1';
          else
          ADDM4K3S5(2)<='0';
          end if;
        if(oVar2S227(0)='1' OR oVar2S228(0)='1' OR oVar2S229(0)='1' )then
          ADDM4K3S5(1)<='1';
          else
          ADDM4K3S5(1)<='0';
          end if;
        if(oVar2S236(0)='1' OR oVar2S237(0)='1' OR oVar2S238(0)='1' )then
          ADDM4K3S5(0)<='1';
          else
          ADDM4K3S5(0)<='0';
          end if;
        if(oVar2S252(0)='1' OR oVar2S253(0)='1' OR oVar2S254(0)='1' )then
          ADDM4K3S6(7)<='1';
          else
          ADDM4K3S6(7)<='0';
          end if;
        if(oVar2S273(0)='1' OR oVar2S274(0)='1' OR oVar2S275(0)='1' )then
          ADDM4K3S6(6)<='1';
          else
          ADDM4K3S6(6)<='0';
          end if;
        if(oVar2S279(0)='1' OR oVar2S280(0)='1' OR oVar2S281(0)='1' )then
          ADDM4K3S6(5)<='1';
          else
          ADDM4K3S6(5)<='0';
          end if;
        if(oVar2S339(0)='1' OR oVar2S340(0)='1' OR oVar2S341(0)='1' )then
          ADDM4K3S6(4)<='1';
          else
          ADDM4K3S6(4)<='0';
          end if;
        if(oVar2S206(0)='1' OR oVar2S207(0)='1' OR oVar2S208(0)='1' )then
          ADDM4K3S6(3)<='1';
          else
          ADDM4K3S6(3)<='0';
          end if;
        if(oVar2S336(0)='1' OR oVar2S337(0)='1' OR oVar2S338(0)='1' )then
          ADDM4K3S6(2)<='1';
          else
          ADDM4K3S6(2)<='0';
          end if;
        if(oVar2S233(0)='1' OR oVar2S234(0)='1' OR oVar2S235(0)='1' )then
          ADDM4K3S6(1)<='1';
          else
          ADDM4K3S6(1)<='0';
          end if;
        if(oVar2S218(0)='1' OR oVar2S219(0)='1' OR oVar2S220(0)='1' )then
          ADDM4K3S6(0)<='1';
          else
          ADDM4K3S6(0)<='0';
          end if;
        if(oVar2S249(0)='1' OR oVar2S250(0)='1' OR oVar2S251(0)='1' )then
          ADDM4K3S7(7)<='1';
          else
          ADDM4K3S7(7)<='0';
          end if;
        if(oVar2S162(0)='1' OR oVar2S163(0)='1' )then
          ADDM4K3S7(6)<='1';
          else
          ADDM4K3S7(6)<='0';
          end if;
        if(oVar2S243(0)='1' OR oVar2S244(0)='1' OR oVar2S245(0)='1' )then
          ADDM4K3S7(5)<='1';
          else
          ADDM4K3S7(5)<='0';
          end if;
        if(oVar2S221(0)='1' OR oVar2S222(0)='1' OR oVar2S223(0)='1' )then
          ADDM4K3S7(4)<='1';
          else
          ADDM4K3S7(4)<='0';
          end if;
        if(oVar2S138(0)='1' OR oVar2S139(0)='1' )then
          ADDM4K3S7(3)<='1';
          else
          ADDM4K3S7(3)<='0';
          end if;
        if(oVar2S203(0)='1' OR oVar2S204(0)='1' )then
          ADDM4K3S7(2)<='1';
          else
          ADDM4K3S7(2)<='0';
          end if;
        if(oVar2S246(0)='1' OR oVar2S247(0)='1' OR oVar2S248(0)='1' )then
          ADDM4K3S7(1)<='1';
          else
          ADDM4K3S7(1)<='0';
          end if;
        if(oVar2S193(0)='1' OR oVar2S194(0)='1' )then
          ADDM4K3S7(0)<='1';
          else
          ADDM4K3S7(0)<='0';
          end if;
        if(oVar2S354(0)='1' OR oVar2S355(0)='1' OR oVar2S356(0)='1' )then
          ADDM4K3S0(7)<='1';
          else
          ADDM4K3S0(7)<='0';
          end if;
        if(oVar2S264(0)='1' OR oVar2S265(0)='1' )then
          ADDM4K3S0(6)<='1';
          else
          ADDM4K3S0(6)<='0';
          end if;
        if(oVar2S215(0)='1' OR oVar2S216(0)='1' )then
          ADDM4K3S0(5)<='1';
          else
          ADDM4K3S0(5)<='0';
          end if;
        if(oVar2S303(0)='1' OR oVar2S304(0)='1' )then
          ADDM4K3S0(4)<='1';
          else
          ADDM4K3S0(4)<='0';
          end if;
        if(oVar2S258(0)='1' OR oVar2S259(0)='1' OR oVar2S260(0)='1' )then
          ADDM4K3S0(3)<='1';
          else
          ADDM4K3S0(3)<='0';
          end if;
        if(oVar2S308(0)='1' OR oVar2S309(0)='1' )then
          ADDM4K3S0(2)<='1';
          else
          ADDM4K3S0(2)<='0';
          end if;
        if(oVar2S357(0)='1' OR oVar2S358(0)='1' )then
          ADDM4K3S0(1)<='1';
          else
          ADDM4K3S0(1)<='0';
          end if;
        if(oVar2S305(0)='1' OR oVar2S306(0)='1' )then
          ADDM4K3S0(0)<='1';
          else
          ADDM4K3S0(0)<='0';
          end if;
        if(oVar2S212(0)='1' OR oVar2S213(0)='1' )then
          ADDM4K3S1(7)<='1';
          else
          ADDM4K3S1(7)<='0';
          end if;
        if(oVar2S320(0)='1' OR oVar2S321(0)='1' )then
          ADDM4K3S1(6)<='1';
          else
          ADDM4K3S1(6)<='0';
          end if;
        if(oVar2S241(0)='1' OR oVar2S242(0)='1' )then
          ADDM4K3S1(5)<='1';
          else
          ADDM4K3S1(5)<='0';
          end if;
        if(oVar2S323(0)='1' OR oVar2S324(0)='1' )then
          ADDM4K3S1(4)<='1';
          else
          ADDM4K3S1(4)<='0';
          end if;
        if(oVar2S369(0)='1' OR oVar2S370(0)='1' OR oVar2S371(0)='1' )then
          ADDM4K3S1(3)<='1';
          else
          ADDM4K3S1(3)<='0';
          end if;
        if(oVar2S261(0)='1' OR oVar2S262(0)='1' )then
          ADDM4K3S1(2)<='1';
          else
          ADDM4K3S1(2)<='0';
          end if;
        if(oVar2S366(0)='1' OR oVar2S367(0)='1' OR oVar2S368(0)='1' )then
          ADDM4K3S1(1)<='1';
          else
          ADDM4K3S1(1)<='0';
          end if;
        if(oVar2S311(0)='1' OR oVar2S312(0)='1' OR oVar2S313(0)='1' )then
          ADDM4K3S1(0)<='1';
          else
          ADDM4K3S1(0)<='0';
          end if;
 end if;
end process;
ADDM4K3S8c : ADDM4K3S8RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S8,
                q    => aVar3S8
    );
ADDM4K3S9c : ADDM4K3S9RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S9,
                q    => aVar3S9
    );
ADDM4K3S12c : ADDM4K3S12RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S12,
                q    => aVar3S12
    );
ADDM4K3S13c : ADDM4K3S13RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S13,
                q    => aVar3S13
    );
ADDM4K3S10c : ADDM4K3S10RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S10,
                q    => aVar3S10
    );
ADDM4K3S11c : ADDM4K3S11RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S11,
                q    => aVar3S11
    );
ADDM4K3S14c : ADDM4K3S14RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S14,
                q    => aVar3S14
    );
ADDM4K3S15c : ADDM4K3S15RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S15,
                q    => aVar3S15
    );
ADDM4K3S2c : ADDM4K3S2RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S2,
                q    => aVar3S2
    );
ADDM4K3S3c : ADDM4K3S3RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S3,
                q    => aVar3S3
    );
ADDM4K3S4c : ADDM4K3S4RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S4,
                q    => aVar3S4
    );
ADDM4K3S5c : ADDM4K3S5RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S5,
                q    => aVar3S5
    );
ADDM4K3S6c : ADDM4K3S6RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S6,
                q    => aVar3S6
    );
ADDM4K3S7c : ADDM4K3S7RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S7,
                q    => aVar3S7
    );
ADDM4K3S0c : ADDM4K3S0RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S0,
                q    => aVar3S0
    );
ADDM4K3S1c : ADDM4K3S1RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S1,
                q    => aVar3S1
    );
Adder_1: Adder_type
port map(
dataa => aVar3S0, 
datab => aVar3S1, 
result => aVar4S0
);

Adder_2: Adder_type
port map(
dataa => aVar3S2, 
datab => aVar3S3, 
result => aVar4S1
);

Adder_3: Adder_type
port map(
dataa => aVar3S4, 
datab => aVar3S5, 
result => aVar4S2
);

Adder_4: Adder_type
port map(
dataa => aVar3S6, 
datab => aVar3S7, 
result => aVar4S3
);

Adder_5: Adder_type
port map(
dataa => aVar3S8, 
datab => aVar3S9, 
result => aVar4S4
);

Adder_6: Adder_type
port map(
dataa => aVar3S10, 
datab => aVar3S11, 
result => aVar4S5
);

Adder_7: Adder_type
port map(
dataa => aVar3S12, 
datab => aVar3S13, 
result => aVar4S6
);

Adder_8: Adder_type
port map(
dataa => aVar3S14, 
datab => aVar3S15, 
result => aVar4S7
);

Adder_9: Adder_type
port map(
dataa => aVar4S0, 
datab => aVar4S1, 
result => aVar5S0
);

Adder_10: Adder_type
port map(
dataa => aVar4S2, 
datab => aVar4S3, 
result => aVar5S1
);

Adder_11: Adder_type
port map(
dataa => aVar4S4, 
datab => aVar4S5, 
result => aVar5S2
);

Adder_12: Adder_type
port map(
dataa => aVar4S6, 
datab => aVar4S7, 
result => aVar5S3
);

Adder_13: Adder_type
port map(
dataa => aVar5S0, 
datab => aVar5S1, 
result => aVar6S0
);

Adder_14: Adder_type
port map(
dataa => aVar5S2, 
datab => aVar5S3, 
result => aVar6S1
);

Adder_15: Adder_type
port map(
dataa => aVar6S0, 
datab => aVar6S1, 
result => aVar7S0
);

	 output (15 downto 0)<= aVar7S0 (15 downto 0) ;
end rtl;
