LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY code_450 IS
   PORT(
      --*************************************************
      -- V1495 Front Panel Ports (PORT A,B,C,G)
      --*************************************************
      A_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In A (32 x LVDS/ECL)
      B_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In B (32 x LVDS/ECL)
      D_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In D (32 x LVDS/ECL)
      E_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In E (32 x LVDS/ECL)
      F_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- OUT F (32 x LVDS/ECL)
      C_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- Out C (32 x LVDS)
      c1            : IN STD_LOGIC                            -- the PLL1 output
   );
END code_450 ;
ARCHITECTURE rtl OF code_450 IS
	signal A     : std_logic_vector(31 downto 0);
	signal B     : std_logic_vector(31 downto 0);
	signal C     : std_logic_vector(31 downto 0);
	signal D     : std_logic_vector(31 downto 0);
	signal E     : std_logic_vector(31 downto 0);
	signal F     : std_logic_vector(31 downto 0);
	signal G     : std_logic_vector(1 downto 0);
	signal output	: std_logic_vector(15 downto 0);
component Adder_type
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		overflow		: OUT STD_LOGIC_VECTOR ;
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
end component;
component  ADDM4K3S8RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S9RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S12RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S13RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S10RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S11RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S14RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S15RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S2RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S3RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S4RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S5RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S6RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S7RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S0RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S1RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

        signal cVar1S0S0P055P030nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S0P055N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S0P055N030N031P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S0P055N030N031N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S0P055N030N031N028: std_logic_vector(   0 downto 0);
        signal cVar1S5S0P055N030N031N028: std_logic_vector(   0 downto 0);
        signal cVar1S6S0N055P059P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S0N055P059P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S8S0N055P059P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S9S0N055P059P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S10S0N055P059N061P058nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S0N055P059N061N058: std_logic_vector(   0 downto 0);
        signal cVar1S12S0N055P059N061N058: std_logic_vector(   0 downto 0);
        signal cVar1S13S0N055P059N061N058: std_logic_vector(   0 downto 0);
        signal cVar1S14S0N055N059P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S0N055N059P052N029: std_logic_vector(   0 downto 0);
        signal cVar1S16S0N055N059P052N029: std_logic_vector(   0 downto 0);
        signal cVar1S17S0N055N059P052N029: std_logic_vector(   0 downto 0);
        signal cVar1S18S0N055N059N052P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S0N055N059N052P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S0N055N059N052P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S0N055N059N052N047: std_logic_vector(   0 downto 0);
        signal cVar1S22S0N055N059N052N047: std_logic_vector(   0 downto 0);
        signal cVar1S23S0N055N059N052N047: std_logic_vector(   0 downto 0);
        signal cVar1S0S1P058P033P060nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S1P058P033N060P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S1P058P033N060P018: std_logic_vector(   0 downto 0);
        signal cVar1S3S1P058N033P031nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S1P058N033N031P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S1P058N033N031N032: std_logic_vector(   0 downto 0);
        signal cVar1S6S1P058N033N031N032: std_logic_vector(   0 downto 0);
        signal cVar1S7S1P058N033N031N032: std_logic_vector(   0 downto 0);
        signal cVar1S8S1N058P051P053P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S1N058P051P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S10S1N058P051P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S1N058P051P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S12S1N058P051N053P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S1N058P051N053N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S1N058P051N053N026: std_logic_vector(   0 downto 0);
        signal cVar1S15S1N058P051N053N026: std_logic_vector(   0 downto 0);
        signal cVar1S16S1N058N051P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S1N058N051P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S18S1N058N051P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S19S1N058N051P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S20S1N058N051N046P064: std_logic_vector(   0 downto 0);
        signal cVar1S21S1N058N051N046P064: std_logic_vector(   0 downto 0);
        signal cVar1S22S1N058N051N046P064: std_logic_vector(   0 downto 0);
        signal cVar1S23S1N058N051N046N064: std_logic_vector(   0 downto 0);
        signal cVar1S24S1N058N051N046N064: std_logic_vector(   0 downto 0);
        signal cVar1S25S1N058N051N046N064: std_logic_vector(   0 downto 0);
        signal cVar1S26S1N058N051N046N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S2P068P019P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S2P068P019P015N066: std_logic_vector(   0 downto 0);
        signal cVar1S2S2P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S3S2P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S4S2P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S5S2P068N019P011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S2P068N019P011N018: std_logic_vector(   0 downto 0);
        signal cVar1S7S2P068N019P011N018: std_logic_vector(   0 downto 0);
        signal cVar1S8S2P068N019P011P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S2P068N019P011P067: std_logic_vector(   0 downto 0);
        signal cVar1S10S2P068N019P011P067: std_logic_vector(   0 downto 0);
        signal cVar1S11S2N068P040P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S2N068P040N038P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S2N068P040N038N023: std_logic_vector(   0 downto 0);
        signal cVar1S14S2N068P040N038N023: std_logic_vector(   0 downto 0);
        signal cVar1S15S2N068P040N038N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S2N068N040P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S2N068N040P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S18S2N068N040P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S19S2N068N040P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S20S2N068N040N050P046: std_logic_vector(   0 downto 0);
        signal cVar1S21S2N068N040N050P046: std_logic_vector(   0 downto 0);
        signal cVar1S22S2N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S23S2N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S24S2N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S0S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S1S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S2S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S3S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S4S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S5S3P068P019P015P017: std_logic_vector(   0 downto 0);
        signal cVar1S6S3P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S7S3P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S8S3P068P019P015P064: std_logic_vector(   0 downto 0);
        signal cVar1S9S3P068N019P018P001: std_logic_vector(   0 downto 0);
        signal cVar1S10S3P068N019P018P001: std_logic_vector(   0 downto 0);
        signal cVar1S11S3P068N019P018P001: std_logic_vector(   0 downto 0);
        signal cVar1S12S3P068N019P018P001: std_logic_vector(   0 downto 0);
        signal cVar1S13S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S14S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S15S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S16S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S17S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S18S3P068N019N018P010: std_logic_vector(   0 downto 0);
        signal cVar1S19S3N068P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S3N068P040N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S3N068P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S22S3N068P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S23S3N068P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S24S3N068N040P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S3N068N040N050P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S3N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S27S3N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S28S3N068N040N050N046: std_logic_vector(   0 downto 0);
        signal cVar1S0S4P040P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S4P040N038P067P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S4P040N038P067N023: std_logic_vector(   0 downto 0);
        signal cVar1S3S4N040P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S4N040P044N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S4N040P044N023N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S4N040P044N023N022: std_logic_vector(   0 downto 0);
        signal cVar1S7S4N040P044N023N022: std_logic_vector(   0 downto 0);
        signal cVar1S8S4N040N044P047P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S4N040N044P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S10S4N040N044P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S11S4N040N044P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S12S4N040N044N047P061: std_logic_vector(   0 downto 0);
        signal cVar1S13S4N040N044N047P061: std_logic_vector(   0 downto 0);
        signal cVar1S14S4N040N044N047P061: std_logic_vector(   0 downto 0);
        signal cVar1S15S4N040N044N047P061: std_logic_vector(   0 downto 0);
        signal cVar1S16S4N040N044N047N061: std_logic_vector(   0 downto 0);
        signal cVar1S17S4N040N044N047N061: std_logic_vector(   0 downto 0);
        signal cVar1S18S4N040N044N047N061: std_logic_vector(   0 downto 0);
        signal cVar1S0S5P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S5P044N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S5P044N023N022P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S5P044N023N022N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S5P044N023N022N025: std_logic_vector(   0 downto 0);
        signal cVar1S5S5N044P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S5N044P040N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S5N044P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S8S5N044P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S9S5N044P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S10S5N044N040P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S5N044N040P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S12S5N044N040P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S13S5N044N040N047P056: std_logic_vector(   0 downto 0);
        signal cVar1S14S5N044N040N047P056: std_logic_vector(   0 downto 0);
        signal cVar1S15S5N044N040N047P056: std_logic_vector(   0 downto 0);
        signal cVar1S16S5N044N040N047P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S5N044N040N047N056: std_logic_vector(   0 downto 0);
        signal cVar1S18S5N044N040N047N056: std_logic_vector(   0 downto 0);
        signal cVar1S19S5N044N040N047N056: std_logic_vector(   0 downto 0);
        signal cVar1S20S5N044N040N047N056: std_logic_vector(   0 downto 0);
        signal cVar1S0S6P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S6P044N023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S6P044N023N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S6P044N023N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S6P044N023N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S6N044P015P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S6N044P015P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S7S6N044P015P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S8S6N044P015P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S6N044P015N050P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S6N044P015N050P056: std_logic_vector(   0 downto 0);
        signal cVar1S11S6N044P015N050P056: std_logic_vector(   0 downto 0);
        signal cVar1S12S6N044P015N050N056: std_logic_vector(   0 downto 0);
        signal cVar1S13S6N044P015N050N056: std_logic_vector(   0 downto 0);
        signal cVar1S14S6N044P015P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S15S6N044P015P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S16S6N044P015P062P035: std_logic_vector(   0 downto 0);
        signal cVar1S17S6N044P015P062N035: std_logic_vector(   0 downto 0);
        signal cVar1S18S6N044P015P062N035: std_logic_vector(   0 downto 0);
        signal cVar1S19S6N044P015N062P058: std_logic_vector(   0 downto 0);
        signal cVar1S20S6N044P015N062P058: std_logic_vector(   0 downto 0);
        signal cVar1S21S6N044P015N062N058: std_logic_vector(   0 downto 0);
        signal cVar1S22S6N044P015N062N058: std_logic_vector(   0 downto 0);
        signal cVar1S23S6N044P015N062N058: std_logic_vector(   0 downto 0);
        signal cVar1S24S6N044P015N062N058: std_logic_vector(   0 downto 0);
        signal cVar1S0S7P050P027P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S7P050P027N048P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S7P050P027N048N009: std_logic_vector(   0 downto 0);
        signal cVar1S3S7P050P027N048N009: std_logic_vector(   0 downto 0);
        signal cVar1S4S7P050N027P052P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S7P050N027P052N008: std_logic_vector(   0 downto 0);
        signal cVar1S6S7P050N027P052N008: std_logic_vector(   0 downto 0);
        signal cVar1S7S7P050N027P052N008: std_logic_vector(   0 downto 0);
        signal cVar1S8S7P050N027N052P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S7P050N027N052P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S7P050N027N052N048: std_logic_vector(   0 downto 0);
        signal cVar1S11S7N050P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S7N050P044N023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S7N050P044N023N004: std_logic_vector(   0 downto 0);
        signal cVar1S14S7N050P044N023N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S7N050P044N023N004: std_logic_vector(   0 downto 0);
        signal cVar1S16S7N050N044P056P031: std_logic_vector(   0 downto 0);
        signal cVar1S17S7N050N044P056P031: std_logic_vector(   0 downto 0);
        signal cVar1S18S7N050N044P056N031: std_logic_vector(   0 downto 0);
        signal cVar1S19S7N050N044P056N031: std_logic_vector(   0 downto 0);
        signal cVar1S20S7N050N044N056P038: std_logic_vector(   0 downto 0);
        signal cVar1S21S7N050N044N056P038: std_logic_vector(   0 downto 0);
        signal cVar1S22S7N050N044N056N038: std_logic_vector(   0 downto 0);
        signal cVar1S23S7N050N044N056N038: std_logic_vector(   0 downto 0);
        signal cVar1S24S7N050N044N056N038: std_logic_vector(   0 downto 0);
        signal cVar1S25S7N050N044N056N038: std_logic_vector(   0 downto 0);
        signal cVar1S0S8P044P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S8P044P023N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S8P044P023N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S8P044N023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S8P044N023N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S8P044N023N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S6S8P044N023N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S7S8P044N023N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S8S8N044P050P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S8N044P050P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S10S8N044P050P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S11S8N044P050P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S12S8N044P050N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S13S8N044P050N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S14S8N044P050N027P026: std_logic_vector(   0 downto 0);
        signal cVar1S15S8N044P050N027N026: std_logic_vector(   0 downto 0);
        signal cVar1S16S8N044P050N027N026: std_logic_vector(   0 downto 0);
        signal cVar1S17S8N044N050P014P051: std_logic_vector(   0 downto 0);
        signal cVar1S18S8N044N050P014P051: std_logic_vector(   0 downto 0);
        signal cVar1S19S8N044N050P014P051: std_logic_vector(   0 downto 0);
        signal cVar1S20S8N044N050P014N051: std_logic_vector(   0 downto 0);
        signal cVar1S21S8N044N050P014N051: std_logic_vector(   0 downto 0);
        signal cVar1S22S8N044N050P014N051: std_logic_vector(   0 downto 0);
        signal cVar1S23S8N044N050P014P032: std_logic_vector(   0 downto 0);
        signal cVar1S24S8N044N050P014P032: std_logic_vector(   0 downto 0);
        signal cVar1S25S8N044N050P014P032: std_logic_vector(   0 downto 0);
        signal cVar1S26S8N044N050P014N032: std_logic_vector(   0 downto 0);
        signal cVar1S27S8N044N050P014N032: std_logic_vector(   0 downto 0);
        signal cVar1S28S8N044N050P014N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S9P051P028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S9P051P028P055P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S9P051N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S9P051N028N029P026: std_logic_vector(   0 downto 0);
        signal cVar1S4S9P051N028N029P026: std_logic_vector(   0 downto 0);
        signal cVar1S5S9P051N028N029P026: std_logic_vector(   0 downto 0);
        signal cVar1S6S9P051N028N029N026: std_logic_vector(   0 downto 0);
        signal cVar1S7S9P051N028N029N026: std_logic_vector(   0 downto 0);
        signal cVar1S8S9N051P022P043P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S9N051P022N043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S9N051P022N043N004: std_logic_vector(   0 downto 0);
        signal cVar1S11S9N051N022P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S9N051N022P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S13S9N051N022P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S14S9N051N022P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S15S9N051N022N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S16S9N051N022N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S17S9N051N022N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S18S9N051N022N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S19S9N051N022N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S20S9N051N022N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S21S9N051N022N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S0S10P017P037P051P063: std_logic_vector(   0 downto 0);
        signal cVar1S1S10P017P037P051P063: std_logic_vector(   0 downto 0);
        signal cVar1S2S10P017P037P051P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S10P017P037N051P048: std_logic_vector(   0 downto 0);
        signal cVar1S4S10P017P037N051P048: std_logic_vector(   0 downto 0);
        signal cVar1S5S10P017P037N051P048: std_logic_vector(   0 downto 0);
        signal cVar1S6S10P017P037N051N048: std_logic_vector(   0 downto 0);
        signal cVar1S7S10P017P037N051N048: std_logic_vector(   0 downto 0);
        signal cVar1S8S10P017P037N051N048: std_logic_vector(   0 downto 0);
        signal cVar1S9S10P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S10S10P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S11S10P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S10P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S10P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S10P017P037N019P063: std_logic_vector(   0 downto 0);
        signal cVar1S15S10P017P037N019P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S10P017P064P019P068: std_logic_vector(   0 downto 0);
        signal cVar1S17S10P017P064P019P068: std_logic_vector(   0 downto 0);
        signal cVar1S18S10P017P064P019P068: std_logic_vector(   0 downto 0);
        signal cVar1S19S10P017P064P019P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S10P017P064P019P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S10P017P064P019P015: std_logic_vector(   0 downto 0);
        signal cVar1S22S10P017P064P019N015: std_logic_vector(   0 downto 0);
        signal cVar1S23S10P017N064P015P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S10P017N064P015P065: std_logic_vector(   0 downto 0);
        signal cVar1S25S10P017N064P015P065: std_logic_vector(   0 downto 0);
        signal cVar1S26S10P017N064P015P065: std_logic_vector(   0 downto 0);
        signal cVar1S27S10P017N064N015P037: std_logic_vector(   0 downto 0);
        signal cVar1S28S10P017N064N015P037: std_logic_vector(   0 downto 0);
        signal cVar1S29S10P017N064N015P037: std_logic_vector(   0 downto 0);
        signal cVar1S30S10P017N064N015P037: std_logic_vector(   0 downto 0);
        signal cVar1S31S10P017N064N015N037: std_logic_vector(   0 downto 0);
        signal cVar1S32S10P017N064N015N037: std_logic_vector(   0 downto 0);
        signal cVar1S33S10P017N064N015N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S11P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S11P048P025N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S11P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S3S11P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S11P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S11P048N025P027P011: std_logic_vector(   0 downto 0);
        signal cVar1S6S11P048N025P027P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S11P048N025P027P011: std_logic_vector(   0 downto 0);
        signal cVar1S8S11P048N025P027P011: std_logic_vector(   0 downto 0);
        signal cVar1S9S11P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S10S11P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S11S11P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S12S11P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S13S11N048P051P028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S11N048P051N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S11N048P051N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S16S11N048P051N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S17S11N048P051N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S18S11N048N051P022P043: std_logic_vector(   0 downto 0);
        signal cVar1S19S11N048N051P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S20S11N048N051P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S21S11N048N051P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S22S11N048N051N022P023: std_logic_vector(   0 downto 0);
        signal cVar1S23S11N048N051N022P023: std_logic_vector(   0 downto 0);
        signal cVar1S24S11N048N051N022P023: std_logic_vector(   0 downto 0);
        signal cVar1S25S11N048N051N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S26S11N048N051N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S27S11N048N051N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S28S11N048N051N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S0S12P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S12P048P025N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S12P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S3S12P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S12P048P025N007N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S12P048N025P027P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S12P048N025N027P067: std_logic_vector(   0 downto 0);
        signal cVar1S7S12P048N025N027P067: std_logic_vector(   0 downto 0);
        signal cVar1S8S12P048N025N027P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S12N048P001P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S12N048P001P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S11S12N048P001P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S12N048P001P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S12N048P001P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S12N048P001N051P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S12N048P001N051P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S12N048P001N051P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S12N048P001N051P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S12N048P001N051P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S12N048P001P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S12N048P001N041P017: std_logic_vector(   0 downto 0);
        signal cVar1S21S12N048P001N041P017: std_logic_vector(   0 downto 0);
        signal cVar1S22S12N048P001N041N017: std_logic_vector(   0 downto 0);
        signal cVar1S0S13P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S13P048P025N007P016nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S13P048N025P027P011nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S13P048N025P027P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S13P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S5S13P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S6S13P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S7S13P048N025N027P007: std_logic_vector(   0 downto 0);
        signal cVar1S8S13N048P051P008P013: std_logic_vector(   0 downto 0);
        signal cVar1S9S13N048P051P008P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S13N048P051N008P028: std_logic_vector(   0 downto 0);
        signal cVar1S11S13N048P051N008P028: std_logic_vector(   0 downto 0);
        signal cVar1S12S13N048P051N008P028: std_logic_vector(   0 downto 0);
        signal cVar1S13S13N048P051N008P028: std_logic_vector(   0 downto 0);
        signal cVar1S14S13N048P051N008N028: std_logic_vector(   0 downto 0);
        signal cVar1S15S13N048P051N008N028: std_logic_vector(   0 downto 0);
        signal cVar1S16S13N048P051N008N028: std_logic_vector(   0 downto 0);
        signal cVar1S17S13N048N051P038P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S13N048N051P038N021: std_logic_vector(   0 downto 0);
        signal cVar1S19S13N048N051P038N021: std_logic_vector(   0 downto 0);
        signal cVar1S20S13N048N051P038N021: std_logic_vector(   0 downto 0);
        signal cVar1S21S13N048N051N038P061: std_logic_vector(   0 downto 0);
        signal cVar1S22S13N048N051N038P061: std_logic_vector(   0 downto 0);
        signal cVar1S23S13N048N051N038P061: std_logic_vector(   0 downto 0);
        signal cVar1S24S13N048N051N038N061: std_logic_vector(   0 downto 0);
        signal cVar1S25S13N048N051N038N061: std_logic_vector(   0 downto 0);
        signal cVar1S26S13N048N051N038N061: std_logic_vector(   0 downto 0);
        signal cVar1S27S13N048N051N038N061: std_logic_vector(   0 downto 0);
        signal cVar1S0S14P017P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S14P017P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S14P017P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S14P017P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S4S14P017P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S14P017P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S6S14P017N048P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S14P017N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S8S14P017N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S9S14P017N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S10S14P017N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S11S14P017N048N044P038: std_logic_vector(   0 downto 0);
        signal cVar1S12S14P017N048N044P038: std_logic_vector(   0 downto 0);
        signal cVar1S13S14P017N048N044P038: std_logic_vector(   0 downto 0);
        signal cVar1S14S14P017N048N044N038: std_logic_vector(   0 downto 0);
        signal cVar1S15S14P017N048N044N038: std_logic_vector(   0 downto 0);
        signal cVar1S16S14P017P064P019P009: std_logic_vector(   0 downto 0);
        signal cVar1S17S14P017P064P019P009: std_logic_vector(   0 downto 0);
        signal cVar1S18S14P017P064P019P009: std_logic_vector(   0 downto 0);
        signal cVar1S19S14P017P064P019P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S14P017P064P019N050: std_logic_vector(   0 downto 0);
        signal cVar1S21S14P017P064P019N050: std_logic_vector(   0 downto 0);
        signal cVar1S22S14P017N064P061P003: std_logic_vector(   0 downto 0);
        signal cVar1S23S14P017N064P061P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S14P017N064P061P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S14P017N064P061P003: std_logic_vector(   0 downto 0);
        signal cVar1S26S14P017N064N061P051: std_logic_vector(   0 downto 0);
        signal cVar1S27S14P017N064N061P051: std_logic_vector(   0 downto 0);
        signal cVar1S28S14P017N064N061P051: std_logic_vector(   0 downto 0);
        signal cVar1S29S14P017N064N061N051: std_logic_vector(   0 downto 0);
        signal cVar1S30S14P017N064N061N051: std_logic_vector(   0 downto 0);
        signal cVar1S0S15P044P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S15P044P023N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S15P044P023N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S15P044P023N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S15P044N023P022P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S15P044N023N022P025: std_logic_vector(   0 downto 0);
        signal cVar1S6S15P044N023N022P025: std_logic_vector(   0 downto 0);
        signal cVar1S7S15P044N023N022P025: std_logic_vector(   0 downto 0);
        signal cVar1S8S15P044N023N022N025: std_logic_vector(   0 downto 0);
        signal cVar1S9S15P044N023N022N025: std_logic_vector(   0 downto 0);
        signal cVar1S10S15N044P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S15N044P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S12S15N044P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S13S15N044P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S14S15N044P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S15S15N044P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S16S15N044P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S17S15N044P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S18S15N044P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S19S15N044N048P007P040: std_logic_vector(   0 downto 0);
        signal cVar1S20S15N044N048P007P040: std_logic_vector(   0 downto 0);
        signal cVar1S21S15N044N048P007P040: std_logic_vector(   0 downto 0);
        signal cVar1S22S15N044N048P007N040: std_logic_vector(   0 downto 0);
        signal cVar1S23S15N044N048P007N040: std_logic_vector(   0 downto 0);
        signal cVar1S24S15N044N048P007N040: std_logic_vector(   0 downto 0);
        signal cVar1S25S15N044N048P007P043: std_logic_vector(   0 downto 0);
        signal cVar1S26S15N044N048P007P043: std_logic_vector(   0 downto 0);
        signal cVar1S27S15N044N048P007P043: std_logic_vector(   0 downto 0);
        signal cVar1S28S15N044N048P007N043: std_logic_vector(   0 downto 0);
        signal cVar1S29S15N044N048P007N043: std_logic_vector(   0 downto 0);
        signal cVar1S0S16P067P048P025P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S16P067P048N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S16P067P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S3S16P067P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S4S16P067P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S16P067N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S6S16P067N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S7S16P067N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S8S16P067N048P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S9S16P067N048P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S10S16P067N048N051P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S16P067N048N051P022: std_logic_vector(   0 downto 0);
        signal cVar1S12S16P067N048N051P022: std_logic_vector(   0 downto 0);
        signal cVar1S13S16P067N048N051N022: std_logic_vector(   0 downto 0);
        signal cVar1S14S16P067N048N051N022: std_logic_vector(   0 downto 0);
        signal cVar1S15S16P067N048N051N022: std_logic_vector(   0 downto 0);
        signal cVar1S16S16P067N048N051N022: std_logic_vector(   0 downto 0);
        signal cVar1S17S16P067P069P018P010: std_logic_vector(   0 downto 0);
        signal cVar1S18S16P067P069P018P010: std_logic_vector(   0 downto 0);
        signal cVar1S19S16P067P069P018P010: std_logic_vector(   0 downto 0);
        signal cVar1S20S16P067P069P018P010: std_logic_vector(   0 downto 0);
        signal cVar1S21S16P067P069N018P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S16P067P069N018P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S16P067P069N018P019: std_logic_vector(   0 downto 0);
        signal cVar1S24S16P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S25S16P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S26S16P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S27S16P067N069P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S16P067N069N052P065: std_logic_vector(   0 downto 0);
        signal cVar1S29S16P067N069N052P065: std_logic_vector(   0 downto 0);
        signal cVar1S30S16P067N069N052N065: std_logic_vector(   0 downto 0);
        signal cVar1S0S17P022P043P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S17P022N043P069P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S17P022N043P069N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S17P022N043P069N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S17N022P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S17N022P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S17N022P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S17N022P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S8S17N022P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S9S17N022P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S10S17N022P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S17N022P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S12S17N022N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S13S17N022N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S14S17N022N048P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S17N022N048P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S16S17N022N048P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S17S17N022N048P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S18S17N022N048N051P038: std_logic_vector(   0 downto 0);
        signal cVar1S19S17N022N048N051P038: std_logic_vector(   0 downto 0);
        signal cVar1S20S17N022N048N051P038: std_logic_vector(   0 downto 0);
        signal cVar1S21S17N022N048N051N038: std_logic_vector(   0 downto 0);
        signal cVar1S22S17N022N048N051N038: std_logic_vector(   0 downto 0);
        signal cVar1S23S17N022N048N051N038: std_logic_vector(   0 downto 0);
        signal cVar1S24S17N022N048N051N038: std_logic_vector(   0 downto 0);
        signal cVar1S0S18P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S18P041N020P021P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S18P041N020N021P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S18P041N020N021P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S18P041N020N021N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S18P041N020N021N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S18N041P039P020P044: std_logic_vector(   0 downto 0);
        signal cVar1S7S18N041P039P020P044: std_logic_vector(   0 downto 0);
        signal cVar1S8S18N041P039P020P044: std_logic_vector(   0 downto 0);
        signal cVar1S9S18N041P039P020N044: std_logic_vector(   0 downto 0);
        signal cVar1S10S18N041P039P020N044: std_logic_vector(   0 downto 0);
        signal cVar1S11S18N041P039P020N044: std_logic_vector(   0 downto 0);
        signal cVar1S12S18N041P039P020N044: std_logic_vector(   0 downto 0);
        signal cVar1S13S18N041P039P020P040: std_logic_vector(   0 downto 0);
        signal cVar1S14S18N041P039P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S15S18N041P039P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S16S18N041P039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S18N041P039N005P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S18N041P039N005N020: std_logic_vector(   0 downto 0);
        signal cVar1S0S19P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S19P041N020P021P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S19P041N020P021N003: std_logic_vector(   0 downto 0);
        signal cVar1S3S19P041N020N021P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S19P041N020N021P022: std_logic_vector(   0 downto 0);
        signal cVar1S5S19P041N020N021N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S19P041N020N021N022: std_logic_vector(   0 downto 0);
        signal cVar1S7S19P041N020N021N022: std_logic_vector(   0 downto 0);
        signal cVar1S8S19N041P039P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S9S19N041P039P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S10S19N041P039P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S11S19N041P039P044N023psss: std_logic_vector(   0 downto 0);
        signal cVar1S12S19N041P039N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S13S19N041P039N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S14S19N041P039N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S15S19N041P039N044P050: std_logic_vector(   0 downto 0);
        signal cVar1S16S19N041P039N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S17S19N041P039N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S18S19N041P039N044N050: std_logic_vector(   0 downto 0);
        signal cVar1S19S19N041P039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S19N041P039N005N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S20P011P029P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S1S20P011P029P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S2S20P011P029P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S3S20P011P029P048N025psss: std_logic_vector(   0 downto 0);
        signal cVar1S4S20P011P029N048P041: std_logic_vector(   0 downto 0);
        signal cVar1S5S20P011P029N048P041: std_logic_vector(   0 downto 0);
        signal cVar1S6S20P011P029N048P041: std_logic_vector(   0 downto 0);
        signal cVar1S7S20P011P029N048N041: std_logic_vector(   0 downto 0);
        signal cVar1S8S20P011P029N048N041: std_logic_vector(   0 downto 0);
        signal cVar1S9S20P011P029N048N041: std_logic_vector(   0 downto 0);
        signal cVar1S10S20P011P029N048N041: std_logic_vector(   0 downto 0);
        signal cVar1S11S20P011P029P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S20P011P029P010N052: std_logic_vector(   0 downto 0);
        signal cVar1S13S20P011P029N010P009: std_logic_vector(   0 downto 0);
        signal cVar1S14S20P011P029N010P009: std_logic_vector(   0 downto 0);
        signal cVar1S15S20P011P029N010N009: std_logic_vector(   0 downto 0);
        signal cVar1S16S20P011P029P060P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S20P011P029P060P014: std_logic_vector(   0 downto 0);
        signal cVar1S18S20P011P029P060P014: std_logic_vector(   0 downto 0);
        signal cVar1S19S20P011P029P060P014: std_logic_vector(   0 downto 0);
        signal cVar1S20S20P011N029P015P033: std_logic_vector(   0 downto 0);
        signal cVar1S21S20P011N029P015P033: std_logic_vector(   0 downto 0);
        signal cVar1S22S20P011N029P015P033: std_logic_vector(   0 downto 0);
        signal cVar1S23S20P011N029P015P033: std_logic_vector(   0 downto 0);
        signal cVar1S24S20P011N029N015P017: std_logic_vector(   0 downto 0);
        signal cVar1S25S20P011N029N015P017: std_logic_vector(   0 downto 0);
        signal cVar1S26S20P011N029N015P017: std_logic_vector(   0 downto 0);
        signal cVar1S27S20P011N029N015N017: std_logic_vector(   0 downto 0);
        signal cVar1S28S20P011N029N015N017: std_logic_vector(   0 downto 0);
        signal cVar1S0S21P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S21P041N020P021P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S21P041N020P021N003: std_logic_vector(   0 downto 0);
        signal cVar1S3S21P041N020N021P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S21P041N020N021N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S21P041N020N021N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S21P041N020N021N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S21N041P039P000P048: std_logic_vector(   0 downto 0);
        signal cVar1S8S21N041P039P000P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S21N041P039P000P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S21N041P039P000N048: std_logic_vector(   0 downto 0);
        signal cVar1S11S21N041P039P000N048: std_logic_vector(   0 downto 0);
        signal cVar1S12S21N041P039P000N048: std_logic_vector(   0 downto 0);
        signal cVar1S13S21N041P039P000P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S21N041P039P000N040: std_logic_vector(   0 downto 0);
        signal cVar1S15S21N041P039P000N040: std_logic_vector(   0 downto 0);
        signal cVar1S16S21N041P039P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S21N041P039N051P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S22P000P041P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S22P000P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S2S22P000P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S3S22P000P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S4S22P000P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S5S22P000P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S6S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S7S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S8S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S9S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S10S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S11S22P000N041P039P012: std_logic_vector(   0 downto 0);
        signal cVar1S12S22P000N041P039P049nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S22P000N041P039N049: std_logic_vector(   0 downto 0);
        signal cVar1S14S22P000N041P039N049: std_logic_vector(   0 downto 0);
        signal cVar1S15S22P000N041P039N049: std_logic_vector(   0 downto 0);
        signal cVar1S16S22P000P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S22P000N040P059P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S22P000N040P059N041: std_logic_vector(   0 downto 0);
        signal cVar1S19S22P000N040P059N041: std_logic_vector(   0 downto 0);
        signal cVar1S0S23P041P020P010nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S23P041N020P005P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S23P041N020P005N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S23P041N020P005N021: std_logic_vector(   0 downto 0);
        signal cVar1S4S23P041N020N005P003: std_logic_vector(   0 downto 0);
        signal cVar1S5S23P041N020N005N003: std_logic_vector(   0 downto 0);
        signal cVar1S6S23N041P055P061P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S23N041P055P061P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S23N041P055P061P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S23N041P055P061P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S23N041P055P061P054nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S23N041P055P061N054: std_logic_vector(   0 downto 0);
        signal cVar1S12S23N041N055P010P039: std_logic_vector(   0 downto 0);
        signal cVar1S13S23N041N055P010P039: std_logic_vector(   0 downto 0);
        signal cVar1S14S23N041N055P010P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S23N041N055P010P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S23N041N055P010P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S23N041N055P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S18S23N041N055P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S19S23N041N055P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S0S24P041P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S24P041N020P005P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S24P041N020P005N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S24P041N020P005N021: std_logic_vector(   0 downto 0);
        signal cVar1S4S24P041N020N005P003: std_logic_vector(   0 downto 0);
        signal cVar1S5S24P041N020N005N003: std_logic_vector(   0 downto 0);
        signal cVar1S6S24P041N020N005N003: std_logic_vector(   0 downto 0);
        signal cVar1S7S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S8S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S9S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S10S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S11S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S12S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S13S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S14S24N041P039P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S15S24N041P039P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S16S24N041P039P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S17S24N041P039P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S18S24N041P039P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S24N041P039N051P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S24N041P039N051N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S25P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S25P041N020P005P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S25P041N020P005N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S25P041N020N005P003: std_logic_vector(   0 downto 0);
        signal cVar1S4S25P041N020N005N003: std_logic_vector(   0 downto 0);
        signal cVar1S5S25P041N020N005N003: std_logic_vector(   0 downto 0);
        signal cVar1S6S25N041P013P031P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S25N041P013P031P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S25N041P013P031N056: std_logic_vector(   0 downto 0);
        signal cVar1S9S25N041P013P031N056: std_logic_vector(   0 downto 0);
        signal cVar1S10S25N041P013N031P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S25N041P013N031P015: std_logic_vector(   0 downto 0);
        signal cVar1S12S25N041P013N031P015: std_logic_vector(   0 downto 0);
        signal cVar1S13S25N041P013N031N015: std_logic_vector(   0 downto 0);
        signal cVar1S14S25N041P013N031N015: std_logic_vector(   0 downto 0);
        signal cVar1S15S25N041N013P031P044: std_logic_vector(   0 downto 0);
        signal cVar1S16S25N041N013P031P044: std_logic_vector(   0 downto 0);
        signal cVar1S17S25N041N013P031N044: std_logic_vector(   0 downto 0);
        signal cVar1S18S25N041N013P031N044: std_logic_vector(   0 downto 0);
        signal cVar1S19S25N041N013P031N044: std_logic_vector(   0 downto 0);
        signal cVar1S20S25N041N013P031P011: std_logic_vector(   0 downto 0);
        signal cVar1S21S25N041N013P031P011: std_logic_vector(   0 downto 0);
        signal cVar1S22S25N041N013P031N011: std_logic_vector(   0 downto 0);
        signal cVar1S0S26P068P041P020P016nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S26P068P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S2S26P068P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S3S26P068P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S4S26P068P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S5S26P068N041P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S6S26P068N041P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S7S26P068N041P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S8S26P068N041P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S9S26P068N041P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S10S26P068N041N024P023: std_logic_vector(   0 downto 0);
        signal cVar1S11S26P068N041N024P023: std_logic_vector(   0 downto 0);
        signal cVar1S12S26P068N041N024P023: std_logic_vector(   0 downto 0);
        signal cVar1S13S26P068N041N024P023: std_logic_vector(   0 downto 0);
        signal cVar1S14S26P068N041N024N023: std_logic_vector(   0 downto 0);
        signal cVar1S15S26P068N041N024N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S26P068N041N024N023: std_logic_vector(   0 downto 0);
        signal cVar1S17S26P068P065P019P061: std_logic_vector(   0 downto 0);
        signal cVar1S18S26P068P065P019P061: std_logic_vector(   0 downto 0);
        signal cVar1S19S26P068P065N019P037: std_logic_vector(   0 downto 0);
        signal cVar1S20S26P068P065N019P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S26P068P065N019P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S26P068P065N019N037: std_logic_vector(   0 downto 0);
        signal cVar1S23S26P068P065N019N037: std_logic_vector(   0 downto 0);
        signal cVar1S24S26P068P065N019N037: std_logic_vector(   0 downto 0);
        signal cVar1S25S26P068P065P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S26S26P068P065P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S27S26P068P065P069P036: std_logic_vector(   0 downto 0);
        signal cVar1S28S26P068P065N069P016: std_logic_vector(   0 downto 0);
        signal cVar1S29S26P068P065N069P016: std_logic_vector(   0 downto 0);
        signal cVar1S30S26P068P065N069N016: std_logic_vector(   0 downto 0);
        signal cVar1S31S26P068P065N069N016: std_logic_vector(   0 downto 0);
        signal cVar1S0S27P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S27P041P020N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S27P041P020N003N002: std_logic_vector(   0 downto 0);
        signal cVar1S3S27P041P020N003N002: std_logic_vector(   0 downto 0);
        signal cVar1S4S27P041N020P068P005: std_logic_vector(   0 downto 0);
        signal cVar1S5S27P041N020P068P005: std_logic_vector(   0 downto 0);
        signal cVar1S6S27P041N020P068N005: std_logic_vector(   0 downto 0);
        signal cVar1S7S27P041N020P068P039: std_logic_vector(   0 downto 0);
        signal cVar1S8S27N041P024P006P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S27N041P024P006N047: std_logic_vector(   0 downto 0);
        signal cVar1S10S27N041P024P006N047: std_logic_vector(   0 downto 0);
        signal cVar1S11S27N041P024P006N047: std_logic_vector(   0 downto 0);
        signal cVar1S12S27N041P024N006P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S27N041P024N006P049: std_logic_vector(   0 downto 0);
        signal cVar1S14S27N041P024N006N049: std_logic_vector(   0 downto 0);
        signal cVar1S15S27N041P024N006N049: std_logic_vector(   0 downto 0);
        signal cVar1S16S27N041N024P023P005: std_logic_vector(   0 downto 0);
        signal cVar1S17S27N041N024P023P005: std_logic_vector(   0 downto 0);
        signal cVar1S18S27N041N024P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S19S27N041N024P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S20S27N041N024P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S21S27N041N024P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S22S27N041N024N023P050: std_logic_vector(   0 downto 0);
        signal cVar1S23S27N041N024N023P050: std_logic_vector(   0 downto 0);
        signal cVar1S24S27N041N024N023P050: std_logic_vector(   0 downto 0);
        signal cVar1S25S27N041N024N023P050: std_logic_vector(   0 downto 0);
        signal cVar1S26S27N041N024N023N050: std_logic_vector(   0 downto 0);
        signal cVar1S27S27N041N024N023N050: std_logic_vector(   0 downto 0);
        signal cVar1S28S27N041N024N023N050: std_logic_vector(   0 downto 0);
        signal cVar1S0S28P024P006P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S28P024P006N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S28P024P006N047N045: std_logic_vector(   0 downto 0);
        signal cVar1S3S28P024P006N047N045: std_logic_vector(   0 downto 0);
        signal cVar1S4S28P024N006P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S5S28P024N006P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S6S28P024N006P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S7S28P024N006P068P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S28N024P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S28N024P040N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S28N024P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S11S28N024P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S12S28N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S13S28N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S14S28N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S28N024N040P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S28N024N040P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S17S28N024N040P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S18S28N024N040N044P042: std_logic_vector(   0 downto 0);
        signal cVar1S19S28N024N040N044P042: std_logic_vector(   0 downto 0);
        signal cVar1S20S28N024N040N044P042: std_logic_vector(   0 downto 0);
        signal cVar1S21S28N024N040N044P042: std_logic_vector(   0 downto 0);
        signal cVar1S22S28N024N040N044P042: std_logic_vector(   0 downto 0);
        signal cVar1S0S29P024P006P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S29P024P006N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S29P024P006N047N045: std_logic_vector(   0 downto 0);
        signal cVar1S3S29P024P006N047N045: std_logic_vector(   0 downto 0);
        signal cVar1S4S29P024N006P068P007: std_logic_vector(   0 downto 0);
        signal cVar1S5S29P024N006P068P007: std_logic_vector(   0 downto 0);
        signal cVar1S6S29P024N006P068N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S29P024N006P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S29P024N006P068N012: std_logic_vector(   0 downto 0);
        signal cVar1S9S29N024P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S29N024P040N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S29N024P040N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S29N024P040N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S13S29N024P040N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S14S29N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S29N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S29N024N040P044P023: std_logic_vector(   0 downto 0);
        signal cVar1S17S29N024N040P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S18S29N024N040P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S19S29N024N040N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S20S29N024N040N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S21S29N024N040N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S22S29N024N040N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S23S29N024N040N044N041: std_logic_vector(   0 downto 0);
        signal cVar1S0S30P067P018P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S30P067P018P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S2S30P067P018P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S30P067P018P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S30P067P018N048P014: std_logic_vector(   0 downto 0);
        signal cVar1S5S30P067P018N048P014: std_logic_vector(   0 downto 0);
        signal cVar1S6S30P067P018N048P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S30P067P018N048P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S30P067P018N048N014: std_logic_vector(   0 downto 0);
        signal cVar1S9S30P067P018N048N014: std_logic_vector(   0 downto 0);
        signal cVar1S10S30P067P018P060P011: std_logic_vector(   0 downto 0);
        signal cVar1S11S30P067P018P060P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S30P067P018P060P011: std_logic_vector(   0 downto 0);
        signal cVar1S13S30P067P018P060N011: std_logic_vector(   0 downto 0);
        signal cVar1S14S30P067P018P060N011: std_logic_vector(   0 downto 0);
        signal cVar1S15S30P067P018P060N011: std_logic_vector(   0 downto 0);
        signal cVar1S16S30P067P018P060P013: std_logic_vector(   0 downto 0);
        signal cVar1S17S30P067P018P060P013: std_logic_vector(   0 downto 0);
        signal cVar1S18S30P067P018P060N013: std_logic_vector(   0 downto 0);
        signal cVar1S19S30P067P018P060N013: std_logic_vector(   0 downto 0);
        signal cVar1S20S30P067P069P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S21S30P067P069P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S22S30P067P069P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S23S30P067P069P018P016: std_logic_vector(   0 downto 0);
        signal cVar1S24S30P067P069N018P019: std_logic_vector(   0 downto 0);
        signal cVar1S25S30P067P069N018P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S30P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S27S30P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S28S30P067P069N018N019: std_logic_vector(   0 downto 0);
        signal cVar1S29S30P067N069P065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S30P067N069P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S31S30P067N069N065P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S32S30P067N069N065N052: std_logic_vector(   0 downto 0);
        signal cVar1S0S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S3S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S4S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S5S31P018P060P054P062: std_logic_vector(   0 downto 0);
        signal cVar1S6S31P018P060P054P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S31P018P060P054N011: std_logic_vector(   0 downto 0);
        signal cVar1S8S31P018P060P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S31P018P060P029N050: std_logic_vector(   0 downto 0);
        signal cVar1S10S31P018P060P029N050: std_logic_vector(   0 downto 0);
        signal cVar1S11S31N018P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S31N018P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S13S31N018P048P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S14S31N018P048N025P036nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S31N018N048P014P034: std_logic_vector(   0 downto 0);
        signal cVar1S16S31N018N048P014N034: std_logic_vector(   0 downto 0);
        signal cVar1S17S31N018N048P014N034: std_logic_vector(   0 downto 0);
        signal cVar1S18S31N018N048P014N034: std_logic_vector(   0 downto 0);
        signal cVar1S19S31N018N048N014P030: std_logic_vector(   0 downto 0);
        signal cVar1S20S31N018N048N014P030: std_logic_vector(   0 downto 0);
        signal cVar1S21S31N018N048N014P030: std_logic_vector(   0 downto 0);
        signal cVar1S22S31N018N048N014P030: std_logic_vector(   0 downto 0);
        signal cVar1S23S31N018N048N014N030: std_logic_vector(   0 downto 0);
        signal cVar1S24S31N018N048N014N030: std_logic_vector(   0 downto 0);
        signal cVar1S25S31N018N048N014N030: std_logic_vector(   0 downto 0);
        signal cVar1S26S31N018N048N014N030: std_logic_vector(   0 downto 0);
        signal cVar1S0S32P015P018P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S32P015P018P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S2S32P015P018P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S32P015P018P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S4S32P015P018N040P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S32P015P018N040P063: std_logic_vector(   0 downto 0);
        signal cVar1S6S32P015P018N040P063: std_logic_vector(   0 downto 0);
        signal cVar1S7S32P015P018N040P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S32P015P018N040N063: std_logic_vector(   0 downto 0);
        signal cVar1S9S32P015P018N040N063: std_logic_vector(   0 downto 0);
        signal cVar1S10S32P015P018N040N063: std_logic_vector(   0 downto 0);
        signal cVar1S11S32P015P018N040N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S15S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S16S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S17S32P015P018P004P062: std_logic_vector(   0 downto 0);
        signal cVar1S18S32P015P018P004P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S32P015P018P004N041: std_logic_vector(   0 downto 0);
        signal cVar1S20S32P015P018P004N041: std_logic_vector(   0 downto 0);
        signal cVar1S21S32P015P018P004N041: std_logic_vector(   0 downto 0);
        signal cVar1S22S32P015P017P060P063: std_logic_vector(   0 downto 0);
        signal cVar1S23S32P015P017P060P063: std_logic_vector(   0 downto 0);
        signal cVar1S24S32P015P017P060P063: std_logic_vector(   0 downto 0);
        signal cVar1S25S32P015P017P060P063: std_logic_vector(   0 downto 0);
        signal cVar1S26S32P015P017N060P018: std_logic_vector(   0 downto 0);
        signal cVar1S27S32P015P017N060P018: std_logic_vector(   0 downto 0);
        signal cVar1S28S32P015P017N060N018: std_logic_vector(   0 downto 0);
        signal cVar1S29S32P015P017N060N018: std_logic_vector(   0 downto 0);
        signal cVar1S30S32P015P017N060N018: std_logic_vector(   0 downto 0);
        signal cVar1S31S32P015P017N060N018: std_logic_vector(   0 downto 0);
        signal cVar1S32S32P015P017P008P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S33S32P015P017P008P066: std_logic_vector(   0 downto 0);
        signal cVar1S34S32P015P017N008P056: std_logic_vector(   0 downto 0);
        signal cVar1S35S32P015P017N008P056: std_logic_vector(   0 downto 0);
        signal cVar1S36S32P015P017N008P056: std_logic_vector(   0 downto 0);
        signal cVar1S0S33P016P063P056P059: std_logic_vector(   0 downto 0);
        signal cVar1S1S33P016P063P056P059: std_logic_vector(   0 downto 0);
        signal cVar1S2S33P016P063P056P059: std_logic_vector(   0 downto 0);
        signal cVar1S3S33P016P063P056P059: std_logic_vector(   0 downto 0);
        signal cVar1S4S33P016P063P056P059: std_logic_vector(   0 downto 0);
        signal cVar1S5S33P016P063P056P062: std_logic_vector(   0 downto 0);
        signal cVar1S6S33P016N063P059P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S33P016N063P059P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S33P016N063P059P014: std_logic_vector(   0 downto 0);
        signal cVar1S9S33P016N063P059N014: std_logic_vector(   0 downto 0);
        signal cVar1S10S33P016N063P059N014: std_logic_vector(   0 downto 0);
        signal cVar1S11S33P016N063P059N014: std_logic_vector(   0 downto 0);
        signal cVar1S12S33P016N063P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S33P016N063P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S33P016N063P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S15S33P016N063P059N032: std_logic_vector(   0 downto 0);
        signal cVar1S16S33N016P034P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S17S33N016P034P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S18S33N016P034P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S19S33N016P034P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S20S33N016P034P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S21S33N016P034N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S22S33N016P034N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S23S33N016P034N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S24S33N016P034N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S25S33N016P034N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S26S33N016P034N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S27S33N016P034N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S28S33N016P034P014P053: std_logic_vector(   0 downto 0);
        signal cVar1S29S33N016P034P014P053: std_logic_vector(   0 downto 0);
        signal cVar1S30S33N016P034P014P053: std_logic_vector(   0 downto 0);
        signal cVar1S31S33N016P034N014P017: std_logic_vector(   0 downto 0);
        signal cVar1S0S34P067P062P008P049: std_logic_vector(   0 downto 0);
        signal cVar1S1S34P067P062P008P049: std_logic_vector(   0 downto 0);
        signal cVar1S2S34P067P062P008N049: std_logic_vector(   0 downto 0);
        signal cVar1S3S34P067P062P008N049: std_logic_vector(   0 downto 0);
        signal cVar1S4S34P067P062P008N049: std_logic_vector(   0 downto 0);
        signal cVar1S5S34P067P062P008N049: std_logic_vector(   0 downto 0);
        signal cVar1S6S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S7S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S8S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S9S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S10S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S11S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S12S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S13S34P067P062N008P035: std_logic_vector(   0 downto 0);
        signal cVar1S14S34P067P062P055P035: std_logic_vector(   0 downto 0);
        signal cVar1S15S34P067P062P055P035: std_logic_vector(   0 downto 0);
        signal cVar1S16S34P067P062P055P035: std_logic_vector(   0 downto 0);
        signal cVar1S17S34P067P062P055N035: std_logic_vector(   0 downto 0);
        signal cVar1S18S34P067P062P055N035: std_logic_vector(   0 downto 0);
        signal cVar1S19S34P067P062P055N035: std_logic_vector(   0 downto 0);
        signal cVar1S20S34P067P062P055P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S34P067P010P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S22S34P067P010P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S23S34P067P010P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S24S34P067P010P069P031: std_logic_vector(   0 downto 0);
        signal cVar1S25S34P067P010N069P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S34P067P010P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S27S34P067P010P015P036: std_logic_vector(   0 downto 0);
        signal cVar1S28S34P067P010N015P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S29S34P067P010N015N050: std_logic_vector(   0 downto 0);
        signal cVar1S0S35P058P035P013P066: std_logic_vector(   0 downto 0);
        signal cVar1S1S35P058P035P013P066: std_logic_vector(   0 downto 0);
        signal cVar1S2S35P058P035P013P066: std_logic_vector(   0 downto 0);
        signal cVar1S3S35P058P035P013P066: std_logic_vector(   0 downto 0);
        signal cVar1S4S35P058P035N013P004: std_logic_vector(   0 downto 0);
        signal cVar1S5S35P058P035N013P004: std_logic_vector(   0 downto 0);
        signal cVar1S6S35P058P035N013P004: std_logic_vector(   0 downto 0);
        signal cVar1S7S35P058P035P060P034: std_logic_vector(   0 downto 0);
        signal cVar1S8S35N058P030P012P031: std_logic_vector(   0 downto 0);
        signal cVar1S9S35N058P030P012P031: std_logic_vector(   0 downto 0);
        signal cVar1S10S35N058P030P012P031: std_logic_vector(   0 downto 0);
        signal cVar1S11S35N058P030N012P010: std_logic_vector(   0 downto 0);
        signal cVar1S12S35N058P030N012P010: std_logic_vector(   0 downto 0);
        signal cVar1S13S35N058P030N012N010: std_logic_vector(   0 downto 0);
        signal cVar1S14S35N058N030P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S15S35N058N030P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S16S35N058N030P024P006: std_logic_vector(   0 downto 0);
        signal cVar1S17S35N058N030P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S18S35N058N030P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S19S35N058N030N024P037: std_logic_vector(   0 downto 0);
        signal cVar1S20S35N058N030N024P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S35N058N030N024P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S35N058N030N024N037: std_logic_vector(   0 downto 0);
        signal cVar1S23S35N058N030N024N037: std_logic_vector(   0 downto 0);
        signal cVar1S24S35N058N030N024N037: std_logic_vector(   0 downto 0);
        signal cVar1S25S35N058N030N024N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S36P037P048P025P067nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S36P037P048N025P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S36P037P048N025P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S36P037P048N025N009: std_logic_vector(   0 downto 0);
        signal cVar1S4S36P037P048N025N009: std_logic_vector(   0 downto 0);
        signal cVar1S5S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S7S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S8S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S9S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S10S36P037N048P046P009: std_logic_vector(   0 downto 0);
        signal cVar1S11S36P037N048P046P044: std_logic_vector(   0 downto 0);
        signal cVar1S12S36P037N048P046P044: std_logic_vector(   0 downto 0);
        signal cVar1S13S36P037N048P046P044: std_logic_vector(   0 downto 0);
        signal cVar1S14S36P037N048P046P044: std_logic_vector(   0 downto 0);
        signal cVar1S15S36P037N048P046N044: std_logic_vector(   0 downto 0);
        signal cVar1S16S36P037P059P005P035: std_logic_vector(   0 downto 0);
        signal cVar1S17S36P037P059P005P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S36P037P059P005N035: std_logic_vector(   0 downto 0);
        signal cVar1S19S36P037P059P005N035: std_logic_vector(   0 downto 0);
        signal cVar1S20S36P037P059P005N035: std_logic_vector(   0 downto 0);
        signal cVar1S21S36P037P059P005P063: std_logic_vector(   0 downto 0);
        signal cVar1S22S36P037P059P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S36P037P059N008P060: std_logic_vector(   0 downto 0);
        signal cVar1S24S36P037P059N008N060: std_logic_vector(   0 downto 0);
        signal cVar1S0S37P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S37P048P025N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S37P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S37P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S37P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S37P048N025P037P017nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S37P048N025P037P017: std_logic_vector(   0 downto 0);
        signal cVar1S7S37P048N025P037P017: std_logic_vector(   0 downto 0);
        signal cVar1S8S37P048N025P037P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S37P048N025P037P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S37P048N025P037N006: std_logic_vector(   0 downto 0);
        signal cVar1S11S37N048P044P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S37N048P044N004P005: std_logic_vector(   0 downto 0);
        signal cVar1S13S37N048P044N004P005: std_logic_vector(   0 downto 0);
        signal cVar1S14S37N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S15S37N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S16S37N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S17S37N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S18S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S19S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S20S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S21S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S22S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S23S37N048N044P046P025: std_logic_vector(   0 downto 0);
        signal cVar1S24S37N048N044P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S0S38P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S38P048P025N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S38P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S38P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S38P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S38P048N025P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S6S38P048N025P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S7S38P048N025P052P027: std_logic_vector(   0 downto 0);
        signal cVar1S8S38P048N025P052N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S38P048N025P052N027: std_logic_vector(   0 downto 0);
        signal cVar1S10S38P048N025P052N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S38P048N025P052P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S38P048N025P052N046: std_logic_vector(   0 downto 0);
        signal cVar1S13S38N048P025P046P018: std_logic_vector(   0 downto 0);
        signal cVar1S14S38N048P025P046P018: std_logic_vector(   0 downto 0);
        signal cVar1S15S38N048P025P046P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S38N048P025P046N018: std_logic_vector(   0 downto 0);
        signal cVar1S17S38N048P025P046N018: std_logic_vector(   0 downto 0);
        signal cVar1S18S38N048P025P046N018: std_logic_vector(   0 downto 0);
        signal cVar1S19S38N048P025P046N018: std_logic_vector(   0 downto 0);
        signal cVar1S20S38N048P025P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S21S38N048P025P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S22S38N048P025P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S23S38N048P025P007P009: std_logic_vector(   0 downto 0);
        signal cVar1S24S38N048P025P007P009: std_logic_vector(   0 downto 0);
        signal cVar1S25S38N048P025P007P009: std_logic_vector(   0 downto 0);
        signal cVar1S26S38N048P025N007P044: std_logic_vector(   0 downto 0);
        signal cVar1S27S38N048P025N007N044: std_logic_vector(   0 downto 0);
        signal cVar1S0S39P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S39P048P025N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S39P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S39P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S39P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S39P048N025P027P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S39P048N025P027N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S39P048N025P027N007: std_logic_vector(   0 downto 0);
        signal cVar1S8S39P048N025P027N007: std_logic_vector(   0 downto 0);
        signal cVar1S9S39P048N025N027P058nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S39P048N025N027N058: std_logic_vector(   0 downto 0);
        signal cVar1S11S39P048N025N027N058: std_logic_vector(   0 downto 0);
        signal cVar1S12S39P048N025N027N058: std_logic_vector(   0 downto 0);
        signal cVar1S13S39N048P044P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S39N048P044N004P005: std_logic_vector(   0 downto 0);
        signal cVar1S15S39N048P044N004P005: std_logic_vector(   0 downto 0);
        signal cVar1S16S39N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S17S39N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S18S39N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S19S39N048P044N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S20S39N048N044P046P052: std_logic_vector(   0 downto 0);
        signal cVar1S21S39N048N044P046P052: std_logic_vector(   0 downto 0);
        signal cVar1S22S39N048N044P046P052: std_logic_vector(   0 downto 0);
        signal cVar1S23S39N048N044P046P052: std_logic_vector(   0 downto 0);
        signal cVar1S24S39N048N044P046N052: std_logic_vector(   0 downto 0);
        signal cVar1S25S39N048N044P046N052: std_logic_vector(   0 downto 0);
        signal cVar1S26S39N048N044P046N052: std_logic_vector(   0 downto 0);
        signal cVar1S27S39N048N044P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S28S39N048N044P046P027: std_logic_vector(   0 downto 0);
        signal cVar1S0S40P018P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S40P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S40P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S40P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S4S40P018P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S40P018P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S6S40P018N048P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S7S40P018N048P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S8S40P018N048P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S9S40P018N048P010P032: std_logic_vector(   0 downto 0);
        signal cVar1S10S40P018N048P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S11S40P018N048P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S12S40P018N048P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S13S40P018N048P010N032: std_logic_vector(   0 downto 0);
        signal cVar1S14S40P018N048P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S15S40P018N048P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S16S40P018N048P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S17S40P018N048P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S18S40P018N048P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S19S40P018N048P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S20S40P018P069P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S21S40P018P069P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S22S40P018P069P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S23S40P018P069N009P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S40P018P069N009P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S40P018P069N009N003: std_logic_vector(   0 downto 0);
        signal cVar1S26S40P018P069N009N003: std_logic_vector(   0 downto 0);
        signal cVar1S27S40P018P069N009N003: std_logic_vector(   0 downto 0);
        signal cVar1S28S40P018P069N009N003: std_logic_vector(   0 downto 0);
        signal cVar1S29S40P018P069P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S41P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S41P048P025N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S41P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S41P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S41P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S41P048N025P052P065: std_logic_vector(   0 downto 0);
        signal cVar1S6S41P048N025P052P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S41P048N025P052P065: std_logic_vector(   0 downto 0);
        signal cVar1S8S41P048N025P052P065: std_logic_vector(   0 downto 0);
        signal cVar1S9S41P048N025P052P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S41P048N025P052N015: std_logic_vector(   0 downto 0);
        signal cVar1S11S41P048N025P052N015: std_logic_vector(   0 downto 0);
        signal cVar1S12S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S13S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S14S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S15S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S16S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S17S41N048P018P059P045: std_logic_vector(   0 downto 0);
        signal cVar1S18S41N048P018P059P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S41N048P018P059N050: std_logic_vector(   0 downto 0);
        signal cVar1S20S41N048P018P059N050: std_logic_vector(   0 downto 0);
        signal cVar1S21S41N048N018P032P028: std_logic_vector(   0 downto 0);
        signal cVar1S22S41N048N018P032P028: std_logic_vector(   0 downto 0);
        signal cVar1S23S41N048N018P032P028: std_logic_vector(   0 downto 0);
        signal cVar1S24S41N048N018N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S25S41N048N018N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S26S41N048N018N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S27S41N048N018N032P056: std_logic_vector(   0 downto 0);
        signal cVar1S28S41N048N018N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S29S41N048N018N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S30S41N048N018N032N056: std_logic_vector(   0 downto 0);
        signal cVar1S0S42P018P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S42P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S42P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S42P018P048N025P027: std_logic_vector(   0 downto 0);
        signal cVar1S4S42P018P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S42P018P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S6S42P018P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S7S42P018N048P038P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S42P018N048P038N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S42P018N048P038N002: std_logic_vector(   0 downto 0);
        signal cVar1S10S42P018N048N038P000: std_logic_vector(   0 downto 0);
        signal cVar1S11S42P018N048N038P000: std_logic_vector(   0 downto 0);
        signal cVar1S12S42P018N048N038P000: std_logic_vector(   0 downto 0);
        signal cVar1S13S42P018N048N038P000: std_logic_vector(   0 downto 0);
        signal cVar1S14S42P018N048N038P000: std_logic_vector(   0 downto 0);
        signal cVar1S15S42P018P048P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S42P018P048P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S42P018P048P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S42P018P048P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S42P018P048P011P013: std_logic_vector(   0 downto 0);
        signal cVar1S20S42P018N048P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S42P018N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S22S42P018N048P044N023: std_logic_vector(   0 downto 0);
        signal cVar1S23S42P018N048N044P004: std_logic_vector(   0 downto 0);
        signal cVar1S24S42P018N048N044P004: std_logic_vector(   0 downto 0);
        signal cVar1S25S42P018N048N044P004: std_logic_vector(   0 downto 0);
        signal cVar1S26S42P018N048N044P004: std_logic_vector(   0 downto 0);
        signal cVar1S27S42P018N048N044P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S43P048P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S43P048P025N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S43P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S43P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S43P048P025N007N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S43P048N025P062P058nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S43P048N025P062N058: std_logic_vector(   0 downto 0);
        signal cVar1S7S43P048N025N062P027: std_logic_vector(   0 downto 0);
        signal cVar1S8S43P048N025N062P027: std_logic_vector(   0 downto 0);
        signal cVar1S9S43P048N025N062P027: std_logic_vector(   0 downto 0);
        signal cVar1S10S43P048N025N062N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S43P048N025N062N027: std_logic_vector(   0 downto 0);
        signal cVar1S12S43N048P022P043P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S43N048P022N043P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S43N048P022N043N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S43N048N022P038P021: std_logic_vector(   0 downto 0);
        signal cVar1S16S43N048N022P038P021: std_logic_vector(   0 downto 0);
        signal cVar1S17S43N048N022P038N021: std_logic_vector(   0 downto 0);
        signal cVar1S18S43N048N022P038N021: std_logic_vector(   0 downto 0);
        signal cVar1S19S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S20S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S21S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S22S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S23S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S24S43N048N022N038P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S44P022P043P037P010nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S44P022P043P037P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S44P022N043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S44P022N043N004P047: std_logic_vector(   0 downto 0);
        signal cVar1S4S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S5S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S6S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S7S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S8S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S44N022P004P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S11S44N022P004P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S12S44N022P004P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S13S44N022P004P043N023: std_logic_vector(   0 downto 0);
        signal cVar1S14S44N022P004P043N023: std_logic_vector(   0 downto 0);
        signal cVar1S15S44N022P004P043N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S44N022P004P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S44N022P004N040P017: std_logic_vector(   0 downto 0);
        signal cVar1S18S44N022P004N040P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S44N022P004N040N017: std_logic_vector(   0 downto 0);
        signal cVar1S20S44N022P004N040N017: std_logic_vector(   0 downto 0);
        signal cVar1S21S44N022P004N040N017: std_logic_vector(   0 downto 0);
        signal cVar1S0S45P022P043P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S45P022P043N019P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S45P022N043P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S45P022N043N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S45P022N043N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S45P022N043N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S45P022N043N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S45N022P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S45N022P047N006P008: std_logic_vector(   0 downto 0);
        signal cVar1S9S45N022P047N006P008: std_logic_vector(   0 downto 0);
        signal cVar1S10S45N022P047N006P008: std_logic_vector(   0 downto 0);
        signal cVar1S11S45N022P047N006N008: std_logic_vector(   0 downto 0);
        signal cVar1S12S45N022P047N006N008: std_logic_vector(   0 downto 0);
        signal cVar1S13S45N022P047N006N008: std_logic_vector(   0 downto 0);
        signal cVar1S14S45N022N047P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S45N022N047P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S45N022N047P051P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S45N022N047P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S18S45N022N047P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S19S45N022N047P051N008: std_logic_vector(   0 downto 0);
        signal cVar1S20S45N022N047N051P049: std_logic_vector(   0 downto 0);
        signal cVar1S21S45N022N047N051P049: std_logic_vector(   0 downto 0);
        signal cVar1S22S45N022N047N051P049: std_logic_vector(   0 downto 0);
        signal cVar1S23S45N022N047N051P049: std_logic_vector(   0 downto 0);
        signal cVar1S24S45N022N047N051P049: std_logic_vector(   0 downto 0);
        signal cVar1S0S46P022P043P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S46P022P043N019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S46P022N043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S46P022N043N004P047: std_logic_vector(   0 downto 0);
        signal cVar1S4S46P022N043N004P047: std_logic_vector(   0 downto 0);
        signal cVar1S5S46N022P048P025P050: std_logic_vector(   0 downto 0);
        signal cVar1S6S46N022P048N025P043: std_logic_vector(   0 downto 0);
        signal cVar1S7S46N022P048N025P043: std_logic_vector(   0 downto 0);
        signal cVar1S8S46N022P048N025P043: std_logic_vector(   0 downto 0);
        signal cVar1S9S46N022N048P037P065: std_logic_vector(   0 downto 0);
        signal cVar1S10S46N022N048P037P065: std_logic_vector(   0 downto 0);
        signal cVar1S11S46N022N048P037P065: std_logic_vector(   0 downto 0);
        signal cVar1S12S46N022N048P037P065: std_logic_vector(   0 downto 0);
        signal cVar1S13S46N022N048P037P065: std_logic_vector(   0 downto 0);
        signal cVar1S14S46N022N048N037P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S46N022N048N037P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S46N022N048N037P023: std_logic_vector(   0 downto 0);
        signal cVar1S17S46N022N048N037N023: std_logic_vector(   0 downto 0);
        signal cVar1S18S46N022N048N037N023: std_logic_vector(   0 downto 0);
        signal cVar1S19S46N022N048N037N023: std_logic_vector(   0 downto 0);
        signal cVar1S20S46N022N048N037N023: std_logic_vector(   0 downto 0);
        signal cVar1S0S47P022P043P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S47P022P043N019P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S47P022P043N019P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S47P022P043N019P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S47P022N043P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S47P022N043N004P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S47P022N043N004P047: std_logic_vector(   0 downto 0);
        signal cVar1S7S47N022P023P005P068: std_logic_vector(   0 downto 0);
        signal cVar1S8S47N022P023P005P068: std_logic_vector(   0 downto 0);
        signal cVar1S9S47N022P023N005P034: std_logic_vector(   0 downto 0);
        signal cVar1S10S47N022P023N005P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S47N022P023N005P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S47N022N023P043P048: std_logic_vector(   0 downto 0);
        signal cVar1S13S47N022N023P043P048: std_logic_vector(   0 downto 0);
        signal cVar1S14S47N022N023P043P048: std_logic_vector(   0 downto 0);
        signal cVar1S15S47N022N023P043N048: std_logic_vector(   0 downto 0);
        signal cVar1S16S47N022N023P043N048: std_logic_vector(   0 downto 0);
        signal cVar1S17S47N022N023P043N048: std_logic_vector(   0 downto 0);
        signal cVar1S18S47N022N023P043N048: std_logic_vector(   0 downto 0);
        signal cVar1S19S47N022N023P043P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S47N022N023P043N006: std_logic_vector(   0 downto 0);
        signal cVar1S21S47N022N023P043N006: std_logic_vector(   0 downto 0);
        signal cVar1S22S47N022N023P043N006: std_logic_vector(   0 downto 0);
        signal cVar1S23S47N022N023P043N006: std_logic_vector(   0 downto 0);
        signal cVar1S0S48P016P065P034P059: std_logic_vector(   0 downto 0);
        signal cVar1S1S48P016P065P034P059: std_logic_vector(   0 downto 0);
        signal cVar1S2S48P016P065P034N059: std_logic_vector(   0 downto 0);
        signal cVar1S3S48P016P065P034N059: std_logic_vector(   0 downto 0);
        signal cVar1S4S48P016P065P034N059: std_logic_vector(   0 downto 0);
        signal cVar1S5S48P016P065P034N059: std_logic_vector(   0 downto 0);
        signal cVar1S6S48P016P065P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S48P016P065P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S48P016P065P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S9S48P016P065P034N014: std_logic_vector(   0 downto 0);
        signal cVar1S10S48P016P065P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S48P016P065P067P063: std_logic_vector(   0 downto 0);
        signal cVar1S12S48P016P065P067P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S48P016P065N067P066: std_logic_vector(   0 downto 0);
        signal cVar1S14S48P016P065N067P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S48P016P065N067P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S48P016P065N067P066: std_logic_vector(   0 downto 0);
        signal cVar1S17S48P016P065N067P066: std_logic_vector(   0 downto 0);
        signal cVar1S18S48P016P063P015P057: std_logic_vector(   0 downto 0);
        signal cVar1S19S48P016P063P015P057: std_logic_vector(   0 downto 0);
        signal cVar1S20S48P016P063P015P057: std_logic_vector(   0 downto 0);
        signal cVar1S21S48P016P063P015P056: std_logic_vector(   0 downto 0);
        signal cVar1S22S48P016P063P015P056: std_logic_vector(   0 downto 0);
        signal cVar1S23S48P016P063P015P056: std_logic_vector(   0 downto 0);
        signal cVar1S24S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S25S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S26S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S27S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S28S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S29S48P016N063P052P061: std_logic_vector(   0 downto 0);
        signal cVar1S30S48P016N063P052P060: std_logic_vector(   0 downto 0);
        signal cVar1S31S48P016N063P052P060: std_logic_vector(   0 downto 0);
        signal cVar1S0S49P023P005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S49P023P005N042P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S49P023N005P034P007: std_logic_vector(   0 downto 0);
        signal cVar1S3S49P023N005P034P007: std_logic_vector(   0 downto 0);
        signal cVar1S4S49P023N005P034N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S49P023N005P034N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S49P023N005P034N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S49N023P022P043P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S49N023P022P043N005: std_logic_vector(   0 downto 0);
        signal cVar1S9S49N023P022P043N005: std_logic_vector(   0 downto 0);
        signal cVar1S10S49N023P022P043N005: std_logic_vector(   0 downto 0);
        signal cVar1S11S49N023P022N043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S49N023P022N043N004: std_logic_vector(   0 downto 0);
        signal cVar1S13S49N023P022N043N004: std_logic_vector(   0 downto 0);
        signal cVar1S14S49N023P022N043N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S49N023N022P016P035: std_logic_vector(   0 downto 0);
        signal cVar1S16S49N023N022P016P035: std_logic_vector(   0 downto 0);
        signal cVar1S17S49N023N022P016P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S49N023N022P016P035: std_logic_vector(   0 downto 0);
        signal cVar1S19S49N023N022N016P028: std_logic_vector(   0 downto 0);
        signal cVar1S20S49N023N022N016P028: std_logic_vector(   0 downto 0);
        signal cVar1S21S49N023N022N016P028: std_logic_vector(   0 downto 0);
        signal cVar1S22S49N023N022N016N028: std_logic_vector(   0 downto 0);
        signal cVar1S23S49N023N022N016N028: std_logic_vector(   0 downto 0);
        signal cVar1S24S49N023N022N016N028: std_logic_vector(   0 downto 0);
        signal cVar1S0S50P023P005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S50P023P005N042P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S50P023N005P034P007: std_logic_vector(   0 downto 0);
        signal cVar1S3S50P023N005P034P007: std_logic_vector(   0 downto 0);
        signal cVar1S4S50P023N005P034N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S50P023N005P034N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S50N023P028P029P010: std_logic_vector(   0 downto 0);
        signal cVar1S7S50N023P028P029N010: std_logic_vector(   0 downto 0);
        signal cVar1S8S50N023P028P029N010: std_logic_vector(   0 downto 0);
        signal cVar1S9S50N023N028P053P025: std_logic_vector(   0 downto 0);
        signal cVar1S10S50N023N028P053P025: std_logic_vector(   0 downto 0);
        signal cVar1S11S50N023N028P053N025: std_logic_vector(   0 downto 0);
        signal cVar1S12S50N023N028P053N025: std_logic_vector(   0 downto 0);
        signal cVar1S13S50N023N028P053N025: std_logic_vector(   0 downto 0);
        signal cVar1S14S50N023N028P053N025: std_logic_vector(   0 downto 0);
        signal cVar1S15S50N023N028P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S16S50N023N028P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S17S50N023N028P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S18S50N023N028P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S19S50N023N028P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S0S51P028P029P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S1S51P028P029P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S2S51P028P029P010P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S51P028P029N010P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S51P028P029N010N008: std_logic_vector(   0 downto 0);
        signal cVar1S5S51N028P023P005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S51N028P023P005N042: std_logic_vector(   0 downto 0);
        signal cVar1S7S51N028P023N005P049: std_logic_vector(   0 downto 0);
        signal cVar1S8S51N028P023N005P049: std_logic_vector(   0 downto 0);
        signal cVar1S9S51N028N023P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S51N028N023P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S11S51N028N023P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S12S51N028N023N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S51N028N023N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S51N028N023N025P024: std_logic_vector(   0 downto 0);
        signal cVar1S15S51N028N023N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S16S51N028N023N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S17S51N028N023N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S0S52P045P043P005P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S52P045P043N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S52P045P043N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S52P045P043N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S52P045P043N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S52P045N043P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S52P045N043P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S7S52P045N043P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S8S52P045N043N047P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S52P045N043N047N048: std_logic_vector(   0 downto 0);
        signal cVar1S10S52P045N043N047N048: std_logic_vector(   0 downto 0);
        signal cVar1S11S52P045N043N047N048: std_logic_vector(   0 downto 0);
        signal cVar1S12S52N045P028P010P055: std_logic_vector(   0 downto 0);
        signal cVar1S13S52N045P028P010N055: std_logic_vector(   0 downto 0);
        signal cVar1S14S52N045P028P010N055: std_logic_vector(   0 downto 0);
        signal cVar1S15S52N045P028N010P011: std_logic_vector(   0 downto 0);
        signal cVar1S16S52N045P028N010P011: std_logic_vector(   0 downto 0);
        signal cVar1S17S52N045P028N010P011: std_logic_vector(   0 downto 0);
        signal cVar1S18S52N045P028N010N011: std_logic_vector(   0 downto 0);
        signal cVar1S19S52N045P028N010N011: std_logic_vector(   0 downto 0);
        signal cVar1S20S52N045N028P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S21S52N045N028P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S22S52N045N028P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S23S52N045N028P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S24S52N045N028N040P025: std_logic_vector(   0 downto 0);
        signal cVar1S25S52N045N028N040P025: std_logic_vector(   0 downto 0);
        signal cVar1S26S52N045N028N040P025: std_logic_vector(   0 downto 0);
        signal cVar1S27S52N045N028N040N025: std_logic_vector(   0 downto 0);
        signal cVar1S28S52N045N028N040N025: std_logic_vector(   0 downto 0);
        signal cVar1S29S52N045N028N040N025: std_logic_vector(   0 downto 0);
        signal cVar1S30S52N045N028N040N025: std_logic_vector(   0 downto 0);
        signal cVar1S0S53P025P007P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S53P025P007P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S53P025N007P046P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S53P025N007P046N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S53P025N007P046N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S53P025N007N046P003: std_logic_vector(   0 downto 0);
        signal cVar1S6S53P025N007N046P003: std_logic_vector(   0 downto 0);
        signal cVar1S7S53N025P028P010P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S53N025P028P010N055: std_logic_vector(   0 downto 0);
        signal cVar1S9S53N025P028P010N055: std_logic_vector(   0 downto 0);
        signal cVar1S10S53N025P028N010P029: std_logic_vector(   0 downto 0);
        signal cVar1S11S53N025P028N010P029: std_logic_vector(   0 downto 0);
        signal cVar1S12S53N025P028N010P029: std_logic_vector(   0 downto 0);
        signal cVar1S13S53N025N028P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S14S53N025N028P040P021: std_logic_vector(   0 downto 0);
        signal cVar1S15S53N025N028P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S16S53N025N028P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S17S53N025N028N040P045: std_logic_vector(   0 downto 0);
        signal cVar1S18S53N025N028N040P045: std_logic_vector(   0 downto 0);
        signal cVar1S19S53N025N028N040P045: std_logic_vector(   0 downto 0);
        signal cVar1S20S53N025N028N040N045: std_logic_vector(   0 downto 0);
        signal cVar1S21S53N025N028N040N045: std_logic_vector(   0 downto 0);
        signal cVar1S22S53N025N028N040N045: std_logic_vector(   0 downto 0);
        signal cVar1S23S53N025N028N040N045: std_logic_vector(   0 downto 0);
        signal cVar1S0S54P018P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S54P018P040N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S54P018P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S54P018P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S54P018P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S54P018N040P045P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S54P018N040P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S54P018N040P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S8S54P018N040P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S9S54P018N040N045P015: std_logic_vector(   0 downto 0);
        signal cVar1S10S54P018N040N045P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S54P018N040N045N015: std_logic_vector(   0 downto 0);
        signal cVar1S12S54P018N040N045N015: std_logic_vector(   0 downto 0);
        signal cVar1S13S54P018N040N045N015: std_logic_vector(   0 downto 0);
        signal cVar1S14S54P018P015P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S15S54P018P015P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S16S54P018P015P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S54P018P015P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S54P018P015N019P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S54P018N015P019P007: std_logic_vector(   0 downto 0);
        signal cVar1S20S54P018N015P019P007: std_logic_vector(   0 downto 0);
        signal cVar1S21S54P018N015P019P007: std_logic_vector(   0 downto 0);
        signal cVar1S22S54P018N015P019P007: std_logic_vector(   0 downto 0);
        signal cVar1S23S54P018N015P019P059: std_logic_vector(   0 downto 0);
        signal cVar1S24S54P018N015P019P059: std_logic_vector(   0 downto 0);
        signal cVar1S25S54P018N015P019N059: std_logic_vector(   0 downto 0);
        signal cVar1S26S54P018N015P019N059: std_logic_vector(   0 downto 0);
        signal cVar1S0S55P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S55P040N002P015P021: std_logic_vector(   0 downto 0);
        signal cVar1S2S55P040N002P015P021: std_logic_vector(   0 downto 0);
        signal cVar1S3S55P040N002P015N021: std_logic_vector(   0 downto 0);
        signal cVar1S4S55P040N002P015N021: std_logic_vector(   0 downto 0);
        signal cVar1S5S55P040N002P015N021: std_logic_vector(   0 downto 0);
        signal cVar1S6S55P040N002P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S55P040N002P015N013: std_logic_vector(   0 downto 0);
        signal cVar1S8S55N040P045P005P068: std_logic_vector(   0 downto 0);
        signal cVar1S9S55N040P045N005P004: std_logic_vector(   0 downto 0);
        signal cVar1S10S55N040P045N005P004: std_logic_vector(   0 downto 0);
        signal cVar1S11S55N040P045N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S12S55N040P045N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S13S55N040P045N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S14S55N040P045N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S55N040N045P015P047: std_logic_vector(   0 downto 0);
        signal cVar1S16S55N040N045P015P047: std_logic_vector(   0 downto 0);
        signal cVar1S17S55N040N045P015P047: std_logic_vector(   0 downto 0);
        signal cVar1S18S55N040N045P015P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S55N040N045P015P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S55N040N045N015P028: std_logic_vector(   0 downto 0);
        signal cVar1S21S55N040N045N015P028: std_logic_vector(   0 downto 0);
        signal cVar1S22S55N040N045N015N028: std_logic_vector(   0 downto 0);
        signal cVar1S23S55N040N045N015N028: std_logic_vector(   0 downto 0);
        signal cVar1S24S55N040N045N015N028: std_logic_vector(   0 downto 0);
        signal cVar1S25S55N040N045N015N028: std_logic_vector(   0 downto 0);
        signal cVar1S0S56P045P005P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S56P045N005P004P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S56P045N005N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S56P045N005N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S56P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S56P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S6S56P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S7S56N045P040P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S56N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S56N045P040N021P066: std_logic_vector(   0 downto 0);
        signal cVar1S10S56N045P040N021P066: std_logic_vector(   0 downto 0);
        signal cVar1S11S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S12S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S13S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S16S56N045N040P018P043: std_logic_vector(   0 downto 0);
        signal cVar1S17S56N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S18S56N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S19S56N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S20S56N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S21S56N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S0S57P045P005P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S57P045N005P004P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S57P045N005N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S57P045N005N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S57P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S57P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S6S57P045N005N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S7S57N045P040P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S57N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S57N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S10S57N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S11S57N045P040N021P020: std_logic_vector(   0 downto 0);
        signal cVar1S12S57N045P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S13S57N045P040N021N020: std_logic_vector(   0 downto 0);
        signal cVar1S14S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S15S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S16S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S17S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S18S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S19S57N045N040P018P060: std_logic_vector(   0 downto 0);
        signal cVar1S20S57N045N040N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S21S57N045N040N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S22S57N045N040N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S23S57N045N040N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S24S57N045N040N018P043: std_logic_vector(   0 downto 0);
        signal cVar1S0S58P045P005P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S58P045N005P021P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S58P045N005P021N006: std_logic_vector(   0 downto 0);
        signal cVar1S3S58P045N005P021N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S58P045N005P021N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S58N045P018P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S58N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S7S58N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S8S58N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S10S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S11S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S12S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S13S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S16S58N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S17S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S19S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S20S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S21S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S22S58N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S23S58N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S24S58N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S25S58N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S26S58N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S0S59P045P022P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S59P045P022N019P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S59P045N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S59P045N022N023P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S59P045N022N023N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S59P045N022N023N006: std_logic_vector(   0 downto 0);
        signal cVar1S6S59P045N022N023N006: std_logic_vector(   0 downto 0);
        signal cVar1S7S59N045P040P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S59N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S59N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S10S59N045P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S11S59N045P040N021P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S59N045P040N021P066: std_logic_vector(   0 downto 0);
        signal cVar1S13S59N045N040P025P007: std_logic_vector(   0 downto 0);
        signal cVar1S14S59N045N040P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S15S59N045N040P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S16S59N045N040P025N007: std_logic_vector(   0 downto 0);
        signal cVar1S17S59N045N040N025P018: std_logic_vector(   0 downto 0);
        signal cVar1S18S59N045N040N025P018: std_logic_vector(   0 downto 0);
        signal cVar1S19S59N045N040N025N018: std_logic_vector(   0 downto 0);
        signal cVar1S20S59N045N040N025N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S59N045N040N025N018: std_logic_vector(   0 downto 0);
        signal cVar1S0S60P045P005P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S60P045N005P021P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S60P045N005P021P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S60P045N005P021P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S60P045N005P021N024psss: std_logic_vector(   0 downto 0);
        signal cVar1S5S60N045P018P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S60N045P018P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S60N045P018P040P002: std_logic_vector(   0 downto 0);
        signal cVar1S8S60N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S60N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S10S60N045P018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S11S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S12S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S13S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S16S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S17S60N045P018N040P043: std_logic_vector(   0 downto 0);
        signal cVar1S18S60N045P018P025P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S60N045P018P025N035: std_logic_vector(   0 downto 0);
        signal cVar1S20S60N045P018P025N035: std_logic_vector(   0 downto 0);
        signal cVar1S21S60N045P018N025P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S60N045P018N025P037: std_logic_vector(   0 downto 0);
        signal cVar1S23S60N045P018N025P037: std_logic_vector(   0 downto 0);
        signal cVar1S24S60N045P018N025P037: std_logic_vector(   0 downto 0);
        signal cVar1S25S60N045P018N025P037: std_logic_vector(   0 downto 0);
        signal cVar1S0S61P045P005P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S61P045N005P021P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S61P045N005P021P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S61P045N005P021N024: std_logic_vector(   0 downto 0);
        signal cVar1S4S61P045N005P021N024: std_logic_vector(   0 downto 0);
        signal cVar1S5S61P045N005P021N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S61N045P018P037P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S61N045P018P037P061: std_logic_vector(   0 downto 0);
        signal cVar1S8S61N045P018P037P061: std_logic_vector(   0 downto 0);
        signal cVar1S9S61N045P018P037N061: std_logic_vector(   0 downto 0);
        signal cVar1S10S61N045P018P037N061: std_logic_vector(   0 downto 0);
        signal cVar1S11S61N045P018P037N061: std_logic_vector(   0 downto 0);
        signal cVar1S12S61N045P018P037P066: std_logic_vector(   0 downto 0);
        signal cVar1S13S61N045P018P037P066: std_logic_vector(   0 downto 0);
        signal cVar1S14S61N045P018P037P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S61N045P018P037P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S61N045N018P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S61N045N018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S18S61N045N018P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S19S61N045N018N040P000: std_logic_vector(   0 downto 0);
        signal cVar1S20S61N045N018N040P000: std_logic_vector(   0 downto 0);
        signal cVar1S21S61N045N018N040P000: std_logic_vector(   0 downto 0);
        signal cVar1S22S61N045N018N040P000: std_logic_vector(   0 downto 0);
        signal cVar1S0S62P045P005P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S62P045N005P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S62P045N005P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S62P045N005P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S62P045N005P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S5S62P045N005P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S62P045N005P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S7S62P045N005P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S8S62N045P018P000P030: std_logic_vector(   0 downto 0);
        signal cVar1S9S62N045P018P000P030: std_logic_vector(   0 downto 0);
        signal cVar1S10S62N045P018P000N030: std_logic_vector(   0 downto 0);
        signal cVar1S11S62N045P018P000N030: std_logic_vector(   0 downto 0);
        signal cVar1S12S62N045P018P000N030: std_logic_vector(   0 downto 0);
        signal cVar1S13S62N045P018P000N030: std_logic_vector(   0 downto 0);
        signal cVar1S14S62N045P018P000P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S62N045P018P000N040: std_logic_vector(   0 downto 0);
        signal cVar1S16S62N045P018P000N040: std_logic_vector(   0 downto 0);
        signal cVar1S17S62N045P018P061P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S62N045P018P061N035: std_logic_vector(   0 downto 0);
        signal cVar1S19S62N045P018P061N035: std_logic_vector(   0 downto 0);
        signal cVar1S20S62N045P018P061N035: std_logic_vector(   0 downto 0);
        signal cVar1S21S62N045P018N061P025: std_logic_vector(   0 downto 0);
        signal cVar1S22S62N045P018N061P025: std_logic_vector(   0 downto 0);
        signal cVar1S23S62N045P018N061N025: std_logic_vector(   0 downto 0);
        signal cVar1S24S62N045P018N061N025: std_logic_vector(   0 downto 0);
        signal cVar1S0S63P045P005P037nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S63P045N005P021P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S63P045N005P021N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S63P045N005P021N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S63P045N005P021N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S6S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S11S63N045P018P019P056: std_logic_vector(   0 downto 0);
        signal cVar1S12S63N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S63N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S63N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S15S63N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S16S63N045P018N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S17S63N045N018P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S18S63N045N018P030P031: std_logic_vector(   0 downto 0);
        signal cVar1S19S63N045N018N030P031: std_logic_vector(   0 downto 0);
        signal cVar1S20S63N045N018N030P031: std_logic_vector(   0 downto 0);
        signal cVar1S21S63N045N018N030P031: std_logic_vector(   0 downto 0);
        signal cVar1S22S63N045N018N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S23S63N045N018N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S24S63N045N018N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S25S63N045N018N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S64P018P069P011P029: std_logic_vector(   0 downto 0);
        signal cVar1S1S64P018P069P011P029: std_logic_vector(   0 downto 0);
        signal cVar1S2S64P018P069P011P029: std_logic_vector(   0 downto 0);
        signal cVar1S3S64P018P069P011N029: std_logic_vector(   0 downto 0);
        signal cVar1S4S64P018P069P011N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S64P018P069P011N029: std_logic_vector(   0 downto 0);
        signal cVar1S6S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S7S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S8S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S9S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S10S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S11S64P018P069N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S12S64P018P069P019P067: std_logic_vector(   0 downto 0);
        signal cVar1S13S64P018P069P019P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S64P018P069P019P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S64P018P069P019N067: std_logic_vector(   0 downto 0);
        signal cVar1S16S64P018P069N019P068: std_logic_vector(   0 downto 0);
        signal cVar1S17S64P018P069N019P068: std_logic_vector(   0 downto 0);
        signal cVar1S18S64P018P069N019N068: std_logic_vector(   0 downto 0);
        signal cVar1S19S64P018P069N019N068: std_logic_vector(   0 downto 0);
        signal cVar1S20S64P018P031P007P013: std_logic_vector(   0 downto 0);
        signal cVar1S21S64P018P031P007P013: std_logic_vector(   0 downto 0);
        signal cVar1S22S64P018P031P007P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S64P018P031P007N013: std_logic_vector(   0 downto 0);
        signal cVar1S24S64P018P031P007N013: std_logic_vector(   0 downto 0);
        signal cVar1S25S64P018N031P007P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S64P018N031P007N051: std_logic_vector(   0 downto 0);
        signal cVar1S27S64P018N031P007N051: std_logic_vector(   0 downto 0);
        signal cVar1S28S64P018N031P007N051: std_logic_vector(   0 downto 0);
        signal cVar1S29S64P018N031N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S30S64P018N031N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S31S64P018N031N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S32S64P018N031N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S33S64P018N031N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S34S64P018N031N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S0S65P018P014P042P068: std_logic_vector(   0 downto 0);
        signal cVar1S1S65P018P014P042P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S65P018P014P042N068: std_logic_vector(   0 downto 0);
        signal cVar1S3S65P018P014P042N068: std_logic_vector(   0 downto 0);
        signal cVar1S4S65P018P014P042P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S65P018P014P042N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S65P018P014P042N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S65P018P014P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S65P018P014N045P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S65P018P014N045N046: std_logic_vector(   0 downto 0);
        signal cVar1S10S65P018P014N045N046: std_logic_vector(   0 downto 0);
        signal cVar1S11S65P018P014N045N046: std_logic_vector(   0 downto 0);
        signal cVar1S12S65P018P014N045N046: std_logic_vector(   0 downto 0);
        signal cVar1S13S65N018P041P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S65N018P041P020N002: std_logic_vector(   0 downto 0);
        signal cVar1S15S65N018P041P020N002: std_logic_vector(   0 downto 0);
        signal cVar1S16S65N018P041N020P023: std_logic_vector(   0 downto 0);
        signal cVar1S17S65N018P041N020N023: std_logic_vector(   0 downto 0);
        signal cVar1S18S65N018P041N020N023: std_logic_vector(   0 downto 0);
        signal cVar1S19S65N018N041P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S20S65N018N041P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S21S65N018N041P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S22S65N018N041P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S23S65N018N041P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S24S65N018N041P039P049nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S65N018N041P039N049: std_logic_vector(   0 downto 0);
        signal cVar1S0S66P018P041P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S66P018P041P020N002: std_logic_vector(   0 downto 0);
        signal cVar1S2S66P018P041P020N002: std_logic_vector(   0 downto 0);
        signal cVar1S3S66P018P041N020P023: std_logic_vector(   0 downto 0);
        signal cVar1S4S66P018P041N020N023: std_logic_vector(   0 downto 0);
        signal cVar1S5S66P018P041N020N023: std_logic_vector(   0 downto 0);
        signal cVar1S6S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S7S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S8S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S9S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S10S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S11S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S12S66P018N041P039P020: std_logic_vector(   0 downto 0);
        signal cVar1S13S66P018N041P039P011: std_logic_vector(   0 downto 0);
        signal cVar1S14S66P018P068P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S66P018P068N057P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S66P018P068N057P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S66P018P068N057P063: std_logic_vector(   0 downto 0);
        signal cVar1S18S66P018P068N057P063: std_logic_vector(   0 downto 0);
        signal cVar1S19S66P018P068N057P063: std_logic_vector(   0 downto 0);
        signal cVar1S20S66P018N068P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S21S66P018N068P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S22S66P018N068P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S23S66P018N068N031P005: std_logic_vector(   0 downto 0);
        signal cVar1S24S66P018N068N031N005: std_logic_vector(   0 downto 0);
        signal cVar1S25S66P018N068N031N005: std_logic_vector(   0 downto 0);
        signal cVar1S26S66P018N068N031N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S67P009P027P063P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S67P009P027P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S67P009P027P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S3S67P009N027P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S67P009N027P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S5S67P009N027P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S6S67P009N027N049P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S67P009N027N049P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S67P009N027N049N014: std_logic_vector(   0 downto 0);
        signal cVar1S9S67P009N027N049N014: std_logic_vector(   0 downto 0);
        signal cVar1S10S67P009N027N049N014: std_logic_vector(   0 downto 0);
        signal cVar1S11S67N009P041P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S67N009P041N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S67N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S14S67N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S15S67N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S16S67N009N041P018P000: std_logic_vector(   0 downto 0);
        signal cVar1S17S67N009N041P018P000: std_logic_vector(   0 downto 0);
        signal cVar1S18S67N009N041P018N000: std_logic_vector(   0 downto 0);
        signal cVar1S19S67N009N041P018N000: std_logic_vector(   0 downto 0);
        signal cVar1S20S67N009N041P018N000: std_logic_vector(   0 downto 0);
        signal cVar1S21S67N009N041P018N000: std_logic_vector(   0 downto 0);
        signal cVar1S22S67N009N041N018P039: std_logic_vector(   0 downto 0);
        signal cVar1S23S67N009N041N018P039: std_logic_vector(   0 downto 0);
        signal cVar1S24S67N009N041N018P039: std_logic_vector(   0 downto 0);
        signal cVar1S25S67N009N041N018P039: std_logic_vector(   0 downto 0);
        signal cVar1S26S67N009N041N018P039: std_logic_vector(   0 downto 0);
        signal cVar1S0S68P009P027P063P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S68P009P027P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S68P009N027P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S68P009N027P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S4S68P009N027P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S5S68P009N027N049P053: std_logic_vector(   0 downto 0);
        signal cVar1S6S68P009N027N049P053: std_logic_vector(   0 downto 0);
        signal cVar1S7S68P009N027N049N053: std_logic_vector(   0 downto 0);
        signal cVar1S8S68P009N027N049N053: std_logic_vector(   0 downto 0);
        signal cVar1S9S68P009N027N049N053: std_logic_vector(   0 downto 0);
        signal cVar1S10S68P009N027N049N053: std_logic_vector(   0 downto 0);
        signal cVar1S11S68N009P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S68N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S13S68N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S14S68N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S15S68N009P041N020P021: std_logic_vector(   0 downto 0);
        signal cVar1S16S68N009P041N020P021: std_logic_vector(   0 downto 0);
        signal cVar1S17S68N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S18S68N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S19S68N009P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S20S68N009N041P016P031: std_logic_vector(   0 downto 0);
        signal cVar1S21S68N009N041P016P031: std_logic_vector(   0 downto 0);
        signal cVar1S22S68N009N041P016P031: std_logic_vector(   0 downto 0);
        signal cVar1S23S68N009N041P016P031: std_logic_vector(   0 downto 0);
        signal cVar1S24S68N009N041P016N031: std_logic_vector(   0 downto 0);
        signal cVar1S25S68N009N041P016N031: std_logic_vector(   0 downto 0);
        signal cVar1S26S68N009N041P016N031: std_logic_vector(   0 downto 0);
        signal cVar1S27S68N009N041P016P059: std_logic_vector(   0 downto 0);
        signal cVar1S28S68N009N041P016P059: std_logic_vector(   0 downto 0);
        signal cVar1S29S68N009N041P016P059: std_logic_vector(   0 downto 0);
        signal cVar1S30S68N009N041P016P059: std_logic_vector(   0 downto 0);
        signal cVar1S31S68N009N041P016P059: std_logic_vector(   0 downto 0);
        signal cVar1S0S69P009P049P060P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S69P009P049P060P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S69P009P049P060P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S69P009N049P053P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S69P009N049P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S69P009N049P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S6S69P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S69P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S8S69P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S9S69P009N049N053N050: std_logic_vector(   0 downto 0);
        signal cVar1S10S69P009N049N053N050: std_logic_vector(   0 downto 0);
        signal cVar1S11S69N009P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S69N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S13S69N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S14S69N009P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S15S69N009P041N020P001nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S69N009P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S17S69N009P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S18S69N009P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S19S69N009N041P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S20S69N009N041P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S21S69N009N041P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S22S69N009N041P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S69N009N041P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S24S69N009N041P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S25S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S26S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S27S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S28S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S29S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S30S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S31S69N009N041N031P054: std_logic_vector(   0 downto 0);
        signal cVar1S0S70P016P018P036P053: std_logic_vector(   0 downto 0);
        signal cVar1S1S70P016P018P036P053: std_logic_vector(   0 downto 0);
        signal cVar1S2S70P016P018P036P053: std_logic_vector(   0 downto 0);
        signal cVar1S3S70P016P018P036N053: std_logic_vector(   0 downto 0);
        signal cVar1S4S70P016P018P036N053: std_logic_vector(   0 downto 0);
        signal cVar1S5S70P016P018P036N053: std_logic_vector(   0 downto 0);
        signal cVar1S6S70P016P018P036N053: std_logic_vector(   0 downto 0);
        signal cVar1S7S70P016P018P036P017: std_logic_vector(   0 downto 0);
        signal cVar1S8S70P016P018P036P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S70P016P018P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S10S70P016P018P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S11S70P016P018P036N017: std_logic_vector(   0 downto 0);
        signal cVar1S12S70P016P018P045P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S70P016P018N045P026: std_logic_vector(   0 downto 0);
        signal cVar1S14S70P016P018N045P026: std_logic_vector(   0 downto 0);
        signal cVar1S15S70P016P018N045P026: std_logic_vector(   0 downto 0);
        signal cVar1S16S70P016P018N045P026: std_logic_vector(   0 downto 0);
        signal cVar1S17S70P016P018N045P026: std_logic_vector(   0 downto 0);
        signal cVar1S18S70P016P035P053P041: std_logic_vector(   0 downto 0);
        signal cVar1S19S70P016P035P053P041: std_logic_vector(   0 downto 0);
        signal cVar1S20S70P016P035P053N041: std_logic_vector(   0 downto 0);
        signal cVar1S21S70P016P035P053N041: std_logic_vector(   0 downto 0);
        signal cVar1S22S70P016P035P053N041: std_logic_vector(   0 downto 0);
        signal cVar1S23S70P016P035P053P037: std_logic_vector(   0 downto 0);
        signal cVar1S24S70P016P035P053N037: std_logic_vector(   0 downto 0);
        signal cVar1S25S70P016P035P053N037: std_logic_vector(   0 downto 0);
        signal cVar1S26S70P016P035P032P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S27S70P016P035N032P034: std_logic_vector(   0 downto 0);
        signal cVar1S0S71P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S71P041P020N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S71P041P020N003N002: std_logic_vector(   0 downto 0);
        signal cVar1S3S71P041P020N003N002: std_logic_vector(   0 downto 0);
        signal cVar1S4S71P041N020P001nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S71P041N020N001P005: std_logic_vector(   0 downto 0);
        signal cVar1S6S71P041N020N001P005: std_logic_vector(   0 downto 0);
        signal cVar1S7S71P041N020N001P005: std_logic_vector(   0 downto 0);
        signal cVar1S8S71P041N020N001N005: std_logic_vector(   0 downto 0);
        signal cVar1S9S71P041N020N001N005: std_logic_vector(   0 downto 0);
        signal cVar1S10S71P041N020N001N005: std_logic_vector(   0 downto 0);
        signal cVar1S11S71N041P049P026P033: std_logic_vector(   0 downto 0);
        signal cVar1S12S71N041P049N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S71N041P049N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S71N041P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S15S71N041P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S16S71N041P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S17S71N041N049P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S18S71N041N049P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S19S71N041N049P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S20S71N041N049P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S21S71N041N049P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S22S71N041N049P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S23S71N041N049P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S24S71N041N049P039P036nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S71N041N049P039N036: std_logic_vector(   0 downto 0);
        signal cVar1S26S71N041N049P039N036: std_logic_vector(   0 downto 0);
        signal cVar1S0S72P016P018P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S72P016P018P023N042: std_logic_vector(   0 downto 0);
        signal cVar1S2S72P016P018P023N042: std_logic_vector(   0 downto 0);
        signal cVar1S3S72P016P018N023P047: std_logic_vector(   0 downto 0);
        signal cVar1S4S72P016P018N023P047: std_logic_vector(   0 downto 0);
        signal cVar1S5S72P016P018N023P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S72P016P018N023N047: std_logic_vector(   0 downto 0);
        signal cVar1S7S72P016P018N023N047: std_logic_vector(   0 downto 0);
        signal cVar1S8S72P016P018N023N047: std_logic_vector(   0 downto 0);
        signal cVar1S9S72P016P018P045P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S72P016P018P045N015: std_logic_vector(   0 downto 0);
        signal cVar1S11S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S15S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S16S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S17S72P016P018N045P013: std_logic_vector(   0 downto 0);
        signal cVar1S18S72P016P033P041P011: std_logic_vector(   0 downto 0);
        signal cVar1S19S72P016P033P041P011: std_logic_vector(   0 downto 0);
        signal cVar1S20S72P016P033N041P009: std_logic_vector(   0 downto 0);
        signal cVar1S21S72P016P033N041P009: std_logic_vector(   0 downto 0);
        signal cVar1S22S72P016P033N041P009: std_logic_vector(   0 downto 0);
        signal cVar1S23S72P016P033N041N009: std_logic_vector(   0 downto 0);
        signal cVar1S24S72P016P033N041N009: std_logic_vector(   0 downto 0);
        signal cVar1S25S72P016P033P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S26S72P016P033P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S27S72P016P033P069N068: std_logic_vector(   0 downto 0);
        signal cVar1S28S72P016P033P069N068: std_logic_vector(   0 downto 0);
        signal cVar1S29S72P016P033P069N068: std_logic_vector(   0 downto 0);
        signal cVar1S30S72P016P033P069P067: std_logic_vector(   0 downto 0);
        signal cVar1S0S73P047P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S73P047P006N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S73P047N006P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S73P047N006P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S4S73P047N006N008P007: std_logic_vector(   0 downto 0);
        signal cVar1S5S73P047N006N008N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S73P047N006N008N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S73P047N006N008N007: std_logic_vector(   0 downto 0);
        signal cVar1S8S73N047P031P013P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S73N047P031P013P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S73N047P031P013N056: std_logic_vector(   0 downto 0);
        signal cVar1S11S73N047P031P013N056: std_logic_vector(   0 downto 0);
        signal cVar1S12S73N047P031P013N056: std_logic_vector(   0 downto 0);
        signal cVar1S13S73N047P031N013P011: std_logic_vector(   0 downto 0);
        signal cVar1S14S73N047P031N013P011: std_logic_vector(   0 downto 0);
        signal cVar1S15S73N047P031N013N011: std_logic_vector(   0 downto 0);
        signal cVar1S16S73N047P031N013N011: std_logic_vector(   0 downto 0);
        signal cVar1S17S73N047N031P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S18S73N047N031P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S19S73N047N031P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S20S73N047N031P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S21S73N047N031P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S22S73N047N031P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S23S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S24S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S25S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S26S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S27S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S28S73N047N031N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S0S74P064P066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S1S74P064P066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S74P064P066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S74P064P066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S4S74P064P066P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S5S74P064P066P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S6S74P064P066P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S7S74P064P066N027P041: std_logic_vector(   0 downto 0);
        signal cVar1S8S74P064P066N027P041: std_logic_vector(   0 downto 0);
        signal cVar1S9S74P064P066N027P041: std_logic_vector(   0 downto 0);
        signal cVar1S10S74P064P066N027P041: std_logic_vector(   0 downto 0);
        signal cVar1S11S74P064P066N027N041: std_logic_vector(   0 downto 0);
        signal cVar1S12S74P064P066N027N041: std_logic_vector(   0 downto 0);
        signal cVar1S13S74P064P066N027N041: std_logic_vector(   0 downto 0);
        signal cVar1S14S74P064P066N027N041: std_logic_vector(   0 downto 0);
        signal cVar1S15S74P064P066P006P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S74P064P066P006P059: std_logic_vector(   0 downto 0);
        signal cVar1S17S74P064P066P006P059: std_logic_vector(   0 downto 0);
        signal cVar1S18S74P064P066P006P035: std_logic_vector(   0 downto 0);
        signal cVar1S19S74P064P066P006P035: std_logic_vector(   0 downto 0);
        signal cVar1S20S74P064P011P042P017nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S74P064P011N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S22S74P064P011N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S23S74P064P011N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S74P064P011N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S74P064P011P017P054nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S74P064P011P017N054: std_logic_vector(   0 downto 0);
        signal cVar1S27S74P064P011P017N054: std_logic_vector(   0 downto 0);
        signal cVar1S28S74P064P011N017P009: std_logic_vector(   0 downto 0);
        signal cVar1S29S74P064P011N017N009: std_logic_vector(   0 downto 0);
        signal cVar1S0S75P029P011P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S75P029P011N051P054: std_logic_vector(   0 downto 0);
        signal cVar1S2S75P029P011N051P054: std_logic_vector(   0 downto 0);
        signal cVar1S3S75P029P011N051N054: std_logic_vector(   0 downto 0);
        signal cVar1S4S75P029N011P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S75P029N011P010N052: std_logic_vector(   0 downto 0);
        signal cVar1S6S75P029N011N010P009: std_logic_vector(   0 downto 0);
        signal cVar1S7S75P029N011N010P009: std_logic_vector(   0 downto 0);
        signal cVar1S8S75P029N011N010P009: std_logic_vector(   0 downto 0);
        signal cVar1S9S75P029N011N010N009: std_logic_vector(   0 downto 0);
        signal cVar1S10S75P029N011N010N009: std_logic_vector(   0 downto 0);
        signal cVar1S11S75N029P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S75N029P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S13S75N029P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S14S75N029P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S15S75N029P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S16S75N029P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S17S75N029P041N020P005: std_logic_vector(   0 downto 0);
        signal cVar1S18S75N029P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S19S75N029P041N020N005: std_logic_vector(   0 downto 0);
        signal cVar1S20S75N029N041P045P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S75N029N041P045N023: std_logic_vector(   0 downto 0);
        signal cVar1S22S75N029N041P045N023: std_logic_vector(   0 downto 0);
        signal cVar1S23S75N029N041P045N023: std_logic_vector(   0 downto 0);
        signal cVar1S24S75N029N041N045P027: std_logic_vector(   0 downto 0);
        signal cVar1S25S75N029N041N045P027: std_logic_vector(   0 downto 0);
        signal cVar1S26S75N029N041N045N027: std_logic_vector(   0 downto 0);
        signal cVar1S27S75N029N041N045N027: std_logic_vector(   0 downto 0);
        signal cVar1S0S76P064P027P066P009: std_logic_vector(   0 downto 0);
        signal cVar1S1S76P064P027P066P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S76P064P027P066N009: std_logic_vector(   0 downto 0);
        signal cVar1S3S76P064P027P066P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S76P064P027P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S5S76P064P027P066P068: std_logic_vector(   0 downto 0);
        signal cVar1S6S76P064N027P041P020: std_logic_vector(   0 downto 0);
        signal cVar1S7S76P064N027P041P020: std_logic_vector(   0 downto 0);
        signal cVar1S8S76P064N027P041P020: std_logic_vector(   0 downto 0);
        signal cVar1S9S76P064N027P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S10S76P064N027P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S11S76P064N027P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S12S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S13S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S14S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S76P064N027N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S18S76P064P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S76P064N042P008P027: std_logic_vector(   0 downto 0);
        signal cVar1S20S76P064N042P008P027: std_logic_vector(   0 downto 0);
        signal cVar1S21S76P064N042P008P027: std_logic_vector(   0 downto 0);
        signal cVar1S22S76P064N042P008P027: std_logic_vector(   0 downto 0);
        signal cVar1S23S76P064N042P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S24S76P064N042P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S0S77P017P064P034P035: std_logic_vector(   0 downto 0);
        signal cVar1S1S77P017P064P034P035: std_logic_vector(   0 downto 0);
        signal cVar1S2S77P017P064P034P035: std_logic_vector(   0 downto 0);
        signal cVar1S3S77P017P064N034P020: std_logic_vector(   0 downto 0);
        signal cVar1S4S77P017P064N034P020: std_logic_vector(   0 downto 0);
        signal cVar1S5S77P017P064N034P020: std_logic_vector(   0 downto 0);
        signal cVar1S6S77P017P064N034N020: std_logic_vector(   0 downto 0);
        signal cVar1S7S77P017P064N034N020: std_logic_vector(   0 downto 0);
        signal cVar1S8S77P017P064N034N020: std_logic_vector(   0 downto 0);
        signal cVar1S9S77P017P064P050P016nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S77P017P064N050P020: std_logic_vector(   0 downto 0);
        signal cVar1S11S77P017P064N050P020: std_logic_vector(   0 downto 0);
        signal cVar1S12S77P017P064N050P020: std_logic_vector(   0 downto 0);
        signal cVar1S13S77N017P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S77N017P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S15S77N017P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S16S77N017P041N020P015: std_logic_vector(   0 downto 0);
        signal cVar1S17S77N017P041N020P015: std_logic_vector(   0 downto 0);
        signal cVar1S18S77N017P041N020P015: std_logic_vector(   0 downto 0);
        signal cVar1S19S77N017P041N020P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S77N017N041P062P027: std_logic_vector(   0 downto 0);
        signal cVar1S21S77N017N041P062P027: std_logic_vector(   0 downto 0);
        signal cVar1S22S77N017N041P062P027: std_logic_vector(   0 downto 0);
        signal cVar1S23S77N017N041P062N027: std_logic_vector(   0 downto 0);
        signal cVar1S24S77N017N041P062N027: std_logic_vector(   0 downto 0);
        signal cVar1S25S77N017N041P062N027: std_logic_vector(   0 downto 0);
        signal cVar1S26S77N017N041P062N027: std_logic_vector(   0 downto 0);
        signal cVar1S27S77N017N041P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S28S77N017N041P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S29S77N017N041P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S30S77N017N041P062P010: std_logic_vector(   0 downto 0);
        signal cVar1S0S78P062P063P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S1S78P062P063P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S2S78P062P063P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S78P062P063P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S78P062P063P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S5S78P062P063P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S6S78P062P063N007P029: std_logic_vector(   0 downto 0);
        signal cVar1S7S78P062P063N007P029: std_logic_vector(   0 downto 0);
        signal cVar1S8S78P062P063N007P029: std_logic_vector(   0 downto 0);
        signal cVar1S9S78P062P063N007N029: std_logic_vector(   0 downto 0);
        signal cVar1S10S78P062P063N007N029: std_logic_vector(   0 downto 0);
        signal cVar1S11S78P062P063N007N029: std_logic_vector(   0 downto 0);
        signal cVar1S12S78P062P063N007N029: std_logic_vector(   0 downto 0);
        signal cVar1S13S78P062P063P035P058: std_logic_vector(   0 downto 0);
        signal cVar1S14S78P062P063P035P058: std_logic_vector(   0 downto 0);
        signal cVar1S15S78P062P063P035P058: std_logic_vector(   0 downto 0);
        signal cVar1S16S78P062P063N035P034: std_logic_vector(   0 downto 0);
        signal cVar1S17S78P062P063N035P034: std_logic_vector(   0 downto 0);
        signal cVar1S18S78P062P063N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S19S78P062P063N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S20S78P062P063N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S21S78P062P026P027P060: std_logic_vector(   0 downto 0);
        signal cVar1S22S78P062P026P027P060: std_logic_vector(   0 downto 0);
        signal cVar1S23S78P062P026P027P060: std_logic_vector(   0 downto 0);
        signal cVar1S24S78P062P026P027N060: std_logic_vector(   0 downto 0);
        signal cVar1S25S78P062P026P027N060: std_logic_vector(   0 downto 0);
        signal cVar1S26S78P062P026P027N060: std_logic_vector(   0 downto 0);
        signal cVar1S27S78P062P026P027N060: std_logic_vector(   0 downto 0);
        signal cVar1S28S78P062P026P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S79P051P008P065P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S79P051P008P065N028: std_logic_vector(   0 downto 0);
        signal cVar1S2S79P051P008P065N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S79P051N008P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S79P051N008N042P009: std_logic_vector(   0 downto 0);
        signal cVar1S5S79P051N008N042P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S79P051N008N042P009: std_logic_vector(   0 downto 0);
        signal cVar1S7S79P051N008N042N009: std_logic_vector(   0 downto 0);
        signal cVar1S8S79P051N008N042N009: std_logic_vector(   0 downto 0);
        signal cVar1S9S79P051N008N042N009: std_logic_vector(   0 downto 0);
        signal cVar1S10S79N051P041P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S79N051P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S12S79N051P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S13S79N051P041P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S14S79N051P041N020P001nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S79N051P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S16S79N051P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S17S79N051P041N020N001: std_logic_vector(   0 downto 0);
        signal cVar1S18S79N051N041P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S19S79N051N041P047P026: std_logic_vector(   0 downto 0);
        signal cVar1S20S79N051N041P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S21S79N051N041P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S22S79N051N041P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S23S79N051N041P047N026: std_logic_vector(   0 downto 0);
        signal cVar1S24S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S25S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S26S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S27S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S28S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S29S79N051N041N047P049: std_logic_vector(   0 downto 0);
        signal cVar1S0S80P040P002P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S80P040P002N021P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S80P040P002N021N041: std_logic_vector(   0 downto 0);
        signal cVar1S3S80P040N002P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S80P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S5S80P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S6S80P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S7S80P040N002N057N004: std_logic_vector(   0 downto 0);
        signal cVar1S8S80P040N002N057N004: std_logic_vector(   0 downto 0);
        signal cVar1S9S80P040N002N057N004: std_logic_vector(   0 downto 0);
        signal cVar1S10S80N040P021P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S11S80N040P021P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S12S80N040P021P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S13S80N040P021P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S14S80N040P021N007P028: std_logic_vector(   0 downto 0);
        signal cVar1S15S80N040P021N007P028: std_logic_vector(   0 downto 0);
        signal cVar1S16S80N040P021N007N028: std_logic_vector(   0 downto 0);
        signal cVar1S17S80N040P021N007N028: std_logic_vector(   0 downto 0);
        signal cVar1S18S80N040P021N007N028: std_logic_vector(   0 downto 0);
        signal cVar1S19S80N040P021N007N028: std_logic_vector(   0 downto 0);
        signal cVar1S20S80N040P021P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S80N040P021N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S22S80N040P021N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S23S80N040P021N042N003: std_logic_vector(   0 downto 0);
        signal cVar1S24S80N040P021N042N003: std_logic_vector(   0 downto 0);
        signal cVar1S0S81P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S81P040N002P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S81P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S3S81P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S4S81P040N002N057P004: std_logic_vector(   0 downto 0);
        signal cVar1S5S81P040N002N057N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S81N040P028P029P053: std_logic_vector(   0 downto 0);
        signal cVar1S7S81N040P028P029P053: std_logic_vector(   0 downto 0);
        signal cVar1S8S81N040P028P029N053: std_logic_vector(   0 downto 0);
        signal cVar1S9S81N040P028P029N053: std_logic_vector(   0 downto 0);
        signal cVar1S10S81N040N028P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S11S81N040N028P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S81N040N028P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S13S81N040N028P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S14S81N040N028P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S15S81N040N028P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S16S81N040N028P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S17S81N040N028N029P007: std_logic_vector(   0 downto 0);
        signal cVar1S18S81N040N028N029P007: std_logic_vector(   0 downto 0);
        signal cVar1S19S81N040N028N029P007: std_logic_vector(   0 downto 0);
        signal cVar1S20S81N040N028N029N007: std_logic_vector(   0 downto 0);
        signal cVar1S21S81N040N028N029N007: std_logic_vector(   0 downto 0);
        signal cVar1S22S81N040N028N029N007: std_logic_vector(   0 downto 0);
        signal cVar1S0S82P062P007P025P009: std_logic_vector(   0 downto 0);
        signal cVar1S1S82P062P007P025P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S82P062P007N025P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S82P062P007N025P003: std_logic_vector(   0 downto 0);
        signal cVar1S4S82P062P007N025N003: std_logic_vector(   0 downto 0);
        signal cVar1S5S82P062P007N025N003: std_logic_vector(   0 downto 0);
        signal cVar1S6S82P062P007N025N003: std_logic_vector(   0 downto 0);
        signal cVar1S7S82P062P007N025N003: std_logic_vector(   0 downto 0);
        signal cVar1S8S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S9S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S10S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S11S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S12S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S82P062N007P015P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S82P062N007P015P029: std_logic_vector(   0 downto 0);
        signal cVar1S16S82P062N007P015N029: std_logic_vector(   0 downto 0);
        signal cVar1S17S82P062N007P015N029: std_logic_vector(   0 downto 0);
        signal cVar1S18S82P062N007P015N029: std_logic_vector(   0 downto 0);
        signal cVar1S19S82P062P026P029P050: std_logic_vector(   0 downto 0);
        signal cVar1S20S82P062P026P029P050: std_logic_vector(   0 downto 0);
        signal cVar1S21S82P062P026P029N050: std_logic_vector(   0 downto 0);
        signal cVar1S22S82P062P026P029N050: std_logic_vector(   0 downto 0);
        signal cVar1S23S82P062P026P029P036: std_logic_vector(   0 downto 0);
        signal cVar1S24S82P062P026P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S83P007P025P046P011nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S83P007P025N046P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S83P007P025N046P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S83P007P025N046P009: std_logic_vector(   0 downto 0);
        signal cVar1S4S83P007N025P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S83P007N025P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S6S83P007N025P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S7S83P007N025P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S83P007N025P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S83P007N025P034P019: std_logic_vector(   0 downto 0);
        signal cVar1S10S83P007N025P034N019: std_logic_vector(   0 downto 0);
        signal cVar1S11S83N007P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S83N007P040N002P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S83N007P040N002N047: std_logic_vector(   0 downto 0);
        signal cVar1S14S83N007P040N002N047: std_logic_vector(   0 downto 0);
        signal cVar1S15S83N007P040N002N047: std_logic_vector(   0 downto 0);
        signal cVar1S16S83N007N040P015P038: std_logic_vector(   0 downto 0);
        signal cVar1S17S83N007N040P015P038: std_logic_vector(   0 downto 0);
        signal cVar1S18S83N007N040N015P034: std_logic_vector(   0 downto 0);
        signal cVar1S19S83N007N040N015P034: std_logic_vector(   0 downto 0);
        signal cVar1S20S83N007N040N015N034: std_logic_vector(   0 downto 0);
        signal cVar1S21S83N007N040N015N034: std_logic_vector(   0 downto 0);
        signal cVar1S22S83N007N040N015N034: std_logic_vector(   0 downto 0);
        signal cVar1S23S83N007N040N015N034: std_logic_vector(   0 downto 0);
        signal cVar1S0S84P040P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S84P040P021N002P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S84P040P021N002P012: std_logic_vector(   0 downto 0);
        signal cVar1S3S84P040P021N002P012: std_logic_vector(   0 downto 0);
        signal cVar1S4S84P040N021P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S84P040N021N057P008: std_logic_vector(   0 downto 0);
        signal cVar1S6S84P040N021N057P008: std_logic_vector(   0 downto 0);
        signal cVar1S7S84P040N021N057P008: std_logic_vector(   0 downto 0);
        signal cVar1S8S84N040P007P025P046: std_logic_vector(   0 downto 0);
        signal cVar1S9S84N040P007P025N046: std_logic_vector(   0 downto 0);
        signal cVar1S10S84N040P007P025N046: std_logic_vector(   0 downto 0);
        signal cVar1S11S84N040P007P025N046: std_logic_vector(   0 downto 0);
        signal cVar1S12S84N040P007N025P055: std_logic_vector(   0 downto 0);
        signal cVar1S13S84N040P007N025P055: std_logic_vector(   0 downto 0);
        signal cVar1S14S84N040P007N025P055: std_logic_vector(   0 downto 0);
        signal cVar1S15S84N040P007N025P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S17S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S18S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S19S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S20S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S21S84N040N007P015P001: std_logic_vector(   0 downto 0);
        signal cVar1S22S84N040N007P015P035: std_logic_vector(   0 downto 0);
        signal cVar1S23S84N040N007P015P035: std_logic_vector(   0 downto 0);
        signal cVar1S24S84N040N007P015P035: std_logic_vector(   0 downto 0);
        signal cVar1S25S84N040N007P015N035: std_logic_vector(   0 downto 0);
        signal cVar1S26S84N040N007P015N035: std_logic_vector(   0 downto 0);
        signal cVar1S27S84N040N007P015N035: std_logic_vector(   0 downto 0);
        signal cVar1S28S84N040N007P015N035: std_logic_vector(   0 downto 0);
        signal cVar1S0S85P015P032P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S85P015P032N005P003: std_logic_vector(   0 downto 0);
        signal cVar1S2S85P015P032N005P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S85P015N032P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S4S85P015N032P011P008: std_logic_vector(   0 downto 0);
        signal cVar1S5S85P015N032N011P000: std_logic_vector(   0 downto 0);
        signal cVar1S6S85P015N032N011P000: std_logic_vector(   0 downto 0);
        signal cVar1S7S85P015N032N011P000: std_logic_vector(   0 downto 0);
        signal cVar1S8S85P015N032N011N000: std_logic_vector(   0 downto 0);
        signal cVar1S9S85P015N032N011N000: std_logic_vector(   0 downto 0);
        signal cVar1S10S85N015P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S85N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S12S85N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S85N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S85N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S85N015N021P044P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S85N015N021P044N004: std_logic_vector(   0 downto 0);
        signal cVar1S17S85N015N021P044N004: std_logic_vector(   0 downto 0);
        signal cVar1S18S85N015N021P044N004: std_logic_vector(   0 downto 0);
        signal cVar1S19S85N015N021N044P005: std_logic_vector(   0 downto 0);
        signal cVar1S20S85N015N021N044P005: std_logic_vector(   0 downto 0);
        signal cVar1S21S85N015N021N044P005: std_logic_vector(   0 downto 0);
        signal cVar1S22S85N015N021N044P005: std_logic_vector(   0 downto 0);
        signal cVar1S23S85N015N021N044P005: std_logic_vector(   0 downto 0);
        signal cVar1S0S86P021P038P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S86P021P038N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S86P021P038N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S86P021P038N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S86P021N038P010P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S86P021N038P010N042: std_logic_vector(   0 downto 0);
        signal cVar1S6S86P021N038P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S86N021P020P039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S86N021P020P039N003: std_logic_vector(   0 downto 0);
        signal cVar1S9S86N021P020P039N003: std_logic_vector(   0 downto 0);
        signal cVar1S10S86N021P020P039N003: std_logic_vector(   0 downto 0);
        signal cVar1S11S86N021P020N039P031: std_logic_vector(   0 downto 0);
        signal cVar1S12S86N021P020N039P031: std_logic_vector(   0 downto 0);
        signal cVar1S13S86N021P020N039P031: std_logic_vector(   0 downto 0);
        signal cVar1S14S86N021P020N039P031: std_logic_vector(   0 downto 0);
        signal cVar1S15S86N021N020P002P015: std_logic_vector(   0 downto 0);
        signal cVar1S16S86N021N020P002P015: std_logic_vector(   0 downto 0);
        signal cVar1S17S86N021N020P002P015: std_logic_vector(   0 downto 0);
        signal cVar1S18S86N021N020P002N015: std_logic_vector(   0 downto 0);
        signal cVar1S19S86N021N020P002N015: std_logic_vector(   0 downto 0);
        signal cVar1S20S86N021N020P002N015: std_logic_vector(   0 downto 0);
        signal cVar1S21S86N021N020P002P004: std_logic_vector(   0 downto 0);
        signal cVar1S22S86N021N020P002P004: std_logic_vector(   0 downto 0);
        signal cVar1S23S86N021N020P002N004: std_logic_vector(   0 downto 0);
        signal cVar1S24S86N021N020P002N004: std_logic_vector(   0 downto 0);
        signal cVar1S0S87P015P055P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S87P015P055P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S2S87P015P055P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S3S87P015P055P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S4S87P015N055P021P020: std_logic_vector(   0 downto 0);
        signal cVar1S5S87P015N055P021P020: std_logic_vector(   0 downto 0);
        signal cVar1S6S87P015N055P021N020: std_logic_vector(   0 downto 0);
        signal cVar1S7S87P015N055P021N020: std_logic_vector(   0 downto 0);
        signal cVar1S8S87P015N055P021N020: std_logic_vector(   0 downto 0);
        signal cVar1S9S87P015N055P021P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S87P015N055P021N066: std_logic_vector(   0 downto 0);
        signal cVar1S11S87P015N055P021N066: std_logic_vector(   0 downto 0);
        signal cVar1S12S87N015P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S87N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S87N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S87N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S16S87N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S87N015P021N038P014: std_logic_vector(   0 downto 0);
        signal cVar1S18S87N015N021P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S87N015N021P020N039: std_logic_vector(   0 downto 0);
        signal cVar1S20S87N015N021P020N039: std_logic_vector(   0 downto 0);
        signal cVar1S21S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S22S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S23S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S24S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S25S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S26S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S27S87N015N021N020P057: std_logic_vector(   0 downto 0);
        signal cVar1S0S88P015P057P055P039: std_logic_vector(   0 downto 0);
        signal cVar1S1S88P015P057P055P039: std_logic_vector(   0 downto 0);
        signal cVar1S2S88P015P057P055N039: std_logic_vector(   0 downto 0);
        signal cVar1S3S88P015P057P055N039: std_logic_vector(   0 downto 0);
        signal cVar1S4S88P015P057P055N039: std_logic_vector(   0 downto 0);
        signal cVar1S5S88P015P057P055N039: std_logic_vector(   0 downto 0);
        signal cVar1S6S88P015P057P055P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S88P015P057P055N069: std_logic_vector(   0 downto 0);
        signal cVar1S8S88P015P057P055N069: std_logic_vector(   0 downto 0);
        signal cVar1S9S88P015P057P055N069: std_logic_vector(   0 downto 0);
        signal cVar1S10S88P015P057P010P055: std_logic_vector(   0 downto 0);
        signal cVar1S11S88P015P057P010P055: std_logic_vector(   0 downto 0);
        signal cVar1S12S88P015P057N010P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S88P015P057N010P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S88P015P057N010N013: std_logic_vector(   0 downto 0);
        signal cVar1S15S88P015P057N010N013: std_logic_vector(   0 downto 0);
        signal cVar1S16S88P015P057N010N013: std_logic_vector(   0 downto 0);
        signal cVar1S17S88P015P057N010N013: std_logic_vector(   0 downto 0);
        signal cVar1S18S88P015P055P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S88P015P055P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S20S88P015P055P061N032: std_logic_vector(   0 downto 0);
        signal cVar1S21S88P015N055P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S88P015N055P020N002: std_logic_vector(   0 downto 0);
        signal cVar1S23S88P015N055N020P009: std_logic_vector(   0 downto 0);
        signal cVar1S24S88P015N055N020P009: std_logic_vector(   0 downto 0);
        signal cVar1S25S88P015N055N020N009: std_logic_vector(   0 downto 0);
        signal cVar1S26S88P015N055N020N009: std_logic_vector(   0 downto 0);
        signal cVar1S0S89P015P013P008P059: std_logic_vector(   0 downto 0);
        signal cVar1S1S89P015P013P008P059: std_logic_vector(   0 downto 0);
        signal cVar1S2S89P015P013P008P059: std_logic_vector(   0 downto 0);
        signal cVar1S3S89P015P013P008N059: std_logic_vector(   0 downto 0);
        signal cVar1S4S89P015P013P008N059: std_logic_vector(   0 downto 0);
        signal cVar1S5S89P015P013P008N059: std_logic_vector(   0 downto 0);
        signal cVar1S6S89P015P013P008P019: std_logic_vector(   0 downto 0);
        signal cVar1S7S89P015P013P008P019: std_logic_vector(   0 downto 0);
        signal cVar1S8S89P015P013P008N019: std_logic_vector(   0 downto 0);
        signal cVar1S9S89P015P013P059P055: std_logic_vector(   0 downto 0);
        signal cVar1S10S89P015P013P059N055: std_logic_vector(   0 downto 0);
        signal cVar1S11S89P015P013P059N055: std_logic_vector(   0 downto 0);
        signal cVar1S12S89P015P013P059N055: std_logic_vector(   0 downto 0);
        signal cVar1S13S89P015P013P059N055: std_logic_vector(   0 downto 0);
        signal cVar1S14S89P015P013P059P061: std_logic_vector(   0 downto 0);
        signal cVar1S15S89P015P013P059P061: std_logic_vector(   0 downto 0);
        signal cVar1S16S89N015P039P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S89N015P039P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S18S89N015P039P020N003: std_logic_vector(   0 downto 0);
        signal cVar1S19S89N015P039N020P017: std_logic_vector(   0 downto 0);
        signal cVar1S20S89N015P039N020P017: std_logic_vector(   0 downto 0);
        signal cVar1S21S89N015N039P044P025: std_logic_vector(   0 downto 0);
        signal cVar1S22S89N015N039P044N025: std_logic_vector(   0 downto 0);
        signal cVar1S23S89N015N039P044N025: std_logic_vector(   0 downto 0);
        signal cVar1S24S89N015N039P044N025: std_logic_vector(   0 downto 0);
        signal cVar1S25S89N015N039N044P038: std_logic_vector(   0 downto 0);
        signal cVar1S26S89N015N039N044P038: std_logic_vector(   0 downto 0);
        signal cVar1S27S89N015N039N044N038: std_logic_vector(   0 downto 0);
        signal cVar1S28S89N015N039N044N038: std_logic_vector(   0 downto 0);
        signal cVar1S29S89N015N039N044N038: std_logic_vector(   0 downto 0);
        signal cVar1S0S90P020P039P010P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S90P020P039P010N003: std_logic_vector(   0 downto 0);
        signal cVar1S2S90P020N039P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S90P020N039N025P031: std_logic_vector(   0 downto 0);
        signal cVar1S4S90P020N039N025P031: std_logic_vector(   0 downto 0);
        signal cVar1S5S90N020P040P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S90N020P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S7S90N020P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S8S90N020P040P021N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S90N020P040N021P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S90N020P040N021N057: std_logic_vector(   0 downto 0);
        signal cVar1S11S90N020N040P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S12S90N020N040P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S13S90N020N040P039P045: std_logic_vector(   0 downto 0);
        signal cVar1S14S90N020N040P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S15S90N020N040P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S16S90N020N040P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S17S90N020N040P039N045: std_logic_vector(   0 downto 0);
        signal cVar1S18S90N020N040P039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S91P020P039P010P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S91P020P039P010N003: std_logic_vector(   0 downto 0);
        signal cVar1S2S91P020N039P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S91P020N039N025P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S91P020N039N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S5S91P020N039N025N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S91N020P045P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S91N020P045P004P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S91N020P045N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S9S91N020P045N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S10S91N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S11S91N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S12S91N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S13S91N020N045P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S91N020N045P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S15S91N020N045P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S16S91N020N045N040P055: std_logic_vector(   0 downto 0);
        signal cVar1S17S91N020N045N040P055: std_logic_vector(   0 downto 0);
        signal cVar1S18S91N020N045N040P055: std_logic_vector(   0 downto 0);
        signal cVar1S19S91N020N045N040N055: std_logic_vector(   0 downto 0);
        signal cVar1S20S91N020N045N040N055: std_logic_vector(   0 downto 0);
        signal cVar1S21S91N020N045N040N055: std_logic_vector(   0 downto 0);
        signal cVar1S0S92P020P039P010P003nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S92P020P039P010N003: std_logic_vector(   0 downto 0);
        signal cVar1S2S92P020P039P010N003: std_logic_vector(   0 downto 0);
        signal cVar1S3S92P020N039P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S92P020N039N025P031: std_logic_vector(   0 downto 0);
        signal cVar1S5S92P020N039N025P031: std_logic_vector(   0 downto 0);
        signal cVar1S6S92N020P045P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S92N020P045P004P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S92N020P045N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S9S92N020P045N004P006: std_logic_vector(   0 downto 0);
        signal cVar1S10S92N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S11S92N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S12S92N020P045N004N006: std_logic_vector(   0 downto 0);
        signal cVar1S13S92N020N045P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S92N020N045P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S15S92N020N045P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S16S92N020N045N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S17S92N020N045N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S18S92N020N045N040P044: std_logic_vector(   0 downto 0);
        signal cVar1S19S92N020N045N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S20S92N020N045N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S21S92N020N045N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S22S92N020N045N040N044: std_logic_vector(   0 downto 0);
        signal cVar1S0S93P040P002P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S93P040P002N021P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S93P040P002N021N041: std_logic_vector(   0 downto 0);
        signal cVar1S3S93P040N002P004P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S93P040N002P004N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S93P040N002P004N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S93P040N002N004P000nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S93P040N002N004N000: std_logic_vector(   0 downto 0);
        signal cVar1S8S93P040N002N004N000: std_logic_vector(   0 downto 0);
        signal cVar1S9S93P040N002N004N000: std_logic_vector(   0 downto 0);
        signal cVar1S10S93N040P045P022P019nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S93N040P045P022N019: std_logic_vector(   0 downto 0);
        signal cVar1S12S93N040P045P022N019: std_logic_vector(   0 downto 0);
        signal cVar1S13S93N040P045P022N019: std_logic_vector(   0 downto 0);
        signal cVar1S14S93N040P045N022P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S93N040P045N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S93N040P045N022N023: std_logic_vector(   0 downto 0);
        signal cVar1S17S93N040N045P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S18S93N040N045P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S19S93N040N045P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S20S93N040N045P020N039: std_logic_vector(   0 downto 0);
        signal cVar1S21S93N040N045P020N039: std_logic_vector(   0 downto 0);
        signal cVar1S22S93N040N045N020P044: std_logic_vector(   0 downto 0);
        signal cVar1S23S93N040N045N020P044: std_logic_vector(   0 downto 0);
        signal cVar1S24S93N040N045N020P044: std_logic_vector(   0 downto 0);
        signal cVar1S25S93N040N045N020N044: std_logic_vector(   0 downto 0);
        signal cVar1S26S93N040N045N020N044: std_logic_vector(   0 downto 0);
        signal cVar1S27S93N040N045N020N044: std_logic_vector(   0 downto 0);
        signal cVar1S28S93N040N045N020N044: std_logic_vector(   0 downto 0);
        signal cVar1S0S94P040P002P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S94P040P002N021P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S94P040P002N021N041: std_logic_vector(   0 downto 0);
        signal cVar1S3S94P040N002P004P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S94P040N002P004N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S94P040N002P004N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S94P040N002N004P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S94N040P044P006P048: std_logic_vector(   0 downto 0);
        signal cVar1S8S94N040P044P006P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S94N040P044N006P023: std_logic_vector(   0 downto 0);
        signal cVar1S10S94N040P044N006P023: std_logic_vector(   0 downto 0);
        signal cVar1S11S94N040P044N006P023: std_logic_vector(   0 downto 0);
        signal cVar1S12S94N040P044N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S13S94N040P044N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S14S94N040P044N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S15S94N040N044P042P020: std_logic_vector(   0 downto 0);
        signal cVar1S16S94N040N044P042P020: std_logic_vector(   0 downto 0);
        signal cVar1S17S94N040N044P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S18S94N040N044P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S19S94N040N044P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S20S94N040N044P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S21S94N040N044P042P058nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S94N040N044P042N058: std_logic_vector(   0 downto 0);
        signal cVar1S23S94N040N044P042N058: std_logic_vector(   0 downto 0);
        signal cVar1S0S95P044P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S95P044P023N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S95P044P023N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S3S95P044P023N005N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S95P044N023P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S95P044N023N051P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S95P044N023N051N057: std_logic_vector(   0 downto 0);
        signal cVar1S7S95P044N023N051N057: std_logic_vector(   0 downto 0);
        signal cVar1S8S95P044N023N051N057: std_logic_vector(   0 downto 0);
        signal cVar1S9S95P044N023N051N057: std_logic_vector(   0 downto 0);
        signal cVar1S10S95N044P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S95N044P040N002P004: std_logic_vector(   0 downto 0);
        signal cVar1S12S95N044P040N002P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S95N044P040N002P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S95N044P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S95N044P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S16S95N044P040N002N004: std_logic_vector(   0 downto 0);
        signal cVar1S17S95N044N040P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S95N044N040P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S19S95N044N040P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S20S95N044N040P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S21S95N044N040N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S22S95N044N040N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S23S95N044N040N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S24S95N044N040N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S25S95N044N040N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S26S95N044N040N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S27S95N044N040N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S28S95N044N040N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S0S96P044P004P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S96P044P004N023P022: std_logic_vector(   0 downto 0);
        signal cVar1S2S96P044N004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S96P044N004N021P005: std_logic_vector(   0 downto 0);
        signal cVar1S4S96P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S5S96P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S6S96P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S7S96P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S8S96N044P016P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S96N044P016P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S96N044P016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S11S96N044P016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S12S96N044P016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S13S96N044P016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S14S96N044P016N012P053: std_logic_vector(   0 downto 0);
        signal cVar1S15S96N044P016N012P053: std_logic_vector(   0 downto 0);
        signal cVar1S16S96N044P016N012N053: std_logic_vector(   0 downto 0);
        signal cVar1S17S96N044P016N012N053: std_logic_vector(   0 downto 0);
        signal cVar1S18S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S19S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S20S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S21S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S22S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S23S96N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S24S96N044P016P052P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S96N044P016P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S26S96N044P016P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S0S97P044P004P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S97P044P004N023P016: std_logic_vector(   0 downto 0);
        signal cVar1S2S97P044N004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S97P044N004N021P005: std_logic_vector(   0 downto 0);
        signal cVar1S4S97P044N004N021P005: std_logic_vector(   0 downto 0);
        signal cVar1S5S97P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S6S97P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S7S97P044N004N021N005: std_logic_vector(   0 downto 0);
        signal cVar1S8S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S11S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S12S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S13S97N044P016P052P059: std_logic_vector(   0 downto 0);
        signal cVar1S14S97N044P016P052P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S97N044P016P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S16S97N044N016P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S97N044N016P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S97N044N016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S19S97N044N016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S20S97N044N016P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S21S97N044N016N012P053: std_logic_vector(   0 downto 0);
        signal cVar1S22S97N044N016N012P053: std_logic_vector(   0 downto 0);
        signal cVar1S23S97N044N016N012P053: std_logic_vector(   0 downto 0);
        signal cVar1S24S97N044N016N012N053: std_logic_vector(   0 downto 0);
        signal cVar1S25S97N044N016N012N053: std_logic_vector(   0 downto 0);
        signal cVar1S26S97N044N016N012N053: std_logic_vector(   0 downto 0);
        signal cVar1S0S98P016P044P004P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S98P016P044P004N023: std_logic_vector(   0 downto 0);
        signal cVar1S2S98P016P044N004P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S98P016P044N004N047: std_logic_vector(   0 downto 0);
        signal cVar1S4S98P016P044N004N047: std_logic_vector(   0 downto 0);
        signal cVar1S5S98P016P044N004N047: std_logic_vector(   0 downto 0);
        signal cVar1S6S98P016N044P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S98P016N044P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S98P016N044P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S9S98P016N044P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S10S98P016N044P012N056: std_logic_vector(   0 downto 0);
        signal cVar1S11S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S12S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S16S98P016N044N012P032: std_logic_vector(   0 downto 0);
        signal cVar1S17S98P016P021P037P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S98P016P021P037N053: std_logic_vector(   0 downto 0);
        signal cVar1S19S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S23S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S24S98P016P021N037P047: std_logic_vector(   0 downto 0);
        signal cVar1S25S98P016P021P069P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S98P016P021P069N038: std_logic_vector(   0 downto 0);
        signal cVar1S27S98P016P021P069N038: std_logic_vector(   0 downto 0);
        signal cVar1S0S99P044P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S99P044N051P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S99P044N051N057P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S99P044N051N057N032: std_logic_vector(   0 downto 0);
        signal cVar1S4S99P044N051N057N032: std_logic_vector(   0 downto 0);
        signal cVar1S5S99P044N051N057N032: std_logic_vector(   0 downto 0);
        signal cVar1S6S99P044N051N057N032: std_logic_vector(   0 downto 0);
        signal cVar1S7S99N044P062P003P039: std_logic_vector(   0 downto 0);
        signal cVar1S8S99N044P062P003P039: std_logic_vector(   0 downto 0);
        signal cVar1S9S99N044P062P003N039: std_logic_vector(   0 downto 0);
        signal cVar1S10S99N044P062P003N039: std_logic_vector(   0 downto 0);
        signal cVar1S11S99N044P062P003N039: std_logic_vector(   0 downto 0);
        signal cVar1S12S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S13S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S14S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S15S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S16S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S17S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S18S99N044P062N003P042: std_logic_vector(   0 downto 0);
        signal cVar1S19S99N044P062P063P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S99N044P062P063N053: std_logic_vector(   0 downto 0);
        signal cVar1S21S99N044P062P063N053: std_logic_vector(   0 downto 0);
        signal cVar1S22S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S23S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S24S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S25S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S26S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S27S99N044P062N063P009: std_logic_vector(   0 downto 0);
        signal cVar1S0S100P015P044P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S100P015P044N004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S100P015P044N004N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S100P015P044N004N021: std_logic_vector(   0 downto 0);
        signal cVar1S4S100P015P044N004N021: std_logic_vector(   0 downto 0);
        signal cVar1S5S100P015N044P062P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S100P015N044P062N045: std_logic_vector(   0 downto 0);
        signal cVar1S7S100P015N044P062N045: std_logic_vector(   0 downto 0);
        signal cVar1S8S100P015N044P062N045: std_logic_vector(   0 downto 0);
        signal cVar1S9S100P015N044P062P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S100P015N044P062P017: std_logic_vector(   0 downto 0);
        signal cVar1S11S100P015N044P062P017: std_logic_vector(   0 downto 0);
        signal cVar1S12S100P015N044P062P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S100P015N044P062N017: std_logic_vector(   0 downto 0);
        signal cVar1S14S100P015N044P062N017: std_logic_vector(   0 downto 0);
        signal cVar1S15S100P015N044P062N017: std_logic_vector(   0 downto 0);
        signal cVar1S16S100P015N044P062N017: std_logic_vector(   0 downto 0);
        signal cVar1S17S100P015P013P056P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S100P015P013P056P032: std_logic_vector(   0 downto 0);
        signal cVar1S19S100P015P013P056N032: std_logic_vector(   0 downto 0);
        signal cVar1S20S100P015P013P056N032: std_logic_vector(   0 downto 0);
        signal cVar1S21S100P015P013P056N032: std_logic_vector(   0 downto 0);
        signal cVar1S22S100P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S23S100P015P013P056N068: std_logic_vector(   0 downto 0);
        signal cVar1S24S100P015P013P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S25S100P015P013N025P066: std_logic_vector(   0 downto 0);
        signal cVar1S26S100P015P013N025P066: std_logic_vector(   0 downto 0);
        signal cVar1S27S100P015P013N025P066: std_logic_vector(   0 downto 0);
        signal cVar1S28S100P015P013N025N066: std_logic_vector(   0 downto 0);
        signal cVar1S29S100P015P013N025N066: std_logic_vector(   0 downto 0);
        signal cVar1S30S100P015P013N025N066: std_logic_vector(   0 downto 0);
        signal cVar1S0S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S1S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S4S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S5S101P015P013P056P068: std_logic_vector(   0 downto 0);
        signal cVar1S6S101P015P013P056P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S101P015P013P056N050: std_logic_vector(   0 downto 0);
        signal cVar1S8S101P015P013P056N050: std_logic_vector(   0 downto 0);
        signal cVar1S9S101P015P013P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S101P015P013N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S101P015P013N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S12S101P015P013N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S13S101P015P013N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S14S101N015P044P025P017: std_logic_vector(   0 downto 0);
        signal cVar1S15S101N015P044P025P017psss: std_logic_vector(   0 downto 0);
        signal cVar1S16S101N015P044N025P005: std_logic_vector(   0 downto 0);
        signal cVar1S17S101N015P044N025N005: std_logic_vector(   0 downto 0);
        signal cVar1S18S101N015P044N025N005: std_logic_vector(   0 downto 0);
        signal cVar1S19S101N015P044N025N005: std_logic_vector(   0 downto 0);
        signal cVar1S20S101N015N044P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S21S101N015N044P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S22S101N015N044P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S23S101N015N044P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S24S101N015N044P016P052: std_logic_vector(   0 downto 0);
        signal cVar1S25S101N015N044N016P012: std_logic_vector(   0 downto 0);
        signal cVar1S26S101N015N044N016P012: std_logic_vector(   0 downto 0);
        signal cVar1S27S101N015N044N016P012: std_logic_vector(   0 downto 0);
        signal cVar1S28S101N015N044N016P012: std_logic_vector(   0 downto 0);
        signal cVar1S29S101N015N044N016N012: std_logic_vector(   0 downto 0);
        signal cVar1S30S101N015N044N016N012: std_logic_vector(   0 downto 0);
        signal cVar1S0S102P016P015P044nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S4S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S5S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S6S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S7S102P016P015N044P032: std_logic_vector(   0 downto 0);
        signal cVar1S8S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S11S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S12S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S14S102P016P015P043P017: std_logic_vector(   0 downto 0);
        signal cVar1S15S102P016P015P043P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S102P016P015P043N005: std_logic_vector(   0 downto 0);
        signal cVar1S17S102P016P021P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S102P016P021P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S19S102P016P021P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S20S102P016P021P012P056: std_logic_vector(   0 downto 0);
        signal cVar1S21S102P016P021P012P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S102P016P021P012N040: std_logic_vector(   0 downto 0);
        signal cVar1S23S102P016P021P012N040: std_logic_vector(   0 downto 0);
        signal cVar1S24S102P016P021P012N040: std_logic_vector(   0 downto 0);
        signal cVar1S25S102P016P021P069P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S102P016P021P069N038: std_logic_vector(   0 downto 0);
        signal cVar1S27S102P016P021P069N038: std_logic_vector(   0 downto 0);
        signal cVar1S0S103P015P017P063P034: std_logic_vector(   0 downto 0);
        signal cVar1S1S103P015P017P063P034: std_logic_vector(   0 downto 0);
        signal cVar1S2S103P015P017P063P034: std_logic_vector(   0 downto 0);
        signal cVar1S3S103P015P017P063P034: std_logic_vector(   0 downto 0);
        signal cVar1S4S103P015P017P063P034: std_logic_vector(   0 downto 0);
        signal cVar1S5S103P015P017P063P035: std_logic_vector(   0 downto 0);
        signal cVar1S6S103P015P017P063N035: std_logic_vector(   0 downto 0);
        signal cVar1S7S103P015P017P063N035: std_logic_vector(   0 downto 0);
        signal cVar1S8S103P015P017P063N035: std_logic_vector(   0 downto 0);
        signal cVar1S9S103P015P017P035P014: std_logic_vector(   0 downto 0);
        signal cVar1S10S103P015P017P035N014: std_logic_vector(   0 downto 0);
        signal cVar1S11S103P015P017P035N014: std_logic_vector(   0 downto 0);
        signal cVar1S12S103P015P017P035N014: std_logic_vector(   0 downto 0);
        signal cVar1S13S103P015P017P035P065: std_logic_vector(   0 downto 0);
        signal cVar1S14S103N015P044P004P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S103N015P044P004N023: std_logic_vector(   0 downto 0);
        signal cVar1S16S103N015P044N004P007: std_logic_vector(   0 downto 0);
        signal cVar1S17S103N015P044N004P007: std_logic_vector(   0 downto 0);
        signal cVar1S18S103N015P044N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S19S103N015P044N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S20S103N015P044N004N007: std_logic_vector(   0 downto 0);
        signal cVar1S21S103N015N044P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S22S103N015N044P031P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S103N015N044P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S24S103N015N044P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S25S103N015N044P031N013: std_logic_vector(   0 downto 0);
        signal cVar1S26S103N015N044N031P030: std_logic_vector(   0 downto 0);
        signal cVar1S27S103N015N044N031P030: std_logic_vector(   0 downto 0);
        signal cVar1S28S103N015N044N031P030: std_logic_vector(   0 downto 0);
        signal cVar1S29S103N015N044N031P030: std_logic_vector(   0 downto 0);
        signal cVar1S30S103N015N044N031N030: std_logic_vector(   0 downto 0);
        signal cVar1S31S103N015N044N031N030: std_logic_vector(   0 downto 0);
        signal cVar1S32S103N015N044N031N030: std_logic_vector(   0 downto 0);
        signal cVar1S0S104P015P005P060P028: std_logic_vector(   0 downto 0);
        signal cVar1S1S104P015P005P060P028: std_logic_vector(   0 downto 0);
        signal cVar1S2S104P015P005P060P028: std_logic_vector(   0 downto 0);
        signal cVar1S3S104P015P005P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S104P015N005P063P052: std_logic_vector(   0 downto 0);
        signal cVar1S5S104P015N005P063N052: std_logic_vector(   0 downto 0);
        signal cVar1S6S104P015N005P063N052: std_logic_vector(   0 downto 0);
        signal cVar1S7S104P015N005P063N052: std_logic_vector(   0 downto 0);
        signal cVar1S8S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S11S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S12S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S14S104P015N005N063P017: std_logic_vector(   0 downto 0);
        signal cVar1S15S104P015P029P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S104P015P029P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S104P015P029P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S104P015N029P056P009: std_logic_vector(   0 downto 0);
        signal cVar1S19S104P015N029P056P009: std_logic_vector(   0 downto 0);
        signal cVar1S20S104P015N029P056P009: std_logic_vector(   0 downto 0);
        signal cVar1S21S104P015N029P056P009: std_logic_vector(   0 downto 0);
        signal cVar1S22S104P015N029P056P009: std_logic_vector(   0 downto 0);
        signal cVar1S23S104P015N029P056P031: std_logic_vector(   0 downto 0);
        signal cVar1S24S104P015N029P056N031: std_logic_vector(   0 downto 0);
        signal cVar1S25S104P015N029P056N031: std_logic_vector(   0 downto 0);
        signal cVar1S26S104P015N029P056N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S105P017P015P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S1S105P017P015P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S105P017P015P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S105P017P015P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S105P017P015P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S105P017P015P018P060nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S105P017P015P018N060: std_logic_vector(   0 downto 0);
        signal cVar1S7S105P017P015P018N060: std_logic_vector(   0 downto 0);
        signal cVar1S8S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S11S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S12S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S13S105P017P015P058P048: std_logic_vector(   0 downto 0);
        signal cVar1S14S105P017P015P058P035: std_logic_vector(   0 downto 0);
        signal cVar1S15S105P017P015P058P035: std_logic_vector(   0 downto 0);
        signal cVar1S16S105N017P015P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S105N017P015P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S18S105N017P015P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S19S105N017P015P034N014: std_logic_vector(   0 downto 0);
        signal cVar1S20S105N017P015P034N014: std_logic_vector(   0 downto 0);
        signal cVar1S21S105N017P015P034N014: std_logic_vector(   0 downto 0);
        signal cVar1S22S105N017P015P034N014: std_logic_vector(   0 downto 0);
        signal cVar1S23S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S24S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S25S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S26S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S27S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S28S105N017P015N034P065: std_logic_vector(   0 downto 0);
        signal cVar1S29S105N017P015P005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S30S105N017P015P005N004: std_logic_vector(   0 downto 0);
        signal cVar1S31S105N017P015P005N004: std_logic_vector(   0 downto 0);
        signal cVar1S32S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S33S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S34S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S35S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S36S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S37S105N017P015N005P043: std_logic_vector(   0 downto 0);
        signal cVar1S0S106P065P015P045P022: std_logic_vector(   0 downto 0);
        signal cVar1S1S106P065P015P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S2S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S3S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S4S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S5S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S6S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S7S106P065P015N045P043: std_logic_vector(   0 downto 0);
        signal cVar1S8S106P065P015P029P060: std_logic_vector(   0 downto 0);
        signal cVar1S9S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S10S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S11S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S12S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S106P065P015N029P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S106P065P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S106P065N052P035P017: std_logic_vector(   0 downto 0);
        signal cVar1S17S106P065N052P035P017: std_logic_vector(   0 downto 0);
        signal cVar1S18S106P065N052P035P017: std_logic_vector(   0 downto 0);
        signal cVar1S19S106P065N052P035N017: std_logic_vector(   0 downto 0);
        signal cVar1S20S106P065N052P035N017: std_logic_vector(   0 downto 0);
        signal cVar1S21S106P065N052P035N017: std_logic_vector(   0 downto 0);
        signal cVar1S22S106P065N052N035P034: std_logic_vector(   0 downto 0);
        signal cVar1S23S106P065N052N035P034: std_logic_vector(   0 downto 0);
        signal cVar1S24S106P065N052N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S25S106P065N052N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S26S106P065N052N035N034: std_logic_vector(   0 downto 0);
        signal cVar1S0S107P052P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S107P052N065P010P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S107P052N065P010P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S107P052N065N010P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S107P052N065N010P067: std_logic_vector(   0 downto 0);
        signal cVar1S5S107P052N065N010N067: std_logic_vector(   0 downto 0);
        signal cVar1S6S107P052N065N010N067: std_logic_vector(   0 downto 0);
        signal cVar1S7S107P052N065N010N067: std_logic_vector(   0 downto 0);
        signal cVar1S8S107P052N065N010N067: std_logic_vector(   0 downto 0);
        signal cVar1S9S107N052P044P025P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S107N052P044P025N005: std_logic_vector(   0 downto 0);
        signal cVar1S11S107N052P044P025N005: std_logic_vector(   0 downto 0);
        signal cVar1S12S107N052P044N025P067nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S107N052P044N025N067: std_logic_vector(   0 downto 0);
        signal cVar1S14S107N052P044N025N067: std_logic_vector(   0 downto 0);
        signal cVar1S15S107N052P044N025N067: std_logic_vector(   0 downto 0);
        signal cVar1S16S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S17S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S18S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S19S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S20S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S21S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S22S107N052N044P058P033: std_logic_vector(   0 downto 0);
        signal cVar1S23S107N052N044P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S24S107N052N044P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S25S107N052N044P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S26S107N052N044P058N033: std_logic_vector(   0 downto 0);
        signal cVar1S0S108P058P033P060P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S108P058P033P060P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S108P058P033P060P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S108P058P033P060N006: std_logic_vector(   0 downto 0);
        signal cVar1S4S108P058P033P060N006: std_logic_vector(   0 downto 0);
        signal cVar1S5S108P058P033P060N006: std_logic_vector(   0 downto 0);
        signal cVar1S6S108P058P033P060P066: std_logic_vector(   0 downto 0);
        signal cVar1S7S108P058P033P060P066: std_logic_vector(   0 downto 0);
        signal cVar1S8S108P058P033P060N066: std_logic_vector(   0 downto 0);
        signal cVar1S9S108P058P033P060N066: std_logic_vector(   0 downto 0);
        signal cVar1S10S108P058P033P060N066: std_logic_vector(   0 downto 0);
        signal cVar1S11S108P058P033P006P051: std_logic_vector(   0 downto 0);
        signal cVar1S12S108P058P033P006P051: std_logic_vector(   0 downto 0);
        signal cVar1S13S108P058P033P006P051: std_logic_vector(   0 downto 0);
        signal cVar1S14S108P058P033P006P017: std_logic_vector(   0 downto 0);
        signal cVar1S15S108P058P006P013P033: std_logic_vector(   0 downto 0);
        signal cVar1S16S108P058P006P013P033: std_logic_vector(   0 downto 0);
        signal cVar1S17S108P058P006P013N033: std_logic_vector(   0 downto 0);
        signal cVar1S18S108P058P006P013N033: std_logic_vector(   0 downto 0);
        signal cVar1S19S108P058P006P013N033: std_logic_vector(   0 downto 0);
        signal cVar1S20S108P058P006N013P014: std_logic_vector(   0 downto 0);
        signal cVar1S21S108P058P006N013P014: std_logic_vector(   0 downto 0);
        signal cVar1S22S108P058P006N013N014: std_logic_vector(   0 downto 0);
        signal cVar1S23S108P058P006N013N014: std_logic_vector(   0 downto 0);
        signal cVar1S24S108P058P006N013N014: std_logic_vector(   0 downto 0);
        signal cVar1S25S108P058P006P017nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S109P045P004P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S109P045N004P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S109P045N004P006N024: std_logic_vector(   0 downto 0);
        signal cVar1S3S109P045N004N006P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S109P045N004N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S5S109P045N004N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S6S109P045N004N006N023: std_logic_vector(   0 downto 0);
        signal cVar1S7S109N045P029P011P054: std_logic_vector(   0 downto 0);
        signal cVar1S8S109N045P029P011P054: std_logic_vector(   0 downto 0);
        signal cVar1S9S109N045P029P011N054: std_logic_vector(   0 downto 0);
        signal cVar1S10S109N045P029P011N054: std_logic_vector(   0 downto 0);
        signal cVar1S11S109N045P029P011N054: std_logic_vector(   0 downto 0);
        signal cVar1S12S109N045P029N011P010: std_logic_vector(   0 downto 0);
        signal cVar1S13S109N045P029N011P010: std_logic_vector(   0 downto 0);
        signal cVar1S14S109N045P029N011N010: std_logic_vector(   0 downto 0);
        signal cVar1S15S109N045P029N011N010: std_logic_vector(   0 downto 0);
        signal cVar1S16S109N045P029N011N010: std_logic_vector(   0 downto 0);
        signal cVar1S17S109N045N029P011P007: std_logic_vector(   0 downto 0);
        signal cVar1S18S109N045N029P011P007: std_logic_vector(   0 downto 0);
        signal cVar1S19S109N045N029P011P007: std_logic_vector(   0 downto 0);
        signal cVar1S20S109N045N029P011N007: std_logic_vector(   0 downto 0);
        signal cVar1S21S109N045N029P011N007: std_logic_vector(   0 downto 0);
        signal cVar1S22S109N045N029P011N007: std_logic_vector(   0 downto 0);
        signal cVar1S23S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S24S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S25S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S26S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S27S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S28S109N045N029P011P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S110P011P029P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S1S110P011P029P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S2S110P011P029P007P025: std_logic_vector(   0 downto 0);
        signal cVar1S3S110P011P029P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S110P011P029P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S5S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S6S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S7S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S8S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S9S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S10S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S11S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S12S110P011P029N007P049: std_logic_vector(   0 downto 0);
        signal cVar1S13S110P011P029P005P010: std_logic_vector(   0 downto 0);
        signal cVar1S14S110P011P029P005P010: std_logic_vector(   0 downto 0);
        signal cVar1S15S110P011P029P005N010: std_logic_vector(   0 downto 0);
        signal cVar1S16S110P011P029P005N010: std_logic_vector(   0 downto 0);
        signal cVar1S17S110P011P029P005N010: std_logic_vector(   0 downto 0);
        signal cVar1S18S110P011P029P054P057: std_logic_vector(   0 downto 0);
        signal cVar1S19S110P011P029P054P057: std_logic_vector(   0 downto 0);
        signal cVar1S20S110P011P029N054P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S110P011P029N054N053: std_logic_vector(   0 downto 0);
        signal cVar1S22S110P011P029N054N053: std_logic_vector(   0 downto 0);
        signal cVar1S23S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S24S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S25S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S26S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S27S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S28S110P011N029P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S29S110P011N029P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S30S110P011N029P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S31S110P011N029P069N068: std_logic_vector(   0 downto 0);
        signal cVar1S32S110P011N029P069N068: std_logic_vector(   0 downto 0);
        signal cVar1S0S111P009P049P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S111P009P049N025P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S111P009N049P053P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S111P009N049P053N029: std_logic_vector(   0 downto 0);
        signal cVar1S4S111P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S5S111P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S6S111P009N049N053P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S111P009N049N053N050: std_logic_vector(   0 downto 0);
        signal cVar1S8S111P009N049N053N050: std_logic_vector(   0 downto 0);
        signal cVar1S9S111N009P044P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S111N009P044N004P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S111N009P044N004N051: std_logic_vector(   0 downto 0);
        signal cVar1S12S111N009P044N004N051: std_logic_vector(   0 downto 0);
        signal cVar1S13S111N009P044N004N051: std_logic_vector(   0 downto 0);
        signal cVar1S14S111N009N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S111N009N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S111N009N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S17S111N009N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S18S111N009N044P042P058nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S111N009N044P042N058: std_logic_vector(   0 downto 0);
        signal cVar1S20S111N009N044P042N058: std_logic_vector(   0 downto 0);
        signal cVar1S0S112P009P049P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S112P009P049N025P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S112P009N049P050P027: std_logic_vector(   0 downto 0);
        signal cVar1S3S112P009N049P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S4S112P009N049P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S112P009N049P050N027: std_logic_vector(   0 downto 0);
        signal cVar1S6S112P009N049N050P053: std_logic_vector(   0 downto 0);
        signal cVar1S7S112P009N049N050P053: std_logic_vector(   0 downto 0);
        signal cVar1S8S112P009N049N050P053: std_logic_vector(   0 downto 0);
        signal cVar1S9S112P009N049N050N053: std_logic_vector(   0 downto 0);
        signal cVar1S10S112P009N049N050N053: std_logic_vector(   0 downto 0);
        signal cVar1S11S112N009P011P053P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S112N009P011P053P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S112N009P011P053P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S112N009P011P053N064: std_logic_vector(   0 downto 0);
        signal cVar1S15S112N009P011P053N064: std_logic_vector(   0 downto 0);
        signal cVar1S16S112N009P011P053P036: std_logic_vector(   0 downto 0);
        signal cVar1S17S112N009P011P053P036: std_logic_vector(   0 downto 0);
        signal cVar1S18S112N009P011P053P036: std_logic_vector(   0 downto 0);
        signal cVar1S19S112N009P011P053P036: std_logic_vector(   0 downto 0);
        signal cVar1S20S112N009P011P029P054: std_logic_vector(   0 downto 0);
        signal cVar1S21S112N009P011P029P054: std_logic_vector(   0 downto 0);
        signal cVar1S22S112N009P011P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S23S112N009P011P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S24S112N009P011P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S25S112N009P011N029P047: std_logic_vector(   0 downto 0);
        signal cVar1S26S112N009P011N029P047: std_logic_vector(   0 downto 0);
        signal cVar1S27S112N009P011N029P047: std_logic_vector(   0 downto 0);
        signal cVar1S28S112N009P011N029N047: std_logic_vector(   0 downto 0);
        signal cVar1S29S112N009P011N029N047: std_logic_vector(   0 downto 0);
        signal cVar1S30S112N009P011N029N047: std_logic_vector(   0 downto 0);
        signal cVar1S0S113P037P066P027P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S113P037P066P027N047: std_logic_vector(   0 downto 0);
        signal cVar1S2S113P037P066P027N047: std_logic_vector(   0 downto 0);
        signal cVar1S3S113P037P066P027P068: std_logic_vector(   0 downto 0);
        signal cVar1S4S113P037N066P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S5S113P037N066P069P068: std_logic_vector(   0 downto 0);
        signal cVar1S6S113P037N066N069P035: std_logic_vector(   0 downto 0);
        signal cVar1S7S113P037N066N069P035: std_logic_vector(   0 downto 0);
        signal cVar1S8S113P037N066N069N035: std_logic_vector(   0 downto 0);
        signal cVar1S9S113P037N066N069N035: std_logic_vector(   0 downto 0);
        signal cVar1S10S113P037N066N069N035: std_logic_vector(   0 downto 0);
        signal cVar1S11S113N037P059P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S113N037P059N043P058: std_logic_vector(   0 downto 0);
        signal cVar1S13S113N037P059N043P058: std_logic_vector(   0 downto 0);
        signal cVar1S14S113N037P059N043P058: std_logic_vector(   0 downto 0);
        signal cVar1S15S113N037N059P009P049: std_logic_vector(   0 downto 0);
        signal cVar1S16S113N037N059P009P049: std_logic_vector(   0 downto 0);
        signal cVar1S17S113N037N059P009P049: std_logic_vector(   0 downto 0);
        signal cVar1S18S113N037N059P009N049: std_logic_vector(   0 downto 0);
        signal cVar1S19S113N037N059P009N049: std_logic_vector(   0 downto 0);
        signal cVar1S20S113N037N059P009N049: std_logic_vector(   0 downto 0);
        signal cVar1S21S113N037N059P009N049: std_logic_vector(   0 downto 0);
        signal cVar1S22S113N037N059N009P054: std_logic_vector(   0 downto 0);
        signal cVar1S23S113N037N059N009P054: std_logic_vector(   0 downto 0);
        signal cVar1S24S113N037N059N009P054: std_logic_vector(   0 downto 0);
        signal cVar1S25S113N037N059N009P054: std_logic_vector(   0 downto 0);
        signal cVar1S26S113N037N059N009N054: std_logic_vector(   0 downto 0);
        signal cVar1S27S113N037N059N009N054: std_logic_vector(   0 downto 0);
        signal cVar1S28S113N037N059N009N054: std_logic_vector(   0 downto 0);
        signal cVar1S0S114P064P037P005P043: std_logic_vector(   0 downto 0);
        signal cVar1S1S114P064P037P005N043: std_logic_vector(   0 downto 0);
        signal cVar1S2S114P064P037P005N043: std_logic_vector(   0 downto 0);
        signal cVar1S3S114P064P037P005N043: std_logic_vector(   0 downto 0);
        signal cVar1S4S114P064P037N005P028: std_logic_vector(   0 downto 0);
        signal cVar1S5S114P064P037N005P028: std_logic_vector(   0 downto 0);
        signal cVar1S6S114P064P037N005P028: std_logic_vector(   0 downto 0);
        signal cVar1S7S114P064P037N005P028: std_logic_vector(   0 downto 0);
        signal cVar1S8S114P064P037N005N028: std_logic_vector(   0 downto 0);
        signal cVar1S9S114P064P037N005N028: std_logic_vector(   0 downto 0);
        signal cVar1S10S114P064P037N005N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S114P064P037N005N028: std_logic_vector(   0 downto 0);
        signal cVar1S12S114P064P037P061P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S114P064P037P061P012: std_logic_vector(   0 downto 0);
        signal cVar1S14S114P064P037P061P012: std_logic_vector(   0 downto 0);
        signal cVar1S15S114P064P037P061P012: std_logic_vector(   0 downto 0);
        signal cVar1S16S114P064P037P061N012: std_logic_vector(   0 downto 0);
        signal cVar1S17S114P064P037P061N012: std_logic_vector(   0 downto 0);
        signal cVar1S18S114P064P037P061P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S114P064P037P061N062: std_logic_vector(   0 downto 0);
        signal cVar1S20S114P064P037P061N062: std_logic_vector(   0 downto 0);
        signal cVar1S21S114P064P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S22S114P064N046P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S114P064N046N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S24S114P064N046N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S25S114P064N046N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S26S114P064N046N042P003: std_logic_vector(   0 downto 0);
        signal cVar1S0S115P049P026P033P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S115P049P026P033N007: std_logic_vector(   0 downto 0);
        signal cVar1S2S115P049P026P033N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S115P049N026P024P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S115P049N026P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S115P049N026P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S115P049N026P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S115P049N026N024P027: std_logic_vector(   0 downto 0);
        signal cVar1S8S115P049N026N024P027: std_logic_vector(   0 downto 0);
        signal cVar1S9S115P049N026N024P027: std_logic_vector(   0 downto 0);
        signal cVar1S10S115P049N026N024N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S115P049N026N024N027: std_logic_vector(   0 downto 0);
        signal cVar1S12S115P049N026N024N027: std_logic_vector(   0 downto 0);
        signal cVar1S13S115N049P064P050P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S115N049P064P050N065: std_logic_vector(   0 downto 0);
        signal cVar1S15S115N049P064P050N065: std_logic_vector(   0 downto 0);
        signal cVar1S16S115N049P064N050P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S115N049P064N050P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S115N049P064N050P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S115N049P064N050P008: std_logic_vector(   0 downto 0);
        signal cVar1S20S115N049P064N050P008: std_logic_vector(   0 downto 0);
        signal cVar1S21S115N049N064P047P028: std_logic_vector(   0 downto 0);
        signal cVar1S22S115N049N064P047P028: std_logic_vector(   0 downto 0);
        signal cVar1S23S115N049N064P047P028: std_logic_vector(   0 downto 0);
        signal cVar1S24S115N049N064P047N028: std_logic_vector(   0 downto 0);
        signal cVar1S25S115N049N064P047N028: std_logic_vector(   0 downto 0);
        signal cVar1S26S115N049N064P047N028: std_logic_vector(   0 downto 0);
        signal cVar1S27S115N049N064P047P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S28S115N049N064P047N069: std_logic_vector(   0 downto 0);
        signal cVar1S29S115N049N064P047N069: std_logic_vector(   0 downto 0);
        signal cVar1S30S115N049N064P047N069: std_logic_vector(   0 downto 0);
        signal cVar1S0S116P060P062P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S1S116P060P062P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S116P060P062P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S116P060P062P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S4S116P060P062P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S5S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S6S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S7S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S8S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S9S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S10S116P060P062N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S11S116P060P062P050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S116P060P062N050P068: std_logic_vector(   0 downto 0);
        signal cVar1S13S116P060P062N050P068: std_logic_vector(   0 downto 0);
        signal cVar1S14S116P060P062N050P068: std_logic_vector(   0 downto 0);
        signal cVar1S15S116P060P062N050P068: std_logic_vector(   0 downto 0);
        signal cVar1S16S116P060P062N050P068: std_logic_vector(   0 downto 0);
        signal cVar1S17S116P060P014P008P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S116P060P014P008N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S116P060P014P008N032: std_logic_vector(   0 downto 0);
        signal cVar1S20S116P060N014P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S21S116P060N014P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S22S116P060N014P033P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S116P060N014P033N013: std_logic_vector(   0 downto 0);
        signal cVar1S24S116P060N014P033N013: std_logic_vector(   0 downto 0);
        signal cVar1S25S116P060N014P033N013: std_logic_vector(   0 downto 0);
        signal cVar1S26S116P060N014N033P066: std_logic_vector(   0 downto 0);
        signal cVar1S27S116P060N014N033P066: std_logic_vector(   0 downto 0);
        signal cVar1S28S116P060N014N033N066: std_logic_vector(   0 downto 0);
        signal cVar1S29S116P060N014N033N066: std_logic_vector(   0 downto 0);
        signal cVar1S30S116P060N014N033N066: std_logic_vector(   0 downto 0);
        signal cVar1S31S116P060N014N033N066: std_logic_vector(   0 downto 0);
        signal cVar1S0S117P049P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S117P049N005P026P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S117P049N005N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S117P049N005N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S117P049N005N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S5S117P049N005N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S117P049N005N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S7S117P049N005N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S8S117N049P024P053P028: std_logic_vector(   0 downto 0);
        signal cVar1S9S117N049P024P053P028: std_logic_vector(   0 downto 0);
        signal cVar1S10S117N049P024P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S117N049P024P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S12S117N049P024P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S13S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S14S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S15S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S16S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S17S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S18S117N049P024N053P051: std_logic_vector(   0 downto 0);
        signal cVar1S19S117N049P024P026P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S117N049P024P026N002: std_logic_vector(   0 downto 0);
        signal cVar1S0S118P049P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S118P049P006N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S118P049N006P007P019: std_logic_vector(   0 downto 0);
        signal cVar1S3S118P049N006P007P019: std_logic_vector(   0 downto 0);
        signal cVar1S4S118P049N006N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S5S118P049N006N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S118P049N006N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S7S118P049N006N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S8S118P049N006N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S9S118N049P052P024P042: std_logic_vector(   0 downto 0);
        signal cVar1S10S118N049P052P024P042: std_logic_vector(   0 downto 0);
        signal cVar1S11S118N049P052P024P042: std_logic_vector(   0 downto 0);
        signal cVar1S12S118N049P052P024N042: std_logic_vector(   0 downto 0);
        signal cVar1S13S118N049P052P024N042: std_logic_vector(   0 downto 0);
        signal cVar1S14S118N049P052P024N042: std_logic_vector(   0 downto 0);
        signal cVar1S15S118N049P052P024P068: std_logic_vector(   0 downto 0);
        signal cVar1S16S118N049P052P024P068: std_logic_vector(   0 downto 0);
        signal cVar1S17S118N049P052P024P068: std_logic_vector(   0 downto 0);
        signal cVar1S18S118N049P052P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S118N049P052N065P067: std_logic_vector(   0 downto 0);
        signal cVar1S20S118N049P052N065P067: std_logic_vector(   0 downto 0);
        signal cVar1S21S118N049P052N065N067: std_logic_vector(   0 downto 0);
        signal cVar1S22S118N049P052N065N067: std_logic_vector(   0 downto 0);
        signal cVar1S23S118N049P052N065N067: std_logic_vector(   0 downto 0);
        signal cVar1S0S119P049P006P007P018nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S119P049P006P007P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S119P049N006P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S119P049N006P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S119P049N006N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S5S119P049N006N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S119P049N006N007P009: std_logic_vector(   0 downto 0);
        signal cVar1S7S119P049N006N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S8S119P049N006N007N009: std_logic_vector(   0 downto 0);
        signal cVar1S9S119N049P042P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S119N049P042N051P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S119N049P042N051P050: std_logic_vector(   0 downto 0);
        signal cVar1S12S119N049P042N051P050: std_logic_vector(   0 downto 0);
        signal cVar1S13S119N049N042P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S119N049N042P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S15S119N049N042P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S16S119N049N042P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S17S119N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S18S119N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S119N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S119N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S120P049P024P010P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S120P049P024P010P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S120P049P024P010N006: std_logic_vector(   0 downto 0);
        signal cVar1S3S120P049N024P026P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S120P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S120P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S120P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S7S120P049N024N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S120P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S120P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S10S120P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S120N049P042P050P004: std_logic_vector(   0 downto 0);
        signal cVar1S12S120N049P042P050P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S120N049P042P050P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S120N049P042P050N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S120N049P042P050N004: std_logic_vector(   0 downto 0);
        signal cVar1S16S120N049P042P050N004: std_logic_vector(   0 downto 0);
        signal cVar1S17S120N049N042P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S120N049N042P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S19S120N049N042P045N022: std_logic_vector(   0 downto 0);
        signal cVar1S20S120N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S120N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S120N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S23S120N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S121P049P024P010P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S121P049P024P010N006: std_logic_vector(   0 downto 0);
        signal cVar1S2S121P049N024P026P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S121P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S121P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S121P049N024P026N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S121P049N024N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S121P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S8S121P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S121P049N024N026N027: std_logic_vector(   0 downto 0);
        signal cVar1S10S121N049P042P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S121N049P042N051P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S121N049N042P045P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S121N049N042P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S14S121N049N042P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S15S121N049N042P045N004: std_logic_vector(   0 downto 0);
        signal cVar1S16S121N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S17S121N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S18S121N049N042N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S122P045P027P024P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S122P045P027P024N013: std_logic_vector(   0 downto 0);
        signal cVar1S2S122P045P027P024N013: std_logic_vector(   0 downto 0);
        signal cVar1S3S122P045P027P024N013: std_logic_vector(   0 downto 0);
        signal cVar1S4S122P045P027N024P025: std_logic_vector(   0 downto 0);
        signal cVar1S5S122P045P027N024P025: std_logic_vector(   0 downto 0);
        signal cVar1S6S122P045P027N024N025: std_logic_vector(   0 downto 0);
        signal cVar1S7S122P045P027N024N025: std_logic_vector(   0 downto 0);
        signal cVar1S8S122P045P027N024N025: std_logic_vector(   0 downto 0);
        signal cVar1S9S122N045P049P024P026: std_logic_vector(   0 downto 0);
        signal cVar1S10S122N045P049P024P026: std_logic_vector(   0 downto 0);
        signal cVar1S11S122N045P049P024P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S122N045P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S13S122N045P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S14S122N045P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S15S122N045P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S16S122N045P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S17S122N045P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S18S122N045N049P047P042: std_logic_vector(   0 downto 0);
        signal cVar1S19S122N045N049P047P042: std_logic_vector(   0 downto 0);
        signal cVar1S20S122N045N049P047P042: std_logic_vector(   0 downto 0);
        signal cVar1S21S122N045N049P047N042: std_logic_vector(   0 downto 0);
        signal cVar1S22S122N045N049P047N042: std_logic_vector(   0 downto 0);
        signal cVar1S23S122N045N049P047N042: std_logic_vector(   0 downto 0);
        signal cVar1S24S122N045N049P047N042: std_logic_vector(   0 downto 0);
        signal cVar1S25S122N045N049P047P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S26S122N045N049P047N064: std_logic_vector(   0 downto 0);
        signal cVar1S27S122N045N049P047N064: std_logic_vector(   0 downto 0);
        signal cVar1S0S123P042P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S123P042N051P050P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S123P042N051P050N039: std_logic_vector(   0 downto 0);
        signal cVar1S3S123P042N051P050N039: std_logic_vector(   0 downto 0);
        signal cVar1S4S123P042N051P050N039: std_logic_vector(   0 downto 0);
        signal cVar1S5S123N042P049P024P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S123N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S123N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S8S123N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S9S123N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S10S123N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S11S123N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S123N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S13S123N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S123N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S15S123N042N049P045P007: std_logic_vector(   0 downto 0);
        signal cVar1S16S123N042N049P045P007: std_logic_vector(   0 downto 0);
        signal cVar1S17S123N042N049P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S18S123N042N049P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S19S123N042N049P045N007: std_logic_vector(   0 downto 0);
        signal cVar1S20S123N042N049N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S123N042N049N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S123N042N049N045P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S124P042P050P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S124P042P050N021P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S124P042P050N021N051: std_logic_vector(   0 downto 0);
        signal cVar1S3S124P042P050N021N051: std_logic_vector(   0 downto 0);
        signal cVar1S4S124P042P050N021N051: std_logic_vector(   0 downto 0);
        signal cVar1S5S124N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S6S124N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S7S124N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S124N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S9S124N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S10S124N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S11S124N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S12S124N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S13S124N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S14S124N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S15S124N042N045P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S16S124N042N045P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S17S124N042N045P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S18S124N042N045N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S19S124N042N045N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S20S124N042N045N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S21S124N042N045N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S22S124N042N045N049P047: std_logic_vector(   0 downto 0);
        signal cVar1S0S125P042P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S125N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S125N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S125N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S125N042P045P027N024psss: std_logic_vector(   0 downto 0);
        signal cVar1S5S125N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S6S125N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S7S125N042N045P049P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S125N042N045P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S9S125N042N045P049N024: std_logic_vector(   0 downto 0);
        signal cVar1S10S125N042N045N049P032: std_logic_vector(   0 downto 0);
        signal cVar1S11S125N042N045N049P032: std_logic_vector(   0 downto 0);
        signal cVar1S12S125N042N045N049N032: std_logic_vector(   0 downto 0);
        signal cVar1S13S125N042N045N049N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S126P042P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S126P042N051P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S126P042N051P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S3S126P042N051P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S4S126P042N051P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S5S126P042N051N023P000nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S126P042N051N023N000: std_logic_vector(   0 downto 0);
        signal cVar1S7S126P042N051N023N000: std_logic_vector(   0 downto 0);
        signal cVar1S8S126N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S126N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S126N042P045P027P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S126N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S12S126N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S13S126N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S14S126N042P045P027N024: std_logic_vector(   0 downto 0);
        signal cVar1S15S126N042N045P049P007: std_logic_vector(   0 downto 0);
        signal cVar1S16S126N042N045P049N007: std_logic_vector(   0 downto 0);
        signal cVar1S17S126N042N045P049N007: std_logic_vector(   0 downto 0);
        signal cVar1S18S126N042N045P049N007: std_logic_vector(   0 downto 0);
        signal cVar1S19S126N042N045P049N007: std_logic_vector(   0 downto 0);
        signal cVar1S20S126N042N045N049P059: std_logic_vector(   0 downto 0);
        signal cVar1S21S126N042N045N049P059: std_logic_vector(   0 downto 0);
        signal cVar1S22S126N042N045N049P059: std_logic_vector(   0 downto 0);
        signal cVar1S23S126N042N045N049P059: std_logic_vector(   0 downto 0);
        signal cVar1S24S126N042N045N049P059: std_logic_vector(   0 downto 0);
        signal cVar1S0S127P042P050P004P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S127P042P050P004N040: std_logic_vector(   0 downto 0);
        signal cVar1S2S127P042P050N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S127P042P050N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S4S127P042P050N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S5S127P042P050N004N005: std_logic_vector(   0 downto 0);
        signal cVar1S6S127N042P049P024P004nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S127N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S8S127N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S9S127N042P049P024N004: std_logic_vector(   0 downto 0);
        signal cVar1S10S127N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S11S127N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S127N042P049N024P026: std_logic_vector(   0 downto 0);
        signal cVar1S13S127N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S127N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S15S127N042P049N024N026: std_logic_vector(   0 downto 0);
        signal cVar1S16S127N042N049P045P024: std_logic_vector(   0 downto 0);
        signal cVar1S17S127N042N049P045P024: std_logic_vector(   0 downto 0);
        signal cVar1S18S127N042N049P045P024: std_logic_vector(   0 downto 0);
        signal cVar1S19S127N042N049P045N024: std_logic_vector(   0 downto 0);
        signal cVar1S20S127N042N049P045N024: std_logic_vector(   0 downto 0);
        signal cVar1S21S127N042N049P045N024: std_logic_vector(   0 downto 0);
        signal cVar1S22S127N042N049P045N024: std_logic_vector(   0 downto 0);
        signal cVar1S23S127N042N049N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S24S127N042N049N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S25S127N042N049N045P020: std_logic_vector(   0 downto 0);
        signal cVar1S26S127N042N049N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S27S127N042N049N045N020: std_logic_vector(   0 downto 0);
        signal cVar1S28S127N042N049N045N020: std_logic_vector(   0 downto 0);
        signal cVar2S3S0P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S0N029P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S0N029N061P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S0P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S0N060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S0N060N033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S0P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S0N063P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S0N063N030P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S0P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S0N027P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S0N027N051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S0P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S0N049P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S0N049N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S0P065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S0N065P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S0N065N043P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S1P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S1N056P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S1P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S1N030P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S1N030N035P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S1P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S1N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S1N026N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S1P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S1N027P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S1N027N054P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S1P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S1N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S1N027N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S1P035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S1N035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S1N035N037P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S1P054P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S1P054N056P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S1N054P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S1N054N042P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S2P013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S2P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S2N066P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S2P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S2P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S2N017P067P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S2P065P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S2P065N052P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S2P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S2P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S2N021P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S2N021N004P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S2P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S2N052P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S2N052N026P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S2P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S2N025P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S2P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S2P060N033P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S2N060psss: std_logic_vector(   0 downto 0);
        signal cVar2S0S3P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S3P013P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S3P013N037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S3P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S3P066P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S3N066P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S3P066P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S3N066P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S3P009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S3P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S3P015N066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S3P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S3P015P016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S3P017P037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S3P017N037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S3N017P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S3N017N016P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S3P036P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S3P036N055P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S3P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S3N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S3N023N022P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S3P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S3N060P051P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S3N060N051P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S4P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S4P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S4N025P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S4N025N024P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S4P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S4N026P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S4N026N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S4P059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S4P059P058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S4N059P063P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S4N059N063P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S4P056P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S4P056N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S4N056psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S5P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S5N024P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S5P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S5N023P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S5N023N000P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S5P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S5P066P064P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S5P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S5P031N013P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S5N031P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S5N031N030P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S5P061P032P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S5P061N032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S5N061P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S5N061N041P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S6P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S6N007P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S6P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S6N026P029P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S6N026N029P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S6P031P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S6N031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S6N031P013P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S6P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S6N040P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S6P012P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S6P012P037P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S6P012P063P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S6P058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S6N058P037P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S6P033P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S6P033P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S6P061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S6P061N059P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S6N061P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S6N061N040P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S7P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S7N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S7P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S7N029P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S7N029N010P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S7P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S7N026P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S7P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S7P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S7N006P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S7N006N007P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S7P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S7N013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S7P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S7P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S7P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S7N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S7P062P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S7P062P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S7N062P066P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S7N062N066P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S8P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S8P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S8N007P042P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S8N007P042P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S8P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S8N048P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S8N048N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S8P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S8N008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S8N008N010P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S8P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S8N029P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S8P028P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S8N028P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S8N028N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S8P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S8P022N043P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S8N022psss: std_logic_vector(   0 downto 0);
        signal cVar2S23S8P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S8P061P013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S8N061P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S8P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S8P065N034P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S8N065P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S9P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S9N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S9N008N009P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S9P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S9N027P057P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S9P010P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S9P025P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S9N025P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S9N025N047P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S9P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S9N027P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S9N027N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S9P038P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S9P038N021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S9N038P009P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S9N038P009P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S10P067P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S10P067N008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S10P067P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S10P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S10N027P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S10N027N025P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S10P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S10P022N043P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S10N022psss: std_logic_vector(   0 downto 0);
        signal cVar2S9S10P066P018P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S10P066P018P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S10N066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S10P068P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S10P068P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S10P068P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S10P016P012P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S10P003P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S10P003N035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S10P066P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S10P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S10P016N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S10P016P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S10P003P035P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S10P067P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S10P067N051P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S10P067P069P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S10P034P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S10P066P012P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S10P066P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S10N066P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S10N066N069P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S10P034P063P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S10N034P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S10N034N031P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S11P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S11N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S11N009N005P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S11P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S11N009P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S11N009N007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S11P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S11P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S11P006N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S11N006P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S11N006N026P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S11P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S11P026N008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S11N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S11P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S11P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S11N044P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S11N044N040P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S11P042P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S11N042P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S11N042N043P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S11P043P007P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S11P043P007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S11P043P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S11P043N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S12P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S12N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S12N009N005P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S12P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S12N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S12N024N026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S12P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S12P008N026P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S12N008psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S12P003P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S12P003P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S12P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S12P026P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S12P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S12P047N026P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S12N047P050P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S12P033P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S12P033N010P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S12P015P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S13P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S13P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S13P006N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S13N006P017P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S13N006P017P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S13P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S13N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S13P010P016P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S13P010P016psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S13N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S13N010N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S13P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S13P029N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S13N029P009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S13P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S13N000P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S13N000N020P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S13P032P066P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S13P032P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S13N032P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S13P055P030P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S13P055N030P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S13N055P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S13N055N022P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S14P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S14N009P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S14N009N007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S14P007P011P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S14P007P011P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S14P022P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S14P022N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S14N022P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S14N022N025P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S14P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S14N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S14N021N020P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S14P003P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S14P003P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S14P035P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S14P035P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S14N035P003P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S14P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S14N056P015P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S14P019P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S14P019N059P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S14P019P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S14P019N014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S14P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S14N028P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S14N028N008P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S14P055P029P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S14N055P048P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S15P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S15N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S15P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S15N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S15N007N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S15P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S15P042P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S15P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S15N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S15N006N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S15P052P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S15P052N050P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S15P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S15P006N024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S15N006P065P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S15P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S15N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S15N002N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S15P042P069P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S15P042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S15P042N064P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S15P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S15N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S15N022N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S15P049P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S15P049N025P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S16P024P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S16P024N006P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S16N024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S16P013P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S16P013N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S16P013psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S16P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S16P036P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S16P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S16N045P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S16N045N041P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S16P038P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S16P038N040P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S16N038P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S16N038P043P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S16P033P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S16P033P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S16P033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S16P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S16P013P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S16P013N065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S16P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S16P016P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S16P016N036P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S16N016P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S16P063P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S16P063P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S16P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S17P066P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S17P066N020P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S17P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S17N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S17N006N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S17P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S17P024P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S17N024P050P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S17N024N050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S17P013P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S17P013N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S17P013P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S17P010P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S17N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S17N010N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S17P021P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S17N021P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S17N021N000P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S17P052P009P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S17P052N009P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S17N052P009P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S17N052P009P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S18P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S18N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S18P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S18N023P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S18P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S18N023P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S18N023N004P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S18P042P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S18P042N050P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S18P042P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S18P042N040P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S18P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S18P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S18N024P037P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S18P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S19P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S19P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S19N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S19P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S19N023P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S19N023N047P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S19P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S19N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S19N005N004P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S19P009P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S19P009N027P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S19N009P008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S19N009N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S19P000P015P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S19P000N015P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S19P000P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S19P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S20P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S20N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S20N007N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S20P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S20N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S20N020N021P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S20P039P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S20P039P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S20P039P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S20P039N064P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S20P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S20P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S20N050P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S20P008P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S20P016P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S20P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S20P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S20N053P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S20P003P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S20N003P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S20N003N055P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S20P069P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S20P035P014P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S20P035N014P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S20P035P012P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S20P054P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S20N054P064P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S21P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S21P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S21N023P022P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S21N023N022P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S21P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S21N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S21N025N027P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S21P051P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S21P051N008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S21N051P055P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S21P015P014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S21N015P017P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S22P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S22N021P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S22P003P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S22N003P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S22N003N022P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S22P030P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S22P030N040P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S22P030P010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S22P030P031P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S22N030P032P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S22N030N032P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S22P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S22N020P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S22N020N064P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S22P018P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S22N018P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S23P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S23N022P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S23P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S23P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S23P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S23P010N028P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S23N010P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S23P029P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S23P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S23P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S23P008N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S23N008P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S23N008N038P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S23P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S23P035P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S23P029P063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S23N029P030P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S24P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S24N022P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S24P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S24P022P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S24N022P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S24P060P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S24P060P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S24P060P035P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S24P060N035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S24P063P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S24P063N014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S24P063P034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S24P001P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S24P056P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S24P056N013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S24N056P014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S24P010P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S25P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S25P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S25P065P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S25P065N022P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S25P016P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S25P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S25P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S25N057P060P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S25P065P019P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S25P065N019psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S25P065P059P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S25P062P017P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S25P062N017P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S25P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S25N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S25P064P037P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S25N064P037P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S25N064N037P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S25P016P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S25P016N054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S25P012P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S26P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S26N039P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S26P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S26N003P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S26P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S26N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S26N047N045P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S26P007P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S26P007N045P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S26P005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S26P005N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S26N005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S26N005N042P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S26P045P043P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S26P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S26P045N022P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S26P045P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S26P045P027P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S26P067P007P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S26P067P007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S26P067P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S26P018P062P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S26N018P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S26N018N069P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S26P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S26N019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S26P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S26P034P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S26P034N064P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S26P014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S26N014P063P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S27P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S27N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S27P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S27N039P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S27P034P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S27P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S27P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S27N045P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S27N045N044P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S27P068P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S27P068N007P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S27P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S27N045P068P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S27P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S27N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S27P042P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S27P042N004P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S27N042P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S27N042N007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S27P009P027P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S27P009N027P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S27N009P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S27N009N026P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S27P005P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S27P005P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S27P005N022P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S28P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S28N044P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S28P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S28N007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S28P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S28P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S28N005P003P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S28P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S28N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S28N005N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S28P025P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S28N025P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S28N025N054P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S28P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S28P021P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S28P021N039P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S28P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S28N058P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S29P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S29N044P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S29P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S29N045P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S29P025P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S29P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S29P021P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S29P021N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S29N021P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S29N021P066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S29P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S29N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S29N005N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S29P025P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S29N025psss: std_logic_vector(   0 downto 0);
        signal cVar2S19S29P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S29P020N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S29N020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S29N020N005P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S29P039P005P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S30P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S30N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S30N027N024P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S30P034P015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S30P034P015P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S30N034P032P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S30N034N032psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S30P030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S30N030psss: std_logic_vector(   0 downto 0);
        signal cVar2S10S30P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S30N003P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S30N003N029P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S30P054P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S30P054N024P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S30P054P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S30P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S30N033P062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S30P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S30N050P035P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S30P060P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S30P060N052P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S30P060P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S30P031P048P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S30P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S30P036P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S30P016P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S30P016N036P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S30N016P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S30P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S30P063P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S31P063P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S31P063P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S31P063P034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S31P064P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S31P064N050P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S31N064P015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S31P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S31P065P013P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S31P030P014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S31P030N014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S31P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S31N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S31P033P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S31P032P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S31N032P008P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S31N032N008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S31P012P016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S31P012P016P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S31N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S31N012N010P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S31P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S31P023N005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S31N023P005P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S31N023P005P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S32P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S32N020P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S32N020N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S32P016P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S32P016P012P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S32N016P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S32N016N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S32P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S32P016P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S32P016P062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S32P016N062P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S32P057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S32P057N017P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S32P057P013P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S32P057N013P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S32P065P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S32P065P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S32P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S32N006P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S32N006N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S32P033P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S32P033P018P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S32N033P035P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S32N033N035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S32P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S32P010P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S32P064P035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S32P064N035P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S32N064P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S32N064N007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S32P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S32P049P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S32N049P014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S32P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S33P034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S33P034P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S33N034P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S33N034N036P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S33P032P057P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S33P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S33P062P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S33P062N004P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S33P062P008P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S33P064P010P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S33N064P066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S33N064N066P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S33P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S33N012P014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S33P069P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S33N069P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S33P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S33N002P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S33N002N003P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S33P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S33N004P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S33P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S33N023P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S33N023N006P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S33P050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S33P050P014P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S33N050P065P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S33N050P065P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S33P066P056P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S33P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S33P066N012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S33P064P035P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S34P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S34N026P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S34P051P016P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S34P051P016P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S34N051P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S34N051N027P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S34P058P033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S34P058N033P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S34N058P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S34N058P060P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S34P063P017P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S34P063N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S34N063P037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S34N063N037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S34P010P011P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S34P010P011P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S34P010P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S34P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S34P016N034P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S34N016P065P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S34P054P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S34P054N052P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S34P054P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S34P058P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S34P069P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S34P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S34P005P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S35P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S35N031P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S35N031N033P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S35P012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S35P031P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S35P031N014P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S35P031P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S35P069P009P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S35P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S35N056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S35N056N057P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S35P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S35N057P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S35P013P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S35P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S35N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S35N047N043P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S35P025P047P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S35P025N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S35P057P052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S35P057P052P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S35P057P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S35P031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S35P031N054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S35N031P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S35N031N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S36P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S36N027P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S36P024P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S36N024P052P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S36P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S36P027P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S36P027N007P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S36P049P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S36N049P052P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S36N049N052P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S36P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S36P025N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S36N025P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S36N025N004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S36P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S36P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S36N014P067P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S36P036P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S36P036P014P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S36P036N014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S36P033P003P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S36P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S36P014P068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S37P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S37N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S37N006N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S37P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S37N060P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S37N060N007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S37P036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S37P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S37N023P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S37P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S37P006N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S37N006P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S37N006N021P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S37P026P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S37P026N049P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S37N026P024P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S37P007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S37P007N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S37N007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S37P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S38P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S38N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S38N009N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S38P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S38N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S38N007N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S38P037P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S38P037N030P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S38P037P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S38P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S38P045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S38P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S38P045N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S38P016P065P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S38P016N065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S38N016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S38N016P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S38P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S38N018P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S38N018N056P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S38P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S38N044P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S38N044N043P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S38P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S38P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S39P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S39N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S39N009N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S39P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S39N006P009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S39N006N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S39P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S39N030P024P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S39N030N024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S39P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S39N023P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S39P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S39P006N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S39N006P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S39N006N021P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S39P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S39P067N015P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S39N067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S39N067N065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S39P018P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S39P018P016P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S39N018P016P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S39P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S39P019N018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S40P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S40N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S40N009N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S40P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S40N058P024P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S40P059P019P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S40P059P019P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S40N059P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S40N059N060P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S40P035P034P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S40P035P034P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S40N035P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S40N035N011P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S40P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S40N055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S40N055N054P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S40P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S40P030N057P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S40N030P029P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S40P028P057P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S40P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S40N007P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S40P066P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S40P066P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S40P015P019P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S40P015P019P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S40P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S40P015N012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S41P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S41N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S41N009N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S41P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S41P050N027P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S41N050P005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S41P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S41P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S41N054P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S41P043P025P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S41P043P025P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S41P043P019P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S41P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S41N022P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S41N022N007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S41P004P061P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S41P004N061P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S41P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S41P065N014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S41P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S41P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S41P013N031P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S41N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S41N013N011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S41P035P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S41P035P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S41N035P024P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S42P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S42N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S42N009N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S42P062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S42N062P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S42N062N006P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S42P015P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S42P015N021P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S42P022P043P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S42P022N043P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S42N022P046P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S42N022P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S42P047P063P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S42P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S42N014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S42N014P017P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S42P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S42P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S42P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S42N046P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S42P042P023P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S42P042P066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S42P017P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S42N017P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S42N017N041P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S43P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S43N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S43N009N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S43P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S43P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S43N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S43N007N006P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S43P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S43N045P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S43P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S43P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S43P049P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S43P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S43N002P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S43P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S43N041P067P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S43P008P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S43P008N049P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S43N008P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S43P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S43N042P017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S43N042N017P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S44P067P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S44P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S44N008P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S44N008P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S44P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S44P047N006P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S44N047P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S44N047N051P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S44P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S44N005P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S44P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S44N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S44N006N007P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S44P012P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S44P012N048P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S44P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S44N044P015P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S44N044N015P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S45P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S45P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S45N033P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S45N033N002P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S45P026P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S45P026N018P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S45N026P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S45P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S45N007P009P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S45N007N009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S45P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S45N028P026P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S45N028N026P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S45P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S45P027N009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S45N027P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S45P023P005P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S45P023N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S45N023P043P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S45P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S45N033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S46P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S46N061P069P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S46P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S46P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S46N045P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S46N045P052P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S46P025P059P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S46P025P059P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S46P025P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S46P062P069P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S46P062N069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S46P005P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S46N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S46N005N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S46P043P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S46P043P045P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S46P043P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S46P043N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S47P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S47N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S47N004N005P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S47P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S47N061P067P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S47P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S47N043P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S47P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S47N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S47N007N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S47P025P050P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S47N025P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S47N025N045P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S47P045P037P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S47P045N037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S47P045P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S47P045N047P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S47P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S47P007N025P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S47N007P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S47N007N059P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S48P055P056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S48P055P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S48P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S48P023N005P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S48N023P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S48N023N028psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S48P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S48N062P059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S48N062N059P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S48P064P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S48P035P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S48N035P062P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S48P034P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S48P034N014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S48N034P035P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S48P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S48N015P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S48P066P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S48P066P018P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S48P066N018P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S48P018P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S48P018N062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S48P018P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S48P004P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S48P004N022P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S48N004P062P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S48P018P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S48P018N015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S48N018P032P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S48P029P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S48P029N017P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S49P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S49N043P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S49P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S49N054P004P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S49N054N004P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S49P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S49N019P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S49N019N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S49P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S49N007P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S49N007N002P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S49P034P063P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S49P034N063P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S49N034P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S49P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S49P010P055P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S49P010N055P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S49N010P029P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S49P059P032P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S49P059N032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S49N059P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S50P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S50N043P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S50P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S50N064P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S50P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S50P008P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S50N008P063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S50P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S50N007P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S50P024P006P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S50P024N006P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S50N024P045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S50N024P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S50P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S50N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S50P026P036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S50N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S50N026N027P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S51P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S51N053P055P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S51N053N055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S51P063P068P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S51P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S51P026P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S51P026N007psss: std_logic_vector(   0 downto 0);
        signal cVar2S10S51P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S51N046P003P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S51P006P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S51P006N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S51N006P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S51P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S51P041N020P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S51N041P039P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S52P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S52N006P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S52N006N007P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S52P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S52N024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S52P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S52N060P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S52N060N044P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S52P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S52P034P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S52P034N054P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S52P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S52N053P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S52N053N057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S52P029P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S52P029N008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S52P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S52N002P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S52P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S52N020P066P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S52P046P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S52P046P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S52N046P007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S52P015P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S52P015P056P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S52N015P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S52N015P005P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S53P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S53N006P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S53P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S53N057P037P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S53P005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S53P005N017P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S53P063P053P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S53P063N053P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S53P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S53P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S53N002P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S53P066P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S53P066N020P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S53P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S53N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S53N022N024P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S53P015P047P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S53P015P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S53N015P018P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S53N015N018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S54P003P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S54N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S54N003N005P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S54P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S54N023P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S54N023N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S54P036P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S54P036P009P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S54P028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S54N028P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S54N028N025P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S54P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S54N027P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S54N027N045P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S54P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S54P006P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S54N006P033P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S54P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S54N025P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S54P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S54N013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S54P007P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S54N007P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S55P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S55N003P005P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S55P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S55N004P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S55N004N050P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S55P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S55P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S55P013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S55P013N022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S55P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S55P006N024P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S55N006P007P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S55N006N007P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S55P042P032P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S55P042N032psss: std_logic_vector(   0 downto 0);
        signal cVar2S17S55P042P016P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S55P042N016P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S55P033P049P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S55P029P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S55P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S55P025P046P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S55P025N046P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S55N025P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S55N025N018P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S56P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S56N024P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S56P007P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S56N007P003P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S56N007N003P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S56P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S56P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S56N020P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S56P015P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S56P015P003P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S56P015P016P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S56P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S56N041P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S56N041N011P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S56P011P029P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S56P011P029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S56P011N029P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S56P026P035P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S56P026N035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S57P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S57N024P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S57P007P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S57N007P014P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S57N007N014P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S57P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S57N003P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S57N003N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S57P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S57P008P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S57P008N060P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S57P011P029P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S57P011P029P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S57P011P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S57P011N053P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S57P001P017P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S57P001N017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S57P008P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S57P008N049P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S57N008P021P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S57P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S57N041P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S58P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S58P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S58N004P007P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S58N004N007P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S58P038P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S58N038P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S58N038N062P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S58P021P038P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S58P021P038P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S58P021P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S58P021N003P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S58P041P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S58P041N005P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S58N041P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S58N041N011P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S58P035P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S58P035N065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S58N035P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S58N035N039P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S58P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S58N064P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S58P028P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S58N028P055P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S58P036P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S58P036N012P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S59P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S59P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S59N044P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S59N044N067P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S59P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S59N003P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S59N003N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S59P018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S59P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S59P046P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S59P046N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S59N046P003P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S59P022P057P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S59P022P057P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S59P030P031P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S59N030P057P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S59N030P057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S60P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S60N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S60N006N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S60P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S60N021P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S60N021N039P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S60P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S60N049P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S60N049N021P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S60P065P030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S60P065N030psss: std_logic_vector(   0 downto 0);
        signal cVar2S13S60P065P066P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S60P065P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S60P041P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S60P041N022P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S60N041P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S60P066P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S60P066N046P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S60P066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S60N066P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S60P066P006P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S60P066N006P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S60P066P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S61P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S61N013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S61P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S61N022P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S61N022N044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S61P017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S61N017P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S61N017N009P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S61P059P068P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S61P059N068psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S61P059P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S61P006P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S61N006P068P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S61P016P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S61N016P024P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S61P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S61N049P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S61P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S61P028N010P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S61N028P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S61P063P060P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S62P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S62N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S62N006N004P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S62P014P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S62P014N022P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S62N014P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S62N014N061P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S62P031P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S62P031N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S62P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S62P031N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S62N031P054P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S62N031P054P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S62P035P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S62P035N013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S62P014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S62P014N034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S62N014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S62P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S62N035P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S62P063P065P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S62P063N065P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S63P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S63P006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S63N006P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S63N006N004psss: std_logic_vector(   0 downto 0);
        signal cVar2S5S63P033P027P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S63P033N027psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S63P033P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S63P033N059P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S63P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S63N064P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S63N064N013P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S63P007P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S63P007N031P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S63P007P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S63P007N049P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S63P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S63P035P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S63P035P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S63P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S63N013P011P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S63N013N011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S63P057P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S63P057N014P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S63P057P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S63P057N028P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S64P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S64N053P054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S64N053N054P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S64P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S64N020P014P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S64N020N014P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S64P045P004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S64P045N004psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S64N045P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S64N045N041P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S64P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S64N009P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S64P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S64N065P017P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S64N065P017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S64P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S64P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S64N059P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S64P035P067P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S64P035P017P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S64P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S64N054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S64N054N057P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S64P057P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S64P057N037P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S64P013P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S64P013N043P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S64P013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S64P068P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S64P068P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S64P066P036P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S64P066N036P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S64N066P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S64N066P036P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S65P037P029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S65P037P024P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S65P012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S65N012P056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S65P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S65N005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S65P031P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S65P031N036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S65N031P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S65N031N032P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S65P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S65N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S65P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S65P009P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S65P009N021P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S65P004P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S65N004psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S65P011P029P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S65P011N029P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S65N011P020P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S65P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S66P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S66N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S66P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S66P009P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S66P009N021P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S66P009P027P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S66P009N027P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S66N009P027P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S66N009P027P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S66P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S66N011P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S66N011N007P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S66P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S66P041P036P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S66P041N036P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S66P017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S66P017P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S66N017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S66P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S66P057P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S66P057N012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S66P069P063P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S66P002P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S66P002N034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S66N002P038P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S67P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S67N019P052P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S67P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S67N025P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S67P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S67N001P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S67P012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S67P012N065P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S67N012P017P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S67P018P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S67P018N007P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S67P018P012P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S67P003P036P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S67P003P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S67P031P013P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S67P031N013P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S67N031P004P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S67N031P004P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S67P020P015P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S67P020N015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S67P020P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S67P020N019P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S67P011P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S68P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S68P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S68N025P019P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S68P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S68N029P051P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S68P015P064P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S68P015P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S68N015P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S68N015N034P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S68P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S68N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S68N002N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S68P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S68N038P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S68P018P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S68P018N007P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S68P018P012P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S68P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S68P054N013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S68N054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S68N054N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S68P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S68P020P039P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S68P020P050P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S68P035P053P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S68P035P029P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S68P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S68P018P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S68N018P069P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S69P013P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S69P013P051P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S69P013psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S69P051P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S69N051P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S69P027P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S69N027P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S69N027N029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S69P051P019P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S69P051N019P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S69P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S69N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S69N002N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S69P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S69P021P040P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S69N021P039P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S69P054P012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S69P054P012psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S69N054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S69N054N057P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S69P054P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S69N054P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S69P039P016P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S69P039N016P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S69P039P011P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S69P011P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S69P011N029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S69N011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S69N011N010P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S70P014P028P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S70P014N028psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S70P014P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S70P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S70P023N005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S70N023P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S70N023N049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S70P037P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S70P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S70P019P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S70P019N065P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S70N019P065P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S70P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S70P047P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S70P047P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S70P047N009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S70P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S70N049P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S70P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S70N040P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S70P042P047P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S70P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S70P042N005P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S70P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S70P036P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S70P036N015P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S70P010P009P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S71P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S71N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S71P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S71N021P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S71N021N022P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S71P039P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S71P039N067P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S71P039P017P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S71P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S71P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S71N006P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S71P027P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S71P027P048P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S71N027P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S71P007P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S71N007P004P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S71N007N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S71P047P016P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S71P047N016P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S71P047P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S71P047N069P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S71P011P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S71P011N020P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S72P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S72N043P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S72P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S72N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S72N006N008P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S72P028P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S72N028P031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S72N028N031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S72P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S72P047P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S72P047N028P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S72P047P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S72P047N009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S72P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S72N031P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S72N031N046P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S72P019P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S72P019P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S72P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S72N029P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S72N029P007P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S72P053P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S72P053P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S72P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S72N013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S72P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S72N007P018P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S72N007N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S72P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S73P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S73P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S73P009P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S73N009P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S73N009N005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S73P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S73P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S73P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S73N057P060P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S73N057N060P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S73P008P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S73P008N055P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S73P055P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S73P055N012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S73P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S73N056P057P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S73N056N057P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S73P010P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S73P010N057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S73N010P013P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S73P019P066P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S73P019N066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S73N019P068P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S73P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S73N032P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S73N032N028P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S74P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S74P017P015P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S74P017P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S74P017N052P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S74P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S74N007P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S74N007N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S74P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S74P020N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S74N020P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S74N020N005P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S74P029P011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S74P029N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S74N029P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S74N029N028P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S74P023P042P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S74P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S74P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S74P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S74N012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S74P029P009P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S74P029P009P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S74P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S74N010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S74P033P062P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S74P033N062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S74P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S74P016P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S75P050P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S75P050P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S75P008P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S75P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S75P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S75N050P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S75N050N053P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S75P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S75N015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S75P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S75N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S75N002N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S75P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S75N021P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S75N021N022P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S75P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S75N001P039P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S75P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S75N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S75N022N024P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S75P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S75N049P066P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S75P028P010P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S75N028P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S76P050P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S76N050P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S76P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S76P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S76N013P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S76P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S76N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S76N003N002P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S76P005P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S76N005P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S76N005N001P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S76P034P063P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S76P034N063P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S76N034P063P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S76N034P063P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S76P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S76N042P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S76P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S76N046P034P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S76N046P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S76P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S76P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S76N019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S77P057P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S77P057P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S77P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S77P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S77N067P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S77N067N003P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S77P039P016P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S77P039N016P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S77P039P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S77P015P052P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S77P015P018P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S77P015N018P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S77P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S77N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S77P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S77N039P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S77N039N043P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S77P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S77P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S77N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S77N009N008P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S77P023P042P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S77P023N042P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S77N023P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S77N023N013P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S77P003P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S77P003N052P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S77P003N034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S77P008P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S78P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S78N049P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S78P011P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S78P011P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S78P011P015P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S78P011N015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S78P011P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S78N011P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S78N011N015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S78P028P053P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S78P028N053P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S78N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S78N028N026P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S78P036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S78P036P034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S78P036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S78P064P006P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S78P064P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S78P036P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S78N036P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S78N036P065P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S78P064P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S78P064P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S78P064N068P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S78P064P059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S78P064P059P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S78N064P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S78N064N052P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S79P026P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S79N026P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S79P053P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S79P053N029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S79N053P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S79P011P053P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S79N011P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S79N011N007P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S79P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S79N002P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S79N002N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S79P021P005P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S79P021N005psss: std_logic_vector(   0 downto 0);
        signal cVar2S17S79N021P039P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S79P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S79N009P024P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S79P024P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S79P024N006psss: std_logic_vector(   0 downto 0);
        signal cVar2S22S79N024P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S79N024N027P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S79P032P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S79P032P011P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S79N032P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S79P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S79N034P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S79N034N033P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S80P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S80P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S80N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S80N023N022P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S80P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S80N000P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S80N000N050P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S80P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S80P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S80P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S80P055P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S80P053P064P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S80N053P002P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S80P029P011P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S80P029N011P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S80N029P062P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S80N029N062psss: std_logic_vector(   0 downto 0);
        signal cVar2S21S80P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S80N019P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S80P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S80N008P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S81P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S81N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S81N023N022P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S81P020P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S81P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S81P014P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S81P068P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S81P068P018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S81P054P057P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S81N054P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S81N054N053P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S81P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S81P010N052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S81N010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S81N010N009P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S81P025P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S81N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S81N025N027P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S81P062P026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S81P062P026P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S81N062P015P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S82P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S82P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S82P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S82P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S82P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S82P049N026P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S82N049P023P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S82N049N023P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S82P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S82P021N002P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S82N021P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S82P012P059P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S82P012N059P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S82N012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S82N012N014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S82P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S82P058P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S82P058P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S82N058P059P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S82P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S82N018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S82P055P027P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S82P055P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S82P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S83P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S83N043P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S83N043N042P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S83P066P027P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S83P066N027psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S83P066P019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S83P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S83N066P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S83P062P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S83P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S83P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S83N039P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S83N039N004P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S83P062P029P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S83P062N029P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S83P014P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S83N014P064P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S83P001P003P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S83P001P003P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S83P001P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S83P001N039P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S84P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S84N003P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S84N003N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S84P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S84N039P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S84N039N060P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S84P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S84P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S84N047P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S84N047N042P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S84P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S84P011P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S84P011N015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S84P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S84P003P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S84P003P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S84P003P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S84P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S84N039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S84N039N003P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S84P065P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S84N065P017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S84N065P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S84P029P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S84P029N051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S84N029P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S84N029N067P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S85P011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S85P011P012P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S85P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S85P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S85P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S85N010P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S85N010N037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S85P038P054P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S85P038P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S85P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S85N042P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S85N042N037P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S85P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S85P025P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S85N025P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S85N025N005P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S85P013P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S85P013N056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S85N013P057P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S85P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S85N049P043P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S86P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S86N003P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S86P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S86P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S86N002P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S86N002N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S86P013P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S86P013N066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S86N013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S86N013N003P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S86P014P055P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S86P014N055P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S86P014P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S86P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S86P005P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S86P005N049P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S86P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S86N019P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S86P006P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S86N006P055P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S87P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S87N067P019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S87N067P019P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S87P033P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S87P033N039P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S87P039P007P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S87P039N007psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S87P039P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S87P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S87N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S87P042P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S87P042N002P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S87N042P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S87N042N003P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S87P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S87P035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S87P035N013P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S87P055P026P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S87P055P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S87P055N069P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S87P030P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S87P030N010P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S87N030P011P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S87N030N011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S88P034P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S88P034N020P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S88P035P003P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S88P035N003psss: std_logic_vector(   0 downto 0);
        signal cVar2S4S88P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S88P035N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S88P053P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S88P053N010P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S88N053P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S88P036P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S88P036P012P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S88P031P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S88N031P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S88P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S88P068N019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S88N068P012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S88N068N012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S88P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S88N057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S88P033P007P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S88P024P005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S88P024N005psss: std_logic_vector(   0 downto 0);
        signal cVar2S25S88P039P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S88P039P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S89P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S89N033P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S89N033P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S89P012P033P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S89N012P032P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S89N012N032P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S89P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S89N063P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S89P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S89P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S89P005P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S89P005P019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S89N005P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S89N005N019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S89P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S89N058P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S89P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S89N002P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S89P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S89N021P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S89P017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S89P005P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S89N005P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S89N005N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S89P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S89N021P017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S89P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S89P027N009P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S89N027P042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S90P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S90P050P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S90P050N024P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S90P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S90N018P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S90N018N004P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S90P003P009P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S90P043P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S90N043P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S90N043N048P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S90P015P013P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S90P015P013P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S90N015P057P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S90N015P057P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S91P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S91P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S91N053P069P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S91P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S91P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S91N024P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S91P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S91N007P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S91N007N051P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S91P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S91N054P003P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S91P010P028P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S91P010N028P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S91N010P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S91P057P043P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S91P057P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S91P057N059P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S92P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S92N002P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S92P035P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S92P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S92P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S92P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S92N024P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S92P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S92N007P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S92N007N051P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S92P003P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S92P003N052P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S92P006P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S92N006P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S92N006N002P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S92P042P023P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S92P042P023P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S92P042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S92P042N064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S93P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S93P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S93N023P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S93P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S93N057P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S93N057N050P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S93P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S93N014P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S93N014N007P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S93P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S93P027P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S93P027N006P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S93P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S93N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S93N003N002P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S93P004P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S93P004N010P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S93P006P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S93N006P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S93N006N004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S93P042P004P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S93P042P004P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S93P042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S93P042N064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S94P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S94P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S94N023P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S94P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S94N042P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S94P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S94N005P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S94N005N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S94P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S94N051P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S94N051N002P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S94P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S94N039P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S94P045P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S94P045N006P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S94N045P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S94N045P004P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S94P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S94N069P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S95P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S95N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S95P006P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S95P006N022P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S95N006P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S95N006N060P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S95P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S95N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S95N023N022P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S95P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S95N000P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S95N000N039P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S95P023P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S95N023P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S95N023N006P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S95P039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S95P039N003P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S95N039P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S95N039N048P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S95P042P016P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S95P042N016P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S95P042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S95P042N064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S96P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S96P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S96P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S96P006N024P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S96N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S96N006N007P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S96P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S96N030P065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S96P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S96P067P065P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S96P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S96P067N034P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S96P028P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S96N028P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S96P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S96P030P031P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S96P047P053P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S96P047P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S96P047N066P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S96P062P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S96P062N060P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S96N062P058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S96P007P010P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S96P007N010P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S97P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S97P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S97N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S97P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S97N057P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S97N057N006P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S97P047P053P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S97P047P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S97P047N066P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S97P065P058P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S97P065P058P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S97P065P063P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S97P007P010P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S97P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S97N030P065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S97P032P014P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S97P032P014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S97N032P054P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S97P028P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S97P028N011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S97N028P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S97P032P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S97P032N041P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S97P032P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S98P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S98P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S98N021P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S98N021N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S98P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S98N030P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S98P041P032P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S98P041N032psss: std_logic_vector(   0 downto 0);
        signal cVar2S10S98P041P018P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S98P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S98P050P014P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S98P050P014P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S98P014P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S98P014N060P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S98N014P058P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S98P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S98P002P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S98P002N009P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S98N002P045P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S98P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S98N006P018P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S98N006N018P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S98P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S98P015N019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S99P004P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S99P004N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S99N004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S99N004N021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S99P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S99N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S99P066P035P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S99P066P035P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S99P066P058P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S99P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S99P008N026P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S99N008P047P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S99N008P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S99P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S99N023P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S99N023N039P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S99P056P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S99P056N060P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S99P056P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S99P056N031P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S99N056P011P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S99N056P011P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S99P033P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S99P033N066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S100P025P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S100N025P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S100N025N005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S100P034P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S100P034N039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S100P034P014P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S100P012P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S100P012N061P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S100P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S100P012N036P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S100P016P014P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S100P016P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S100N016P014P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S100N016N014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S100P012P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S100P012N057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S100P068P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S100P068P066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S100P068P066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S100P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S100P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S100P035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S100P035N037P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S100P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S100P024P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S100N024P031P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S100N024N031P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S101P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S101P021P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S101P066P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S101P066N067P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S101P066P017P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S101P066N017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S101P014P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S101P014N029P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S101P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S101N052P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S101N052N027P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S101P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S101P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S101P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S101P004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S101N004P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S101N004N021P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S101P019P047P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S101P019P047P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S101P019P010P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S101P019P010P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S101P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S101P056P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S101P056N030P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S101N056P032P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S101N056N032P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S101P002P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S101N002P032P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S102P031P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S102P031N056P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S102N031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S102N031P054P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S102P012P014P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S102P012P014P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S102N012P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S102P035P002P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S102N035P063P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S102N035P063P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S102P036P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S102P036P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S102N036P068P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S102N036N068P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S102P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S102P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S102N019P011P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S102P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S102N005P013P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S102P000P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S102P000N010P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S102N000P032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S102P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S102N008P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S103P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S103P036P011P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S103P036N011P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S103P059P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S103N059P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S103P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S103P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S103P069N014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S103N069P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S103P001P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S103P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S103P065N034P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S103P065P011P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S103P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S103P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S103P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S103N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S103P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S103N059P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S103N059P014P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S103P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S103N054P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S103P011P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S103P011N057P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S103N011P055P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S103P060P010P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S103P060N010P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S103P060P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S103P060N066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S103P057P010P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S103P057P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S103P057N060P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S104P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S104P065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S104P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S104P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S104P026P035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S104P026N035P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S104P026P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S104P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S104P013N031P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S104N013P061P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S104P008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S104P008N047P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S104N008P047P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S104N008P047P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S104P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S104P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S104P019N012P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S104P054P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S104N054P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S104N054P026P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S104P054P049P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S104P054N049P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S104P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S104P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S104N068P012P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S104N068N012P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S105P005P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S105N005psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S105P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S105N008P011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S105N008N011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S105P061P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S105P061N035P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S105P029P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S105P029N050P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S105N029P024P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S105N029N024P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S105P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S105N025P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S105P013P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S105N013P012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S105P066P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S105P066N059P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S105P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S105P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S105P016P036P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S105N016P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S105N016N035P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S105P062P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S105P062N039P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S105P062N064P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S105P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S105P067P063P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S105N067P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S105P012P069P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S105P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S105P014P048P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S33S105P014N048P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S34S105P014P009P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S35S105P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S36S105N016P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S37S105N016N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S106P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S106P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S106P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S106P052P008P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S106P052N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S106P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S106N022P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S106N022N049P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S106P036P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S106P055P012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S106N055P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S106N055P021P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S106P021P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S106N021P018P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S106N021P018P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S106P037P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S106P037P036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S106P037P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S106P015P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S106P015N067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S106N015P062P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S106P059P024P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S106P059P068P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S106P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S106N036P067P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S106N036N067P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S107P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S107N069P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S107P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S107N015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S107P009P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S107P009N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S107N009P008P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S107N009N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S107P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S107N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S107P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S107N054P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S107N054N023P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S107P006P047P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S107P006N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S107N006P060P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S107P006P035P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S107P013P010P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S107N013P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S107N013N012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S107P056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S107P056N012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S107N056P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S107N056N014P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S108P024P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S108P024P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S108N024psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S108P029P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S108P029N011P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S108N029psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S108P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S108N063P010P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S108P062P064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S108P062P064P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S108N062P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S108P069P066P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S108P069N066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S108P069P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S108P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S108P010P012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S108P010P012psss: std_logic_vector(   0 downto 0);
        signal cVar2S17S108P031P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S108N031P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S108N031N064P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S108P009P015P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S108P009P015P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S108P012P015P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S108P012P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S108N012P015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S109P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S109P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S109N050P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S109N050N007P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S109P057P050P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S109P057P050P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S109P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S109N053P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S109N053N055P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S109P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S109N052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S109P009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S109P009N050P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S109N009P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S109P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S109P025N046P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S109N025P028P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S109P047P009P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S109P047P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S109P047N006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S109P031P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S109P031N054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S109N031P013P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S109N031N013P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S109P037P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S109N037P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S110P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S110N046P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S110N046N047P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S110P028P009P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S110P028N009psss: std_logic_vector(   0 downto 0);
        signal cVar2S5S110P009P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S110P009P027P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S110P009P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S110P009N050P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S110P006P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S110P006N024P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S110N006P009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S110N006N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S110P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S110N052P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S110P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S110N009P013P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S110N009N013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S110P050P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S110P050P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S110P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S110N055P052P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S110P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S110P047N026P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S110N047P020P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S110N047N020P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S110P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S110N056P057P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S110P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S110N012P009P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S110P018P035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S32S110N018P014P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S111P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S111P003P063P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S111P027P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S111N027P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S111N027N029P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S111P007P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S111N007P027P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S111P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S111N021P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S111N021N011P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S111P068P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S111N068P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S111P004P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S111P004N043P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S111P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S111N023P021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S112P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S112P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S112P029P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S112N029P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S112N029N066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S112P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S112N029P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S112N029N035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S112P051P010P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S112P051P010P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S112P034P060P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S112P034P060P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S112P034P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S112P037P059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S112P037N059psss: std_logic_vector(   0 downto 0);
        signal cVar2S16S112P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S112N042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S112N042N005P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S112P019P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S112P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S112N017P014P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S112P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S112N053P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S112N053N055P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S112P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S112N026P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S112N026N066P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S112P020P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S112P020N041P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S112N020P039P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S113P048P042P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S113P048P017P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S113P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S113P060P064P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S113P060P064P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S113P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S113P062P064P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S113P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S113N021P018P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S113N021N018P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S113P000P055P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S113P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S113N067P060P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S113P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S113N025P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S113N025P019P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S113P057P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S113P057N028P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S113N057P027P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S113N057N027P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S113P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S113P010P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S113N010P011P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S113N010N011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S113P031P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S113P031N016P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S113P031P058P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S114P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S114P007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S114N007P069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S114N007P069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S114P053P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S114P053P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S114N053P012P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S114N053N012P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S114P029P054P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S114P029N054P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S114N029P026P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S114N029N026P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S114P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S114P013P016P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S114N013P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S114N013N056P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S114P068P000P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S114N068P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S114P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S114N069P016P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S114P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S114N036P011P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S114P007P036P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S114P007N036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S115P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S115N011P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S115P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S115N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S115N006N005P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S115P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S115P048P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S115P048P047P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S115P047P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S115P047N033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S115P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S115P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S115N018P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S115P005P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S115P005P059P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S115P005P019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S115P010P019P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S115P010N019P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S115P053P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S115N053P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S115N053N057P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S115P029P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S115N029P005P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S115N029N005P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S115P045P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S115P045N004P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S115N045P014P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S116P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S116N004P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S116N004N006psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S116P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S116N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S116P064P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S116P064P042P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S116P064P066P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S116P045P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S116P045N004P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S116N045P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S116P007P025P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S116P007P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S116P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S116N057P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S116N057N026P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S116P015P012P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S116P015P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S116P019P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S116P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S116P019N018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S116P015P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S116P015N067P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S116N015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S116P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S116N016P058P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S116P031P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S116P031N010P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S116N031P035P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S116N031N035P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S117P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S117N004P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S117N004N006P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S117P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S117N027P047P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S117N027P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S117P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S117P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S117P026P066P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S117N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S117N026N029P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S117P025P048P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S117P025N048P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S117N025P046P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S117N025P046P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S117P052P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S117P052N017P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S117P068P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S118P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S118P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S118P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S118N025P068P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S118P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S118N005P008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S118N005N008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S118P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S118N058P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S118N058N039P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S118P005P004P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S118P005P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S118P005N014P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S118P057P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S118P057N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S118P016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S118P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S118N015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S118P010P003P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S118N010P009P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S118N010N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S119P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S119P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S119P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S119N025P051P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S119N025P051P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S119P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S119N005P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S119P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S119N004P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S119N004N039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S119P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S119N048P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S119N048N063P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S119P023P020P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S119P023P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S119P023N056P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S119P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S120P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S120P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S120P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S120P008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S120N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S120N008N011P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S120P047P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S120P047N034P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S120P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S120P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S120N023P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S120N023N040P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S120P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S120N002P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S120N002N058P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S120P023P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S120N023P003P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S120P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S120P023P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S120P023N056P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S120P026P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S121P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S121P008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S121N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S121N008N011P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S121P047P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S121P047N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S121P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S121P013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S121P014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S121N014P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S121N014N051P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S121P012P056P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S121N012P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S121P026P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S122P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S122N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S122N006N004P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S122P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S122N043P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S122P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S122N022P023P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S122N022N023P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S122P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S122N004P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S122N004P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S122P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S122N007P008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S122N007N008P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S122P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S122N027P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S122N027P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S122P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S122N051P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S122N051N004P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S122P012P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S122P012N056P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S122N012P032P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S122N012P032P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S122P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S122N069P014P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S123P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S123N004P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S123N004N025P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S123P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S123N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S123N006N005P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S123P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S123N007P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S123N007N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S123P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S123N027P047P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S123N027P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S123P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S123N022P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S123P004P013P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S123N004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S123N004N006P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S123P009P050P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S123P009N050P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S123P026P014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S124P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S124N025P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S124N025N058P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S124P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S124N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S124N006N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S124P025P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S124P025N043P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S124N025P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S124N025N001P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S124P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S124N004P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S124N004N006P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S124P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S124N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S124N026N027P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S124P019P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S124P019P046P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S124N019P016P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S124N019N016psss: std_logic_vector(   0 downto 0);
        signal cVar2S22S124P026P014P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S125P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S125N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S125N006N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S125P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S125N004P006P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S125N004N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S125P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S125N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S125P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S125P030N057P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S125P059P038P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S125P059N038P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S126P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S126N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S126N004N007P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S126P050P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S126P050N039P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S126P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S126N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S126N006N004P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S126P025P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S126P025N043P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S126N025P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S126N025N036P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S126P006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S126P009P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S126P009P051P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S126N009P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S126N009N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S126P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S126P043P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S126P043N003P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S126P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S126N043P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S127P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S127P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S127N053P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S127N053N002P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S127P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S127N006P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S127N006N005P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S127P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S127N007P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S127N007N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S127P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S127N027P047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S127N027P047P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S127P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S127N006P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S127N006N004P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S127P025P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S127P025N043P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S127N025P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S127N025N011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S127P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S127N003P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S127N003N048P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S127P039P047P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S127P039P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S127P039N021P016nsss: std_logic_vector(   0 downto 0);
        signal oVar1S0: std_logic_vector(   0 downto 0);
        signal oVar1S1: std_logic_vector(   0 downto 0);
        signal oVar1S2: std_logic_vector(   0 downto 0);
        signal oVar1S3: std_logic_vector(   0 downto 0);
        signal oVar1S4: std_logic_vector(   0 downto 0);
        signal oVar1S5: std_logic_vector(   0 downto 0);
        signal oVar1S7: std_logic_vector(   0 downto 0);
        signal oVar1S8: std_logic_vector(   0 downto 0);
        signal oVar1S9: std_logic_vector(   0 downto 0);
        signal oVar1S10: std_logic_vector(   0 downto 0);
        signal oVar1S11: std_logic_vector(   0 downto 0);
        signal oVar1S12: std_logic_vector(   0 downto 0);
        signal oVar1S13: std_logic_vector(   0 downto 0);
        signal oVar1S14: std_logic_vector(   0 downto 0);
        signal oVar1S15: std_logic_vector(   0 downto 0);
        signal oVar1S16: std_logic_vector(   0 downto 0);
        signal oVar1S17: std_logic_vector(   0 downto 0);
        signal oVar1S18: std_logic_vector(   0 downto 0);
        signal oVar1S19: std_logic_vector(   0 downto 0);
        signal oVar1S20: std_logic_vector(   0 downto 0);
        signal oVar1S21: std_logic_vector(   0 downto 0);
        signal oVar1S22: std_logic_vector(   0 downto 0);
        signal oVar1S23: std_logic_vector(   0 downto 0);
        signal oVar1S24: std_logic_vector(   0 downto 0);
        signal oVar1S25: std_logic_vector(   0 downto 0);
        signal oVar1S26: std_logic_vector(   0 downto 0);
        signal oVar1S27: std_logic_vector(   0 downto 0);
        signal oVar1S28: std_logic_vector(   0 downto 0);
        signal oVar1S29: std_logic_vector(   0 downto 0);
        signal oVar1S30: std_logic_vector(   0 downto 0);
        signal oVar1S31: std_logic_vector(   0 downto 0);
        signal oVar1S32: std_logic_vector(   0 downto 0);
        signal oVar1S33: std_logic_vector(   0 downto 0);
        signal oVar1S34: std_logic_vector(   0 downto 0);
        signal oVar1S35: std_logic_vector(   0 downto 0);
        signal oVar1S36: std_logic_vector(   0 downto 0);
        signal oVar1S37: std_logic_vector(   0 downto 0);
        signal oVar1S38: std_logic_vector(   0 downto 0);
        signal oVar1S39: std_logic_vector(   0 downto 0);
        signal oVar1S40: std_logic_vector(   0 downto 0);
        signal oVar1S41: std_logic_vector(   0 downto 0);
        signal oVar1S42: std_logic_vector(   0 downto 0);
        signal oVar1S43: std_logic_vector(   0 downto 0);
        signal oVar1S44: std_logic_vector(   0 downto 0);
        signal oVar1S45: std_logic_vector(   0 downto 0);
        signal oVar1S46: std_logic_vector(   0 downto 0);
        signal oVar1S47: std_logic_vector(   0 downto 0);
        signal oVar1S48: std_logic_vector(   0 downto 0);
        signal oVar1S49: std_logic_vector(   0 downto 0);
        signal oVar1S50: std_logic_vector(   0 downto 0);
        signal oVar1S51: std_logic_vector(   0 downto 0);
        signal oVar1S52: std_logic_vector(   0 downto 0);
        signal oVar1S53: std_logic_vector(   0 downto 0);
        signal oVar1S54: std_logic_vector(   0 downto 0);
        signal oVar1S55: std_logic_vector(   0 downto 0);
        signal oVar1S56: std_logic_vector(   0 downto 0);
        signal oVar1S57: std_logic_vector(   0 downto 0);
        signal oVar1S58: std_logic_vector(   0 downto 0);
        signal oVar1S59: std_logic_vector(   0 downto 0);
        signal oVar1S60: std_logic_vector(   0 downto 0);
        signal oVar1S61: std_logic_vector(   0 downto 0);
        signal oVar1S62: std_logic_vector(   0 downto 0);
        signal oVar1S63: std_logic_vector(   0 downto 0);
        signal oVar1S64: std_logic_vector(   0 downto 0);
        signal oVar1S65: std_logic_vector(   0 downto 0);
        signal oVar1S66: std_logic_vector(   0 downto 0);
        signal oVar1S67: std_logic_vector(   0 downto 0);
        signal oVar1S68: std_logic_vector(   0 downto 0);
        signal oVar1S69: std_logic_vector(   0 downto 0);
        signal oVar1S70: std_logic_vector(   0 downto 0);
        signal oVar1S71: std_logic_vector(   0 downto 0);
        signal oVar1S72: std_logic_vector(   0 downto 0);
        signal oVar1S73: std_logic_vector(   0 downto 0);
        signal oVar1S74: std_logic_vector(   0 downto 0);
        signal oVar1S75: std_logic_vector(   0 downto 0);
        signal oVar1S76: std_logic_vector(   0 downto 0);
        signal oVar1S77: std_logic_vector(   0 downto 0);
        signal oVar1S78: std_logic_vector(   0 downto 0);
        signal oVar1S79: std_logic_vector(   0 downto 0);
        signal oVar1S80: std_logic_vector(   0 downto 0);
        signal oVar1S81: std_logic_vector(   0 downto 0);
        signal oVar1S82: std_logic_vector(   0 downto 0);
        signal oVar1S83: std_logic_vector(   0 downto 0);
        signal oVar1S84: std_logic_vector(   0 downto 0);
        signal oVar1S85: std_logic_vector(   0 downto 0);
        signal oVar1S86: std_logic_vector(   0 downto 0);
        signal oVar1S87: std_logic_vector(   0 downto 0);
        signal oVar1S88: std_logic_vector(   0 downto 0);
        signal oVar1S89: std_logic_vector(   0 downto 0);
        signal oVar1S90: std_logic_vector(   0 downto 0);
        signal oVar1S91: std_logic_vector(   0 downto 0);
        signal oVar1S92: std_logic_vector(   0 downto 0);
        signal oVar1S93: std_logic_vector(   0 downto 0);
        signal oVar1S94: std_logic_vector(   0 downto 0);
        signal oVar1S95: std_logic_vector(   0 downto 0);
        signal oVar1S96: std_logic_vector(   0 downto 0);
        signal oVar1S97: std_logic_vector(   0 downto 0);
        signal oVar1S99: std_logic_vector(   0 downto 0);
        signal oVar1S100: std_logic_vector(   0 downto 0);
        signal oVar1S101: std_logic_vector(   0 downto 0);
        signal oVar1S102: std_logic_vector(   0 downto 0);
        signal oVar1S103: std_logic_vector(   0 downto 0);
        signal oVar1S104: std_logic_vector(   0 downto 0);
        signal oVar1S105: std_logic_vector(   0 downto 0);
        signal oVar1S106: std_logic_vector(   0 downto 0);
        signal oVar1S107: std_logic_vector(   0 downto 0);
        signal oVar1S108: std_logic_vector(   0 downto 0);
        signal oVar1S109: std_logic_vector(   0 downto 0);
        signal oVar1S110: std_logic_vector(   0 downto 0);
        signal oVar1S111: std_logic_vector(   0 downto 0);
        signal oVar1S112: std_logic_vector(   0 downto 0);
        signal oVar1S113: std_logic_vector(   0 downto 0);
        signal oVar1S114: std_logic_vector(   0 downto 0);
        signal oVar1S115: std_logic_vector(   0 downto 0);
        signal oVar1S116: std_logic_vector(   0 downto 0);
        signal oVar1S117: std_logic_vector(   0 downto 0);
        signal oVar1S118: std_logic_vector(   0 downto 0);
        signal oVar1S119: std_logic_vector(   0 downto 0);
        signal oVar1S120: std_logic_vector(   0 downto 0);
        signal oVar1S121: std_logic_vector(   0 downto 0);
        signal oVar1S122: std_logic_vector(   0 downto 0);
        signal oVar1S123: std_logic_vector(   0 downto 0);
        signal oVar1S124: std_logic_vector(   0 downto 0);
        signal oVar1S125: std_logic_vector(   0 downto 0);
        signal oVar1S126: std_logic_vector(   0 downto 0);
        signal oVar1S127: std_logic_vector(   0 downto 0);
        signal oVar1S128: std_logic_vector(   0 downto 0);
        signal oVar1S129: std_logic_vector(   0 downto 0);
        signal oVar1S130: std_logic_vector(   0 downto 0);
        signal oVar1S131: std_logic_vector(   0 downto 0);
        signal oVar1S132: std_logic_vector(   0 downto 0);
        signal oVar1S133: std_logic_vector(   0 downto 0);
        signal oVar1S134: std_logic_vector(   0 downto 0);
        signal oVar1S135: std_logic_vector(   0 downto 0);
        signal oVar1S136: std_logic_vector(   0 downto 0);
        signal oVar1S137: std_logic_vector(   0 downto 0);
        signal oVar1S138: std_logic_vector(   0 downto 0);
        signal oVar1S139: std_logic_vector(   0 downto 0);
        signal oVar1S140: std_logic_vector(   0 downto 0);
        signal oVar1S141: std_logic_vector(   0 downto 0);
        signal oVar1S142: std_logic_vector(   0 downto 0);
        signal oVar1S143: std_logic_vector(   0 downto 0);
        signal oVar1S144: std_logic_vector(   0 downto 0);
        signal oVar1S145: std_logic_vector(   0 downto 0);
        signal oVar1S146: std_logic_vector(   0 downto 0);
        signal oVar1S147: std_logic_vector(   0 downto 0);
        signal oVar1S148: std_logic_vector(   0 downto 0);
        signal oVar1S149: std_logic_vector(   0 downto 0);
        signal oVar1S150: std_logic_vector(   0 downto 0);
        signal oVar1S151: std_logic_vector(   0 downto 0);
        signal oVar1S152: std_logic_vector(   0 downto 0);
        signal oVar1S153: std_logic_vector(   0 downto 0);
        signal oVar1S154: std_logic_vector(   0 downto 0);
        signal oVar1S155: std_logic_vector(   0 downto 0);
        signal oVar1S156: std_logic_vector(   0 downto 0);
        signal oVar1S157: std_logic_vector(   0 downto 0);
        signal oVar1S158: std_logic_vector(   0 downto 0);
        signal oVar1S160: std_logic_vector(   0 downto 0);
        signal oVar1S161: std_logic_vector(   0 downto 0);
        signal oVar1S162: std_logic_vector(   0 downto 0);
        signal oVar1S163: std_logic_vector(   0 downto 0);
        signal oVar1S164: std_logic_vector(   0 downto 0);
        signal oVar1S166: std_logic_vector(   0 downto 0);
        signal oVar1S167: std_logic_vector(   0 downto 0);
        signal oVar1S168: std_logic_vector(   0 downto 0);
        signal oVar1S169: std_logic_vector(   0 downto 0);
        signal oVar1S170: std_logic_vector(   0 downto 0);
        signal oVar1S171: std_logic_vector(   0 downto 0);
        signal oVar1S172: std_logic_vector(   0 downto 0);
        signal oVar1S173: std_logic_vector(   0 downto 0);
        signal oVar1S174: std_logic_vector(   0 downto 0);
        signal oVar1S175: std_logic_vector(   0 downto 0);
        signal oVar1S176: std_logic_vector(   0 downto 0);
        signal oVar1S177: std_logic_vector(   0 downto 0);
        signal oVar1S178: std_logic_vector(   0 downto 0);
        signal oVar1S179: std_logic_vector(   0 downto 0);
        signal oVar1S180: std_logic_vector(   0 downto 0);
        signal oVar1S181: std_logic_vector(   0 downto 0);
        signal oVar1S182: std_logic_vector(   0 downto 0);
        signal oVar1S183: std_logic_vector(   0 downto 0);
        signal oVar1S184: std_logic_vector(   0 downto 0);
        signal oVar1S185: std_logic_vector(   0 downto 0);
        signal oVar1S187: std_logic_vector(   0 downto 0);
        signal oVar1S188: std_logic_vector(   0 downto 0);
        signal oVar1S189: std_logic_vector(   0 downto 0);
        signal oVar1S190: std_logic_vector(   0 downto 0);
        signal oVar1S191: std_logic_vector(   0 downto 0);
        signal oVar1S192: std_logic_vector(   0 downto 0);
        signal oVar1S193: std_logic_vector(   0 downto 0);
        signal oVar1S194: std_logic_vector(   0 downto 0);
        signal oVar1S195: std_logic_vector(   0 downto 0);
        signal oVar1S196: std_logic_vector(   0 downto 0);
        signal oVar1S197: std_logic_vector(   0 downto 0);
        signal oVar1S198: std_logic_vector(   0 downto 0);
        signal oVar1S199: std_logic_vector(   0 downto 0);
        signal oVar1S200: std_logic_vector(   0 downto 0);
        signal oVar1S201: std_logic_vector(   0 downto 0);
        signal oVar1S202: std_logic_vector(   0 downto 0);
        signal oVar1S203: std_logic_vector(   0 downto 0);
        signal oVar1S204: std_logic_vector(   0 downto 0);
        signal oVar1S205: std_logic_vector(   0 downto 0);
        signal oVar1S206: std_logic_vector(   0 downto 0);
        signal oVar1S208: std_logic_vector(   0 downto 0);
        signal oVar1S209: std_logic_vector(   0 downto 0);
        signal oVar1S210: std_logic_vector(   0 downto 0);
        signal oVar1S211: std_logic_vector(   0 downto 0);
        signal oVar1S212: std_logic_vector(   0 downto 0);
        signal oVar1S213: std_logic_vector(   0 downto 0);
        signal oVar1S214: std_logic_vector(   0 downto 0);
        signal oVar1S215: std_logic_vector(   0 downto 0);
        signal oVar1S216: std_logic_vector(   0 downto 0);
        signal oVar1S217: std_logic_vector(   0 downto 0);
        signal oVar1S218: std_logic_vector(   0 downto 0);
        signal oVar1S219: std_logic_vector(   0 downto 0);
        signal oVar1S220: std_logic_vector(   0 downto 0);
        signal oVar1S221: std_logic_vector(   0 downto 0);
        signal oVar1S222: std_logic_vector(   0 downto 0);
        signal oVar1S223: std_logic_vector(   0 downto 0);
        signal oVar1S224: std_logic_vector(   0 downto 0);
        signal oVar1S225: std_logic_vector(   0 downto 0);
        signal oVar1S226: std_logic_vector(   0 downto 0);
        signal oVar1S227: std_logic_vector(   0 downto 0);
        signal oVar1S228: std_logic_vector(   0 downto 0);
        signal oVar1S229: std_logic_vector(   0 downto 0);
        signal oVar1S230: std_logic_vector(   0 downto 0);
        signal oVar1S231: std_logic_vector(   0 downto 0);
        signal oVar1S232: std_logic_vector(   0 downto 0);
        signal oVar1S233: std_logic_vector(   0 downto 0);
        signal oVar1S234: std_logic_vector(   0 downto 0);
        signal oVar1S235: std_logic_vector(   0 downto 0);
        signal oVar1S236: std_logic_vector(   0 downto 0);
        signal oVar1S237: std_logic_vector(   0 downto 0);
        signal oVar1S238: std_logic_vector(   0 downto 0);
        signal oVar1S239: std_logic_vector(   0 downto 0);
        signal oVar1S240: std_logic_vector(   0 downto 0);
        signal oVar1S241: std_logic_vector(   0 downto 0);
        signal oVar1S243: std_logic_vector(   0 downto 0);
        signal oVar1S244: std_logic_vector(   0 downto 0);
        signal oVar1S245: std_logic_vector(   0 downto 0);
        signal oVar1S246: std_logic_vector(   0 downto 0);
        signal oVar1S247: std_logic_vector(   0 downto 0);
        signal oVar1S248: std_logic_vector(   0 downto 0);
        signal oVar1S249: std_logic_vector(   0 downto 0);
        signal oVar1S250: std_logic_vector(   0 downto 0);
        signal oVar1S251: std_logic_vector(   0 downto 0);
        signal oVar1S252: std_logic_vector(   0 downto 0);
        signal oVar1S253: std_logic_vector(   0 downto 0);
        signal oVar1S254: std_logic_vector(   0 downto 0);
        signal oVar1S255: std_logic_vector(   0 downto 0);
        signal oVar1S256: std_logic_vector(   0 downto 0);
        signal oVar1S257: std_logic_vector(   0 downto 0);
        signal oVar1S258: std_logic_vector(   0 downto 0);
        signal oVar1S259: std_logic_vector(   0 downto 0);
        signal oVar1S260: std_logic_vector(   0 downto 0);
        signal oVar1S261: std_logic_vector(   0 downto 0);
        signal oVar1S262: std_logic_vector(   0 downto 0);
        signal oVar1S263: std_logic_vector(   0 downto 0);
        signal oVar1S264: std_logic_vector(   0 downto 0);
        signal oVar1S265: std_logic_vector(   0 downto 0);
        signal oVar1S266: std_logic_vector(   0 downto 0);
        signal oVar1S267: std_logic_vector(   0 downto 0);
        signal oVar1S268: std_logic_vector(   0 downto 0);
        signal oVar1S269: std_logic_vector(   0 downto 0);
        signal oVar1S270: std_logic_vector(   0 downto 0);
        signal oVar1S271: std_logic_vector(   0 downto 0);
        signal oVar1S272: std_logic_vector(   0 downto 0);
        signal oVar1S273: std_logic_vector(   0 downto 0);
        signal oVar1S274: std_logic_vector(   0 downto 0);
        signal oVar1S275: std_logic_vector(   0 downto 0);
        signal oVar1S276: std_logic_vector(   0 downto 0);
        signal oVar1S277: std_logic_vector(   0 downto 0);
        signal oVar1S278: std_logic_vector(   0 downto 0);
        signal oVar1S280: std_logic_vector(   0 downto 0);
        signal oVar1S281: std_logic_vector(   0 downto 0);
        signal oVar1S282: std_logic_vector(   0 downto 0);
        signal oVar1S283: std_logic_vector(   0 downto 0);
        signal oVar1S284: std_logic_vector(   0 downto 0);
        signal oVar1S285: std_logic_vector(   0 downto 0);
        signal oVar1S286: std_logic_vector(   0 downto 0);
        signal oVar1S287: std_logic_vector(   0 downto 0);
        signal oVar1S288: std_logic_vector(   0 downto 0);
        signal oVar1S289: std_logic_vector(   0 downto 0);
        signal oVar1S290: std_logic_vector(   0 downto 0);
        signal oVar1S291: std_logic_vector(   0 downto 0);
        signal oVar1S292: std_logic_vector(   0 downto 0);
        signal oVar1S293: std_logic_vector(   0 downto 0);
        signal oVar1S294: std_logic_vector(   0 downto 0);
        signal oVar1S295: std_logic_vector(   0 downto 0);
        signal oVar1S296: std_logic_vector(   0 downto 0);
        signal oVar1S297: std_logic_vector(   0 downto 0);
        signal oVar1S298: std_logic_vector(   0 downto 0);
        signal oVar1S299: std_logic_vector(   0 downto 0);
        signal oVar1S300: std_logic_vector(   0 downto 0);
        signal oVar1S301: std_logic_vector(   0 downto 0);
        signal oVar1S302: std_logic_vector(   0 downto 0);
        signal oVar1S303: std_logic_vector(   0 downto 0);
        signal oVar1S304: std_logic_vector(   0 downto 0);
        signal oVar1S305: std_logic_vector(   0 downto 0);
        signal oVar1S306: std_logic_vector(   0 downto 0);
        signal oVar1S307: std_logic_vector(   0 downto 0);
        signal oVar1S308: std_logic_vector(   0 downto 0);
        signal oVar1S309: std_logic_vector(   0 downto 0);
        signal oVar1S310: std_logic_vector(   0 downto 0);
        signal oVar1S312: std_logic_vector(   0 downto 0);
        signal oVar1S313: std_logic_vector(   0 downto 0);
        signal oVar1S314: std_logic_vector(   0 downto 0);
        signal oVar1S315: std_logic_vector(   0 downto 0);
        signal oVar1S316: std_logic_vector(   0 downto 0);
        signal oVar1S317: std_logic_vector(   0 downto 0);
        signal oVar1S318: std_logic_vector(   0 downto 0);
        signal oVar1S319: std_logic_vector(   0 downto 0);
        signal oVar1S320: std_logic_vector(   0 downto 0);
        signal oVar1S321: std_logic_vector(   0 downto 0);
        signal oVar1S322: std_logic_vector(   0 downto 0);
        signal oVar1S323: std_logic_vector(   0 downto 0);
        signal oVar1S324: std_logic_vector(   0 downto 0);
        signal oVar1S325: std_logic_vector(   0 downto 0);
        signal oVar1S326: std_logic_vector(   0 downto 0);
        signal oVar1S327: std_logic_vector(   0 downto 0);
        signal oVar1S328: std_logic_vector(   0 downto 0);
        signal oVar1S329: std_logic_vector(   0 downto 0);
        signal oVar1S330: std_logic_vector(   0 downto 0);
        signal oVar1S331: std_logic_vector(   0 downto 0);
        signal oVar1S332: std_logic_vector(   0 downto 0);
        signal oVar1S333: std_logic_vector(   0 downto 0);
        signal oVar1S334: std_logic_vector(   0 downto 0);
        signal oVar1S335: std_logic_vector(   0 downto 0);
        signal oVar1S336: std_logic_vector(   0 downto 0);
        signal oVar1S337: std_logic_vector(   0 downto 0);
        signal oVar1S338: std_logic_vector(   0 downto 0);
        signal oVar1S339: std_logic_vector(   0 downto 0);
        signal oVar1S340: std_logic_vector(   0 downto 0);
        signal oVar1S341: std_logic_vector(   0 downto 0);
        signal oVar1S342: std_logic_vector(   0 downto 0);
        signal oVar1S343: std_logic_vector(   0 downto 0);
        signal oVar1S345: std_logic_vector(   0 downto 0);
        signal oVar1S346: std_logic_vector(   0 downto 0);
        signal oVar1S347: std_logic_vector(   0 downto 0);
        signal oVar1S348: std_logic_vector(   0 downto 0);
        signal oVar1S349: std_logic_vector(   0 downto 0);
        signal oVar1S350: std_logic_vector(   0 downto 0);
        signal oVar1S351: std_logic_vector(   0 downto 0);
        signal oVar1S352: std_logic_vector(   0 downto 0);
        signal oVar1S354: std_logic_vector(   0 downto 0);
        signal oVar1S355: std_logic_vector(   0 downto 0);
        signal oVar1S356: std_logic_vector(   0 downto 0);
        signal oVar1S357: std_logic_vector(   0 downto 0);
        signal oVar1S358: std_logic_vector(   0 downto 0);
        signal oVar1S359: std_logic_vector(   0 downto 0);
        signal oVar1S360: std_logic_vector(   0 downto 0);
        signal oVar1S361: std_logic_vector(   0 downto 0);
        signal oVar1S362: std_logic_vector(   0 downto 0);
        signal oVar1S363: std_logic_vector(   0 downto 0);
        signal oVar1S364: std_logic_vector(   0 downto 0);
        signal oVar1S365: std_logic_vector(   0 downto 0);
        signal oVar1S367: std_logic_vector(   0 downto 0);
        signal oVar1S368: std_logic_vector(   0 downto 0);
        signal oVar1S369: std_logic_vector(   0 downto 0);
        signal oVar1S370: std_logic_vector(   0 downto 0);
        signal oVar1S371: std_logic_vector(   0 downto 0);
        signal oVar1S372: std_logic_vector(   0 downto 0);
        signal oVar1S373: std_logic_vector(   0 downto 0);
        signal oVar1S374: std_logic_vector(   0 downto 0);
        signal oVar1S375: std_logic_vector(   0 downto 0);
        signal oVar1S376: std_logic_vector(   0 downto 0);
        signal oVar1S377: std_logic_vector(   0 downto 0);
        signal oVar1S378: std_logic_vector(   0 downto 0);
        signal oVar1S379: std_logic_vector(   0 downto 0);
        signal oVar1S380: std_logic_vector(   0 downto 0);
        signal oVar1S381: std_logic_vector(   0 downto 0);
        signal oVar1S382: std_logic_vector(   0 downto 0);
        signal oVar1S383: std_logic_vector(   0 downto 0);
        signal oVar1S384: std_logic_vector(   0 downto 0);
        signal oVar1S385: std_logic_vector(   0 downto 0);
        signal oVar1S387: std_logic_vector(   0 downto 0);
        signal oVar1S388: std_logic_vector(   0 downto 0);
        signal oVar1S389: std_logic_vector(   0 downto 0);
        signal oVar1S390: std_logic_vector(   0 downto 0);
        signal oVar1S391: std_logic_vector(   0 downto 0);
        signal oVar1S392: std_logic_vector(   0 downto 0);
        signal oVar1S393: std_logic_vector(   0 downto 0);
        signal oVar1S394: std_logic_vector(   0 downto 0);
        signal oVar1S395: std_logic_vector(   0 downto 0);
        signal oVar1S396: std_logic_vector(   0 downto 0);
        signal oVar1S397: std_logic_vector(   0 downto 0);
        signal oVar1S398: std_logic_vector(   0 downto 0);
        signal oVar1S399: std_logic_vector(   0 downto 0);
        signal oVar1S400: std_logic_vector(   0 downto 0);
        signal oVar1S401: std_logic_vector(   0 downto 0);
        signal oVar1S402: std_logic_vector(   0 downto 0);
        signal oVar1S403: std_logic_vector(   0 downto 0);
        signal oVar1S404: std_logic_vector(   0 downto 0);
        signal oVar1S405: std_logic_vector(   0 downto 0);
        signal oVar1S406: std_logic_vector(   0 downto 0);
        signal oVar1S407: std_logic_vector(   0 downto 0);
        signal oVar1S408: std_logic_vector(   0 downto 0);
        signal oVar1S409: std_logic_vector(   0 downto 0);
        signal oVar1S410: std_logic_vector(   0 downto 0);
        signal oVar1S411: std_logic_vector(   0 downto 0);
        signal oVar1S412: std_logic_vector(   0 downto 0);
        signal oVar1S413: std_logic_vector(   0 downto 0);
        signal oVar1S414: std_logic_vector(   0 downto 0);
        signal oVar1S415: std_logic_vector(   0 downto 0);
        signal oVar1S416: std_logic_vector(   0 downto 0);
        signal oVar1S417: std_logic_vector(   0 downto 0);
        signal oVar1S418: std_logic_vector(   0 downto 0);
        signal oVar1S419: std_logic_vector(   0 downto 0);
        signal oVar1S420: std_logic_vector(   0 downto 0);
        signal oVar1S421: std_logic_vector(   0 downto 0);
        signal oVar1S422: std_logic_vector(   0 downto 0);
        signal oVar1S423: std_logic_vector(   0 downto 0);
        signal oVar1S424: std_logic_vector(   0 downto 0);
        signal oVar1S425: std_logic_vector(   0 downto 0);
        signal oVar1S426: std_logic_vector(   0 downto 0);
        signal oVar1S427: std_logic_vector(   0 downto 0);
        signal oVar1S428: std_logic_vector(   0 downto 0);
        signal oVar1S429: std_logic_vector(   0 downto 0);
        signal oVar1S430: std_logic_vector(   0 downto 0);
        signal oVar1S431: std_logic_vector(   0 downto 0);
        signal oVar1S432: std_logic_vector(   0 downto 0);
        signal oVar1S433: std_logic_vector(   0 downto 0);
        signal oVar1S434: std_logic_vector(   0 downto 0);
        signal oVar1S435: std_logic_vector(   0 downto 0);
        signal oVar1S436: std_logic_vector(   0 downto 0);
        signal oVar1S437: std_logic_vector(   0 downto 0);
        signal oVar1S438: std_logic_vector(   0 downto 0);
        signal oVar1S439: std_logic_vector(   0 downto 0);
        signal oVar1S440: std_logic_vector(   0 downto 0);
        signal oVar1S441: std_logic_vector(   0 downto 0);
        signal oVar1S442: std_logic_vector(   0 downto 0);
        signal oVar1S443: std_logic_vector(   0 downto 0);
        signal oVar1S444: std_logic_vector(   0 downto 0);
        signal oVar1S445: std_logic_vector(   0 downto 0);
        signal oVar1S446: std_logic_vector(   0 downto 0);
        signal oVar1S447: std_logic_vector(   0 downto 0);
        signal oVar1S448: std_logic_vector(   0 downto 0);
        signal oVar1S449: std_logic_vector(   0 downto 0);
        signal oVar1S450: std_logic_vector(   0 downto 0);
        signal oVar1S451: std_logic_vector(   0 downto 0);
        signal oVar1S452: std_logic_vector(   0 downto 0);
        signal oVar1S453: std_logic_vector(   0 downto 0);
        signal oVar1S454: std_logic_vector(   0 downto 0);
        signal oVar1S455: std_logic_vector(   0 downto 0);
        signal oVar1S456: std_logic_vector(   0 downto 0);
        signal oVar1S457: std_logic_vector(   0 downto 0);
        signal oVar1S458: std_logic_vector(   0 downto 0);
        signal oVar1S459: std_logic_vector(   0 downto 0);
        signal oVar1S460: std_logic_vector(   0 downto 0);
        signal oVar1S461: std_logic_vector(   0 downto 0);
        signal oVar1S462: std_logic_vector(   0 downto 0);
        signal oVar1S463: std_logic_vector(   0 downto 0);
        signal oVar1S464: std_logic_vector(   0 downto 0);
        signal oVar1S465: std_logic_vector(   0 downto 0);
        signal oVar1S466: std_logic_vector(   0 downto 0);
        signal oVar1S467: std_logic_vector(   0 downto 0);
        signal oVar1S468: std_logic_vector(   0 downto 0);
        signal oVar1S469: std_logic_vector(   0 downto 0);
        signal oVar1S470: std_logic_vector(   0 downto 0);
        signal oVar1S471: std_logic_vector(   0 downto 0);
        signal oVar1S472: std_logic_vector(   0 downto 0);
        signal oVar1S473: std_logic_vector(   0 downto 0);
        signal oVar1S474: std_logic_vector(   0 downto 0);
        signal oVar1S475: std_logic_vector(   0 downto 0);
        signal oVar1S476: std_logic_vector(   0 downto 0);
        signal oVar1S477: std_logic_vector(   0 downto 0);
        signal oVar1S478: std_logic_vector(   0 downto 0);
        signal oVar1S479: std_logic_vector(   0 downto 0);
        signal oVar1S480: std_logic_vector(   0 downto 0);
        signal oVar1S481: std_logic_vector(   0 downto 0);
        signal oVar1S482: std_logic_vector(   0 downto 0);
        signal oVar1S483: std_logic_vector(   0 downto 0);
        signal oVar1S484: std_logic_vector(   0 downto 0);
        signal oVar1S485: std_logic_vector(   0 downto 0);
        signal oVar1S486: std_logic_vector(   0 downto 0);
        signal oVar1S487: std_logic_vector(   0 downto 0);
        signal oVar1S488: std_logic_vector(   0 downto 0);
        signal oVar1S489: std_logic_vector(   0 downto 0);
        signal oVar1S490: std_logic_vector(   0 downto 0);
        signal oVar1S491: std_logic_vector(   0 downto 0);
        signal oVar1S493: std_logic_vector(   0 downto 0);
        signal oVar1S494: std_logic_vector(   0 downto 0);
        signal oVar1S495: std_logic_vector(   0 downto 0);
        signal oVar1S496: std_logic_vector(   0 downto 0);
        signal oVar1S497: std_logic_vector(   0 downto 0);
        signal oVar1S498: std_logic_vector(   0 downto 0);
        signal oVar1S499: std_logic_vector(   0 downto 0);
        signal oVar1S500: std_logic_vector(   0 downto 0);
        signal oVar1S502: std_logic_vector(   0 downto 0);
        signal oVar1S503: std_logic_vector(   0 downto 0);
        signal oVar1S504: std_logic_vector(   0 downto 0);
        signal oVar1S505: std_logic_vector(   0 downto 0);
        signal oVar1S506: std_logic_vector(   0 downto 0);
        signal oVar1S507: std_logic_vector(   0 downto 0);
        signal oVar1S508: std_logic_vector(   0 downto 0);
        signal oVar1S510: std_logic_vector(   0 downto 0);
        signal oVar1S511: std_logic_vector(   0 downto 0);
        signal oVar1S512: std_logic_vector(   0 downto 0);
        signal oVar1S513: std_logic_vector(   0 downto 0);
        signal oVar1S514: std_logic_vector(   0 downto 0);
        signal oVar1S515: std_logic_vector(   0 downto 0);
        signal oVar1S516: std_logic_vector(   0 downto 0);
        signal oVar1S517: std_logic_vector(   0 downto 0);
        signal oVar1S518: std_logic_vector(   0 downto 0);
        signal oVar1S519: std_logic_vector(   0 downto 0);
        signal oVar1S520: std_logic_vector(   0 downto 0);
        signal oVar1S521: std_logic_vector(   0 downto 0);
        signal oVar1S522: std_logic_vector(   0 downto 0);
        signal oVar1S523: std_logic_vector(   0 downto 0);
        signal oVar1S524: std_logic_vector(   0 downto 0);
        signal oVar1S525: std_logic_vector(   0 downto 0);
        signal oVar1S526: std_logic_vector(   0 downto 0);
        signal oVar1S527: std_logic_vector(   0 downto 0);
        signal oVar1S528: std_logic_vector(   0 downto 0);
        signal oVar1S529: std_logic_vector(   0 downto 0);
        signal oVar1S530: std_logic_vector(   0 downto 0);
        signal oVar1S531: std_logic_vector(   0 downto 0);
        signal oVar1S532: std_logic_vector(   0 downto 0);
        signal oVar1S533: std_logic_vector(   0 downto 0);
        signal oVar1S534: std_logic_vector(   0 downto 0);
        signal oVar1S535: std_logic_vector(   0 downto 0);
        signal oVar1S536: std_logic_vector(   0 downto 0);
        signal oVar1S537: std_logic_vector(   0 downto 0);
        signal oVar1S538: std_logic_vector(   0 downto 0);
        signal oVar1S539: std_logic_vector(   0 downto 0);
        signal oVar1S540: std_logic_vector(   0 downto 0);
        signal oVar1S541: std_logic_vector(   0 downto 0);
        signal oVar1S542: std_logic_vector(   0 downto 0);
        signal oVar1S543: std_logic_vector(   0 downto 0);
        signal oVar1S544: std_logic_vector(   0 downto 0);
        signal oVar1S545: std_logic_vector(   0 downto 0);
        signal oVar1S546: std_logic_vector(   0 downto 0);
        signal oVar1S547: std_logic_vector(   0 downto 0);
        signal oVar1S549: std_logic_vector(   0 downto 0);
        signal oVar1S550: std_logic_vector(   0 downto 0);
        signal oVar1S551: std_logic_vector(   0 downto 0);
        signal oVar1S552: std_logic_vector(   0 downto 0);
        signal oVar1S553: std_logic_vector(   0 downto 0);
        signal oVar1S554: std_logic_vector(   0 downto 0);
        signal oVar1S555: std_logic_vector(   0 downto 0);
        signal oVar1S556: std_logic_vector(   0 downto 0);
        signal oVar1S557: std_logic_vector(   0 downto 0);
        signal oVar1S558: std_logic_vector(   0 downto 0);
        signal oVar1S559: std_logic_vector(   0 downto 0);
        signal oVar1S560: std_logic_vector(   0 downto 0);
        signal oVar1S561: std_logic_vector(   0 downto 0);
        signal oVar1S562: std_logic_vector(   0 downto 0);
        signal oVar1S563: std_logic_vector(   0 downto 0);
        signal oVar1S564: std_logic_vector(   0 downto 0);
        signal oVar1S565: std_logic_vector(   0 downto 0);
        signal oVar1S566: std_logic_vector(   0 downto 0);
        signal oVar1S567: std_logic_vector(   0 downto 0);
        signal oVar1S568: std_logic_vector(   0 downto 0);
        signal oVar1S569: std_logic_vector(   0 downto 0);
        signal oVar1S570: std_logic_vector(   0 downto 0);
        signal oVar1S571: std_logic_vector(   0 downto 0);
        signal oVar1S572: std_logic_vector(   0 downto 0);
        signal oVar1S573: std_logic_vector(   0 downto 0);
        signal oVar1S574: std_logic_vector(   0 downto 0);
        signal oVar1S575: std_logic_vector(   0 downto 0);
        signal oVar1S576: std_logic_vector(   0 downto 0);
        signal oVar1S577: std_logic_vector(   0 downto 0);
        signal oVar1S578: std_logic_vector(   0 downto 0);
        signal oVar1S579: std_logic_vector(   0 downto 0);
        signal oVar1S580: std_logic_vector(   0 downto 0);
        signal oVar1S581: std_logic_vector(   0 downto 0);
        signal oVar1S582: std_logic_vector(   0 downto 0);
        signal oVar1S583: std_logic_vector(   0 downto 0);
        signal oVar1S584: std_logic_vector(   0 downto 0);
        signal oVar1S585: std_logic_vector(   0 downto 0);
        signal oVar1S586: std_logic_vector(   0 downto 0);
        signal oVar1S587: std_logic_vector(   0 downto 0);
        signal oVar1S588: std_logic_vector(   0 downto 0);
        signal oVar1S589: std_logic_vector(   0 downto 0);
        signal oVar1S590: std_logic_vector(   0 downto 0);
        signal oVar1S591: std_logic_vector(   0 downto 0);
        signal oVar1S592: std_logic_vector(   0 downto 0);
        signal oVar1S593: std_logic_vector(   0 downto 0);
        signal oVar1S594: std_logic_vector(   0 downto 0);
        signal oVar1S595: std_logic_vector(   0 downto 0);
        signal oVar1S596: std_logic_vector(   0 downto 0);
        signal oVar1S597: std_logic_vector(   0 downto 0);
        signal oVar1S598: std_logic_vector(   0 downto 0);
        signal oVar1S599: std_logic_vector(   0 downto 0);
        signal oVar1S600: std_logic_vector(   0 downto 0);
        signal oVar1S601: std_logic_vector(   0 downto 0);
        signal oVar1S602: std_logic_vector(   0 downto 0);
        signal oVar1S603: std_logic_vector(   0 downto 0);
        signal oVar1S604: std_logic_vector(   0 downto 0);
        signal oVar1S605: std_logic_vector(   0 downto 0);
        signal oVar1S607: std_logic_vector(   0 downto 0);
        signal oVar1S608: std_logic_vector(   0 downto 0);
        signal oVar1S609: std_logic_vector(   0 downto 0);
        signal oVar1S610: std_logic_vector(   0 downto 0);
        signal oVar1S611: std_logic_vector(   0 downto 0);
        signal oVar1S612: std_logic_vector(   0 downto 0);
        signal oVar1S613: std_logic_vector(   0 downto 0);
        signal oVar1S614: std_logic_vector(   0 downto 0);
        signal oVar1S615: std_logic_vector(   0 downto 0);
        signal oVar1S616: std_logic_vector(   0 downto 0);
        signal oVar1S617: std_logic_vector(   0 downto 0);
        signal oVar1S618: std_logic_vector(   0 downto 0);
        signal oVar1S619: std_logic_vector(   0 downto 0);
        signal oVar1S620: std_logic_vector(   0 downto 0);
        signal oVar1S622: std_logic_vector(   0 downto 0);
        signal oVar1S623: std_logic_vector(   0 downto 0);
        signal oVar1S624: std_logic_vector(   0 downto 0);
        signal oVar1S625: std_logic_vector(   0 downto 0);
        signal oVar1S626: std_logic_vector(   0 downto 0);
        signal oVar1S627: std_logic_vector(   0 downto 0);
        signal oVar1S628: std_logic_vector(   0 downto 0);
        signal oVar1S629: std_logic_vector(   0 downto 0);
        signal oVar1S630: std_logic_vector(   0 downto 0);
        signal oVar1S631: std_logic_vector(   0 downto 0);
        signal oVar1S632: std_logic_vector(   0 downto 0);
        signal oVar1S633: std_logic_vector(   0 downto 0);
        signal oVar1S634: std_logic_vector(   0 downto 0);
        signal oVar1S635: std_logic_vector(   0 downto 0);
        signal oVar1S637: std_logic_vector(   0 downto 0);
        signal oVar1S638: std_logic_vector(   0 downto 0);
        signal oVar1S639: std_logic_vector(   0 downto 0);
        signal oVar1S640: std_logic_vector(   0 downto 0);
        signal oVar1S641: std_logic_vector(   0 downto 0);
        signal oVar1S642: std_logic_vector(   0 downto 0);
        signal oVar1S643: std_logic_vector(   0 downto 0);
        signal oVar1S644: std_logic_vector(   0 downto 0);
        signal oVar1S645: std_logic_vector(   0 downto 0);
        signal oVar1S646: std_logic_vector(   0 downto 0);
        signal oVar1S647: std_logic_vector(   0 downto 0);
        signal oVar1S648: std_logic_vector(   0 downto 0);
        signal oVar1S649: std_logic_vector(   0 downto 0);
        signal oVar1S650: std_logic_vector(   0 downto 0);
        signal oVar1S651: std_logic_vector(   0 downto 0);
        signal oVar1S652: std_logic_vector(   0 downto 0);
        signal oVar1S653: std_logic_vector(   0 downto 0);
        signal oVar1S654: std_logic_vector(   0 downto 0);
        signal oVar1S655: std_logic_vector(   0 downto 0);
        signal oVar1S656: std_logic_vector(   0 downto 0);
        signal oVar1S657: std_logic_vector(   0 downto 0);
        signal oVar1S658: std_logic_vector(   0 downto 0);
        signal oVar1S659: std_logic_vector(   0 downto 0);
        signal oVar1S660: std_logic_vector(   0 downto 0);
        signal oVar1S661: std_logic_vector(   0 downto 0);
        signal oVar1S662: std_logic_vector(   0 downto 0);
        signal oVar1S663: std_logic_vector(   0 downto 0);
        signal oVar1S664: std_logic_vector(   0 downto 0);
        signal oVar1S665: std_logic_vector(   0 downto 0);
        signal oVar1S666: std_logic_vector(   0 downto 0);
        signal oVar1S667: std_logic_vector(   0 downto 0);
        signal oVar1S668: std_logic_vector(   0 downto 0);
        signal oVar1S669: std_logic_vector(   0 downto 0);
        signal oVar1S670: std_logic_vector(   0 downto 0);
        signal oVar1S671: std_logic_vector(   0 downto 0);
        signal oVar1S672: std_logic_vector(   0 downto 0);
        signal oVar1S673: std_logic_vector(   0 downto 0);
        signal oVar1S674: std_logic_vector(   0 downto 0);
        signal oVar1S675: std_logic_vector(   0 downto 0);
        signal oVar1S676: std_logic_vector(   0 downto 0);
        signal oVar1S677: std_logic_vector(   0 downto 0);
        signal oVar1S678: std_logic_vector(   0 downto 0);
        signal oVar1S679: std_logic_vector(   0 downto 0);
        signal oVar1S680: std_logic_vector(   0 downto 0);
        signal oVar1S681: std_logic_vector(   0 downto 0);
        signal oVar1S682: std_logic_vector(   0 downto 0);
        signal oVar1S684: std_logic_vector(   0 downto 0);
        signal oVar1S685: std_logic_vector(   0 downto 0);
        signal oVar1S686: std_logic_vector(   0 downto 0);
        signal oVar1S687: std_logic_vector(   0 downto 0);
        signal oVar1S688: std_logic_vector(   0 downto 0);
        signal oVar1S689: std_logic_vector(   0 downto 0);
        signal oVar1S690: std_logic_vector(   0 downto 0);
        signal oVar1S691: std_logic_vector(   0 downto 0);
        signal oVar1S692: std_logic_vector(   0 downto 0);
        signal oVar1S693: std_logic_vector(   0 downto 0);
        signal oVar1S694: std_logic_vector(   0 downto 0);
        signal oVar1S695: std_logic_vector(   0 downto 0);
        signal oVar1S696: std_logic_vector(   0 downto 0);
        signal oVar1S697: std_logic_vector(   0 downto 0);
        signal oVar1S698: std_logic_vector(   0 downto 0);
        signal oVar1S699: std_logic_vector(   0 downto 0);
        signal oVar1S700: std_logic_vector(   0 downto 0);
        signal oVar1S701: std_logic_vector(   0 downto 0);
        signal oVar1S702: std_logic_vector(   0 downto 0);
        signal oVar1S703: std_logic_vector(   0 downto 0);
        signal oVar1S704: std_logic_vector(   0 downto 0);
        signal oVar1S705: std_logic_vector(   0 downto 0);
        signal oVar1S706: std_logic_vector(   0 downto 0);
        signal oVar1S707: std_logic_vector(   0 downto 0);
        signal oVar1S708: std_logic_vector(   0 downto 0);
        signal oVar1S709: std_logic_vector(   0 downto 0);
        signal oVar1S710: std_logic_vector(   0 downto 0);
        signal oVar1S711: std_logic_vector(   0 downto 0);
        signal oVar1S712: std_logic_vector(   0 downto 0);
        signal oVar1S714: std_logic_vector(   0 downto 0);
        signal oVar1S715: std_logic_vector(   0 downto 0);
        signal oVar1S716: std_logic_vector(   0 downto 0);
        signal oVar1S717: std_logic_vector(   0 downto 0);
        signal oVar1S718: std_logic_vector(   0 downto 0);
        signal oVar1S719: std_logic_vector(   0 downto 0);
        signal oVar1S720: std_logic_vector(   0 downto 0);
        signal oVar1S722: std_logic_vector(   0 downto 0);
        signal oVar1S723: std_logic_vector(   0 downto 0);
        signal oVar1S724: std_logic_vector(   0 downto 0);
        signal oVar1S725: std_logic_vector(   0 downto 0);
        signal oVar1S726: std_logic_vector(   0 downto 0);
        signal oVar1S727: std_logic_vector(   0 downto 0);
        signal oVar1S728: std_logic_vector(   0 downto 0);
        signal oVar1S729: std_logic_vector(   0 downto 0);
        signal oVar1S730: std_logic_vector(   0 downto 0);
        signal oVar1S731: std_logic_vector(   0 downto 0);
        signal oVar1S732: std_logic_vector(   0 downto 0);
        signal oVar1S733: std_logic_vector(   0 downto 0);
        signal oVar1S734: std_logic_vector(   0 downto 0);
        signal oVar1S735: std_logic_vector(   0 downto 0);
        signal oVar1S736: std_logic_vector(   0 downto 0);
        signal oVar1S737: std_logic_vector(   0 downto 0);
        signal oVar1S738: std_logic_vector(   0 downto 0);
        signal oVar1S739: std_logic_vector(   0 downto 0);
        signal oVar1S740: std_logic_vector(   0 downto 0);
        signal oVar1S741: std_logic_vector(   0 downto 0);
        signal oVar1S742: std_logic_vector(   0 downto 0);
        signal oVar1S743: std_logic_vector(   0 downto 0);
        signal oVar1S744: std_logic_vector(   0 downto 0);
        signal oVar1S746: std_logic_vector(   0 downto 0);
        signal oVar1S747: std_logic_vector(   0 downto 0);
        signal oVar1S748: std_logic_vector(   0 downto 0);
        signal oVar1S749: std_logic_vector(   0 downto 0);
        signal oVar1S750: std_logic_vector(   0 downto 0);
        signal oVar1S751: std_logic_vector(   0 downto 0);
        signal oVar1S752: std_logic_vector(   0 downto 0);
        signal oVar1S753: std_logic_vector(   0 downto 0);
        signal oVar1S754: std_logic_vector(   0 downto 0);
        signal oVar1S755: std_logic_vector(   0 downto 0);
        signal oVar1S756: std_logic_vector(   0 downto 0);
        signal oVar1S757: std_logic_vector(   0 downto 0);
        signal oVar1S758: std_logic_vector(   0 downto 0);
        signal oVar1S759: std_logic_vector(   0 downto 0);
        signal oVar1S760: std_logic_vector(   0 downto 0);
        signal oVar1S761: std_logic_vector(   0 downto 0);
        signal oVar1S762: std_logic_vector(   0 downto 0);
        signal oVar1S763: std_logic_vector(   0 downto 0);
        signal oVar1S764: std_logic_vector(   0 downto 0);
        signal oVar1S765: std_logic_vector(   0 downto 0);
        signal oVar1S766: std_logic_vector(   0 downto 0);
        signal oVar1S767: std_logic_vector(   0 downto 0);
        signal oVar1S768: std_logic_vector(   0 downto 0);
        signal oVar1S769: std_logic_vector(   0 downto 0);
        signal oVar1S770: std_logic_vector(   0 downto 0);
        signal oVar1S771: std_logic_vector(   0 downto 0);
        signal oVar1S772: std_logic_vector(   0 downto 0);
        signal oVar1S773: std_logic_vector(   0 downto 0);
        signal oVar1S774: std_logic_vector(   0 downto 0);
        signal oVar1S775: std_logic_vector(   0 downto 0);
        signal oVar1S776: std_logic_vector(   0 downto 0);
        signal oVar1S777: std_logic_vector(   0 downto 0);
        signal oVar1S778: std_logic_vector(   0 downto 0);
        signal oVar1S779: std_logic_vector(   0 downto 0);
        signal oVar1S780: std_logic_vector(   0 downto 0);
        signal oVar1S781: std_logic_vector(   0 downto 0);
        signal oVar1S782: std_logic_vector(   0 downto 0);
        signal oVar1S783: std_logic_vector(   0 downto 0);
        signal oVar1S784: std_logic_vector(   0 downto 0);
        signal oVar1S785: std_logic_vector(   0 downto 0);
        signal oVar1S786: std_logic_vector(   0 downto 0);
        signal oVar1S787: std_logic_vector(   0 downto 0);
        signal oVar1S788: std_logic_vector(   0 downto 0);
        signal oVar1S789: std_logic_vector(   0 downto 0);
        signal oVar1S790: std_logic_vector(   0 downto 0);
        signal oVar1S791: std_logic_vector(   0 downto 0);
        signal oVar1S792: std_logic_vector(   0 downto 0);
        signal oVar1S793: std_logic_vector(   0 downto 0);
        signal oVar1S794: std_logic_vector(   0 downto 0);
        signal oVar1S795: std_logic_vector(   0 downto 0);
        signal oVar1S796: std_logic_vector(   0 downto 0);
        signal oVar1S797: std_logic_vector(   0 downto 0);
        signal oVar1S798: std_logic_vector(   0 downto 0);
        signal oVar1S799: std_logic_vector(   0 downto 0);
        signal oVar1S800: std_logic_vector(   0 downto 0);
        signal oVar1S801: std_logic_vector(   0 downto 0);
        signal oVar1S802: std_logic_vector(   0 downto 0);
        signal oVar1S803: std_logic_vector(   0 downto 0);
        signal oVar1S804: std_logic_vector(   0 downto 0);
        signal oVar1S805: std_logic_vector(   0 downto 0);
        signal oVar1S806: std_logic_vector(   0 downto 0);
        signal oVar1S807: std_logic_vector(   0 downto 0);
        signal oVar1S808: std_logic_vector(   0 downto 0);
        signal oVar1S809: std_logic_vector(   0 downto 0);
        signal oVar1S810: std_logic_vector(   0 downto 0);
        signal oVar1S811: std_logic_vector(   0 downto 0);
        signal oVar1S812: std_logic_vector(   0 downto 0);
        signal oVar1S813: std_logic_vector(   0 downto 0);
        signal oVar1S814: std_logic_vector(   0 downto 0);
        signal oVar1S815: std_logic_vector(   0 downto 0);
        signal oVar1S816: std_logic_vector(   0 downto 0);
        signal oVar1S817: std_logic_vector(   0 downto 0);
        signal oVar1S818: std_logic_vector(   0 downto 0);
        signal oVar1S819: std_logic_vector(   0 downto 0);
        signal oVar1S820: std_logic_vector(   0 downto 0);
        signal oVar1S821: std_logic_vector(   0 downto 0);
        signal oVar1S822: std_logic_vector(   0 downto 0);
        signal oVar1S823: std_logic_vector(   0 downto 0);
        signal oVar1S824: std_logic_vector(   0 downto 0);
        signal oVar1S825: std_logic_vector(   0 downto 0);
        signal oVar1S826: std_logic_vector(   0 downto 0);
        signal oVar1S827: std_logic_vector(   0 downto 0);
        signal oVar1S828: std_logic_vector(   0 downto 0);
        signal oVar1S829: std_logic_vector(   0 downto 0);
        signal oVar1S830: std_logic_vector(   0 downto 0);
        signal oVar1S831: std_logic_vector(   0 downto 0);
        signal oVar1S832: std_logic_vector(   0 downto 0);
        signal oVar1S833: std_logic_vector(   0 downto 0);
        signal oVar1S834: std_logic_vector(   0 downto 0);
        signal oVar1S835: std_logic_vector(   0 downto 0);
        signal oVar1S836: std_logic_vector(   0 downto 0);
        signal oVar1S837: std_logic_vector(   0 downto 0);
        signal oVar1S838: std_logic_vector(   0 downto 0);
        signal oVar1S839: std_logic_vector(   0 downto 0);
        signal oVar1S840: std_logic_vector(   0 downto 0);
        signal oVar1S841: std_logic_vector(   0 downto 0);
        signal oVar1S842: std_logic_vector(   0 downto 0);
        signal oVar1S843: std_logic_vector(   0 downto 0);
        signal oVar1S844: std_logic_vector(   0 downto 0);
        signal oVar1S845: std_logic_vector(   0 downto 0);
        signal oVar1S846: std_logic_vector(   0 downto 0);
        signal oVar1S847: std_logic_vector(   0 downto 0);
        signal oVar1S848: std_logic_vector(   0 downto 0);
        signal oVar1S849: std_logic_vector(   0 downto 0);
        signal oVar1S850: std_logic_vector(   0 downto 0);
        signal oVar1S851: std_logic_vector(   0 downto 0);
        signal oVar1S852: std_logic_vector(   0 downto 0);
        signal oVar1S853: std_logic_vector(   0 downto 0);
        signal oVar1S854: std_logic_vector(   0 downto 0);
        signal oVar1S856: std_logic_vector(   0 downto 0);
        signal oVar1S857: std_logic_vector(   0 downto 0);
        signal oVar1S858: std_logic_vector(   0 downto 0);
        signal oVar1S859: std_logic_vector(   0 downto 0);
        signal oVar1S860: std_logic_vector(   0 downto 0);
        signal oVar1S861: std_logic_vector(   0 downto 0);
        signal oVar1S862: std_logic_vector(   0 downto 0);
        signal oVar1S863: std_logic_vector(   0 downto 0);
        signal oVar1S864: std_logic_vector(   0 downto 0);
        signal oVar1S865: std_logic_vector(   0 downto 0);
        signal oVar1S866: std_logic_vector(   0 downto 0);
        signal oVar1S867: std_logic_vector(   0 downto 0);
        signal oVar1S869: std_logic_vector(   0 downto 0);
        signal oVar1S870: std_logic_vector(   0 downto 0);
        signal oVar1S871: std_logic_vector(   0 downto 0);
        signal oVar1S872: std_logic_vector(   0 downto 0);
        signal oVar1S873: std_logic_vector(   0 downto 0);
        signal oVar1S874: std_logic_vector(   0 downto 0);
        signal oVar1S875: std_logic_vector(   0 downto 0);
        signal oVar1S876: std_logic_vector(   0 downto 0);
        signal oVar1S877: std_logic_vector(   0 downto 0);
        signal oVar1S878: std_logic_vector(   0 downto 0);
        signal oVar1S879: std_logic_vector(   0 downto 0);
        signal oVar1S880: std_logic_vector(   0 downto 0);
        signal oVar1S882: std_logic_vector(   0 downto 0);
        signal oVar1S883: std_logic_vector(   0 downto 0);
        signal oVar1S884: std_logic_vector(   0 downto 0);
        signal oVar1S885: std_logic_vector(   0 downto 0);
        signal oVar1S886: std_logic_vector(   0 downto 0);
        signal oVar1S887: std_logic_vector(   0 downto 0);
        signal oVar1S888: std_logic_vector(   0 downto 0);
        signal oVar1S889: std_logic_vector(   0 downto 0);
        signal oVar1S890: std_logic_vector(   0 downto 0);
        signal oVar1S891: std_logic_vector(   0 downto 0);
        signal oVar1S892: std_logic_vector(   0 downto 0);
        signal oVar1S893: std_logic_vector(   0 downto 0);
        signal oVar1S895: std_logic_vector(   0 downto 0);
        signal oVar1S896: std_logic_vector(   0 downto 0);
        signal oVar1S897: std_logic_vector(   0 downto 0);
        signal oVar1S898: std_logic_vector(   0 downto 0);
        signal oVar1S899: std_logic_vector(   0 downto 0);
        signal oVar1S900: std_logic_vector(   0 downto 0);
        signal oVar1S901: std_logic_vector(   0 downto 0);
        signal oVar1S902: std_logic_vector(   0 downto 0);
        signal oVar1S903: std_logic_vector(   0 downto 0);
        signal oVar1S904: std_logic_vector(   0 downto 0);
        signal oVar1S905: std_logic_vector(   0 downto 0);
        signal oVar1S906: std_logic_vector(   0 downto 0);
        signal oVar1S907: std_logic_vector(   0 downto 0);
        signal oVar1S908: std_logic_vector(   0 downto 0);
        signal oVar1S909: std_logic_vector(   0 downto 0);
        signal oVar1S910: std_logic_vector(   0 downto 0);
        signal oVar1S911: std_logic_vector(   0 downto 0);
        signal oVar1S912: std_logic_vector(   0 downto 0);
        signal oVar1S913: std_logic_vector(   0 downto 0);
        signal oVar1S914: std_logic_vector(   0 downto 0);
        signal oVar1S915: std_logic_vector(   0 downto 0);
        signal oVar1S916: std_logic_vector(   0 downto 0);
        signal oVar1S917: std_logic_vector(   0 downto 0);
        signal oVar1S918: std_logic_vector(   0 downto 0);
        signal oVar1S919: std_logic_vector(   0 downto 0);
        signal oVar1S920: std_logic_vector(   0 downto 0);
        signal oVar1S921: std_logic_vector(   0 downto 0);
        signal oVar1S922: std_logic_vector(   0 downto 0);
        signal oVar1S923: std_logic_vector(   0 downto 0);
        signal oVar1S924: std_logic_vector(   0 downto 0);
        signal oVar1S925: std_logic_vector(   0 downto 0);
        signal oVar2S0: std_logic_vector(   0 downto 0);
        signal oVar2S1: std_logic_vector(   0 downto 0);
        signal oVar2S2: std_logic_vector(   0 downto 0);
        signal oVar2S3: std_logic_vector(   0 downto 0);
        signal oVar2S4: std_logic_vector(   0 downto 0);
        signal oVar2S5: std_logic_vector(   0 downto 0);
        signal oVar2S6: std_logic_vector(   0 downto 0);
        signal oVar2S7: std_logic_vector(   0 downto 0);
        signal oVar2S9: std_logic_vector(   0 downto 0);
        signal oVar2S10: std_logic_vector(   0 downto 0);
        signal oVar2S11: std_logic_vector(   0 downto 0);
        signal oVar2S12: std_logic_vector(   0 downto 0);
        signal oVar2S13: std_logic_vector(   0 downto 0);
        signal oVar2S14: std_logic_vector(   0 downto 0);
        signal oVar2S15: std_logic_vector(   0 downto 0);
        signal oVar2S16: std_logic_vector(   0 downto 0);
        signal oVar2S17: std_logic_vector(   0 downto 0);
        signal oVar2S18: std_logic_vector(   0 downto 0);
        signal oVar2S20: std_logic_vector(   0 downto 0);
        signal oVar2S21: std_logic_vector(   0 downto 0);
        signal oVar2S22: std_logic_vector(   0 downto 0);
        signal oVar2S23: std_logic_vector(   0 downto 0);
        signal oVar2S24: std_logic_vector(   0 downto 0);
        signal oVar2S25: std_logic_vector(   0 downto 0);
        signal oVar2S26: std_logic_vector(   0 downto 0);
        signal oVar2S28: std_logic_vector(   0 downto 0);
        signal oVar2S29: std_logic_vector(   0 downto 0);
        signal oVar2S30: std_logic_vector(   0 downto 0);
        signal oVar2S31: std_logic_vector(   0 downto 0);
        signal oVar2S33: std_logic_vector(   0 downto 0);
        signal oVar2S34: std_logic_vector(   0 downto 0);
        signal oVar2S36: std_logic_vector(   0 downto 0);
        signal oVar2S37: std_logic_vector(   0 downto 0);
        signal oVar2S39: std_logic_vector(   0 downto 0);
        signal oVar2S40: std_logic_vector(   0 downto 0);
        signal oVar2S42: std_logic_vector(   0 downto 0);
        signal oVar2S43: std_logic_vector(   0 downto 0);
        signal oVar2S44: std_logic_vector(   0 downto 0);
        signal oVar2S45: std_logic_vector(   0 downto 0);
        signal oVar2S46: std_logic_vector(   0 downto 0);
        signal oVar2S47: std_logic_vector(   0 downto 0);
        signal oVar2S48: std_logic_vector(   0 downto 0);
        signal oVar2S49: std_logic_vector(   0 downto 0);
        signal oVar2S51: std_logic_vector(   0 downto 0);
        signal oVar2S52: std_logic_vector(   0 downto 0);
        signal oVar2S53: std_logic_vector(   0 downto 0);
        signal oVar2S54: std_logic_vector(   0 downto 0);
        signal oVar2S55: std_logic_vector(   0 downto 0);
        signal oVar2S56: std_logic_vector(   0 downto 0);
        signal oVar2S57: std_logic_vector(   0 downto 0);
        signal oVar2S58: std_logic_vector(   0 downto 0);
        signal oVar2S59: std_logic_vector(   0 downto 0);
        signal oVar2S60: std_logic_vector(   0 downto 0);
        signal oVar2S61: std_logic_vector(   0 downto 0);
        signal oVar2S62: std_logic_vector(   0 downto 0);
        signal oVar2S64: std_logic_vector(   0 downto 0);
        signal oVar2S65: std_logic_vector(   0 downto 0);
        signal oVar2S67: std_logic_vector(   0 downto 0);
        signal oVar2S68: std_logic_vector(   0 downto 0);
        signal oVar2S69: std_logic_vector(   0 downto 0);
        signal oVar2S70: std_logic_vector(   0 downto 0);
        signal oVar2S71: std_logic_vector(   0 downto 0);
        signal oVar2S72: std_logic_vector(   0 downto 0);
        signal oVar2S73: std_logic_vector(   0 downto 0);
        signal oVar2S74: std_logic_vector(   0 downto 0);
        signal oVar2S75: std_logic_vector(   0 downto 0);
        signal oVar2S76: std_logic_vector(   0 downto 0);
        signal oVar2S77: std_logic_vector(   0 downto 0);
        signal oVar2S78: std_logic_vector(   0 downto 0);
        signal oVar2S79: std_logic_vector(   0 downto 0);
        signal oVar2S80: std_logic_vector(   0 downto 0);
        signal oVar2S82: std_logic_vector(   0 downto 0);
        signal oVar2S83: std_logic_vector(   0 downto 0);
        signal oVar2S85: std_logic_vector(   0 downto 0);
        signal oVar2S86: std_logic_vector(   0 downto 0);
        signal oVar2S87: std_logic_vector(   0 downto 0);
        signal oVar2S88: std_logic_vector(   0 downto 0);
        signal oVar2S89: std_logic_vector(   0 downto 0);
        signal oVar2S90: std_logic_vector(   0 downto 0);
        signal oVar2S91: std_logic_vector(   0 downto 0);
        signal oVar2S92: std_logic_vector(   0 downto 0);
        signal oVar2S94: std_logic_vector(   0 downto 0);
        signal oVar2S95: std_logic_vector(   0 downto 0);
        signal oVar2S97: std_logic_vector(   0 downto 0);
        signal oVar2S98: std_logic_vector(   0 downto 0);
        signal oVar2S100: std_logic_vector(   0 downto 0);
        signal oVar2S101: std_logic_vector(   0 downto 0);
        signal oVar2S103: std_logic_vector(   0 downto 0);
        signal oVar2S104: std_logic_vector(   0 downto 0);
        signal oVar2S106: std_logic_vector(   0 downto 0);
        signal oVar2S107: std_logic_vector(   0 downto 0);
        signal oVar2S108: std_logic_vector(   0 downto 0);
        signal oVar2S109: std_logic_vector(   0 downto 0);
        signal oVar2S110: std_logic_vector(   0 downto 0);
        signal oVar2S111: std_logic_vector(   0 downto 0);
        signal oVar2S112: std_logic_vector(   0 downto 0);
        signal oVar2S113: std_logic_vector(   0 downto 0);
        signal oVar2S114: std_logic_vector(   0 downto 0);
        signal oVar2S115: std_logic_vector(   0 downto 0);
        signal oVar2S116: std_logic_vector(   0 downto 0);
        signal oVar2S117: std_logic_vector(   0 downto 0);
        signal oVar2S119: std_logic_vector(   0 downto 0);
        signal oVar2S120: std_logic_vector(   0 downto 0);
        signal oVar2S121: std_logic_vector(   0 downto 0);
        signal oVar2S122: std_logic_vector(   0 downto 0);
        signal oVar2S123: std_logic_vector(   0 downto 0);
        signal oVar2S124: std_logic_vector(   0 downto 0);
        signal oVar2S125: std_logic_vector(   0 downto 0);
        signal oVar2S126: std_logic_vector(   0 downto 0);
        signal oVar2S128: std_logic_vector(   0 downto 0);
        signal oVar2S129: std_logic_vector(   0 downto 0);
        signal oVar2S130: std_logic_vector(   0 downto 0);
        signal oVar2S131: std_logic_vector(   0 downto 0);
        signal oVar2S132: std_logic_vector(   0 downto 0);
        signal oVar2S133: std_logic_vector(   0 downto 0);
        signal oVar2S134: std_logic_vector(   0 downto 0);
        signal oVar2S135: std_logic_vector(   0 downto 0);
        signal oVar2S136: std_logic_vector(   0 downto 0);
        signal oVar2S137: std_logic_vector(   0 downto 0);
        signal oVar2S138: std_logic_vector(   0 downto 0);
        signal oVar2S139: std_logic_vector(   0 downto 0);
        signal oVar2S140: std_logic_vector(   0 downto 0);
        signal oVar2S141: std_logic_vector(   0 downto 0);
        signal oVar2S142: std_logic_vector(   0 downto 0);
        signal oVar2S143: std_logic_vector(   0 downto 0);
        signal oVar2S144: std_logic_vector(   0 downto 0);
        signal oVar2S145: std_logic_vector(   0 downto 0);
        signal oVar2S146: std_logic_vector(   0 downto 0);
        signal oVar2S147: std_logic_vector(   0 downto 0);
        signal oVar2S148: std_logic_vector(   0 downto 0);
        signal oVar2S149: std_logic_vector(   0 downto 0);
        signal oVar2S150: std_logic_vector(   0 downto 0);
        signal oVar2S151: std_logic_vector(   0 downto 0);
        signal oVar2S152: std_logic_vector(   0 downto 0);
        signal oVar2S153: std_logic_vector(   0 downto 0);
        signal oVar2S154: std_logic_vector(   0 downto 0);
        signal oVar2S155: std_logic_vector(   0 downto 0);
        signal oVar2S156: std_logic_vector(   0 downto 0);
        signal oVar2S157: std_logic_vector(   0 downto 0);
        signal oVar2S158: std_logic_vector(   0 downto 0);
        signal oVar2S159: std_logic_vector(   0 downto 0);
        signal oVar2S160: std_logic_vector(   0 downto 0);
        signal oVar2S162: std_logic_vector(   0 downto 0);
        signal oVar2S163: std_logic_vector(   0 downto 0);
        signal oVar2S165: std_logic_vector(   0 downto 0);
        signal oVar2S166: std_logic_vector(   0 downto 0);
        signal oVar2S168: std_logic_vector(   0 downto 0);
        signal oVar2S169: std_logic_vector(   0 downto 0);
        signal oVar2S170: std_logic_vector(   0 downto 0);
        signal oVar2S171: std_logic_vector(   0 downto 0);
        signal oVar2S173: std_logic_vector(   0 downto 0);
        signal oVar2S174: std_logic_vector(   0 downto 0);
        signal oVar2S176: std_logic_vector(   0 downto 0);
        signal oVar2S177: std_logic_vector(   0 downto 0);
        signal oVar2S179: std_logic_vector(   0 downto 0);
        signal oVar2S180: std_logic_vector(   0 downto 0);
        signal oVar2S182: std_logic_vector(   0 downto 0);
        signal oVar2S183: std_logic_vector(   0 downto 0);
        signal oVar2S184: std_logic_vector(   0 downto 0);
        signal oVar2S185: std_logic_vector(   0 downto 0);
        signal oVar2S187: std_logic_vector(   0 downto 0);
        signal oVar2S188: std_logic_vector(   0 downto 0);
        signal oVar2S190: std_logic_vector(   0 downto 0);
        signal oVar2S191: std_logic_vector(   0 downto 0);
        signal oVar2S193: std_logic_vector(   0 downto 0);
        signal oVar2S194: std_logic_vector(   0 downto 0);
        signal oVar2S195: std_logic_vector(   0 downto 0);
        signal oVar2S196: std_logic_vector(   0 downto 0);
        signal oVar2S197: std_logic_vector(   0 downto 0);
        signal oVar2S198: std_logic_vector(   0 downto 0);
        signal oVar2S199: std_logic_vector(   0 downto 0);
        signal oVar2S200: std_logic_vector(   0 downto 0);
        signal oVar2S201: std_logic_vector(   0 downto 0);
        signal oVar2S202: std_logic_vector(   0 downto 0);
        signal oVar2S204: std_logic_vector(   0 downto 0);
        signal oVar2S205: std_logic_vector(   0 downto 0);
        signal oVar2S206: std_logic_vector(   0 downto 0);
        signal oVar2S207: std_logic_vector(   0 downto 0);
        signal oVar2S208: std_logic_vector(   0 downto 0);
        signal oVar2S209: std_logic_vector(   0 downto 0);
        signal oVar2S211: std_logic_vector(   0 downto 0);
        signal oVar2S212: std_logic_vector(   0 downto 0);
        signal oVar2S213: std_logic_vector(   0 downto 0);
        signal oVar2S214: std_logic_vector(   0 downto 0);
        signal oVar2S216: std_logic_vector(   0 downto 0);
        signal oVar2S217: std_logic_vector(   0 downto 0);
        signal oVar2S218: std_logic_vector(   0 downto 0);
        signal oVar2S219: std_logic_vector(   0 downto 0);
        signal oVar2S220: std_logic_vector(   0 downto 0);
        signal oVar2S221: std_logic_vector(   0 downto 0);
        signal oVar2S222: std_logic_vector(   0 downto 0);
        signal oVar2S223: std_logic_vector(   0 downto 0);
        signal oVar2S225: std_logic_vector(   0 downto 0);
        signal oVar2S226: std_logic_vector(   0 downto 0);
        signal oVar2S227: std_logic_vector(   0 downto 0);
        signal oVar2S228: std_logic_vector(   0 downto 0);
        signal oVar2S230: std_logic_vector(   0 downto 0);
        signal oVar2S231: std_logic_vector(   0 downto 0);
        signal oVar2S232: std_logic_vector(   0 downto 0);
        signal oVar2S233: std_logic_vector(   0 downto 0);
        signal oVar2S234: std_logic_vector(   0 downto 0);
        signal oVar2S235: std_logic_vector(   0 downto 0);
        signal oVar2S237: std_logic_vector(   0 downto 0);
        signal oVar2S238: std_logic_vector(   0 downto 0);
        signal oVar2S240: std_logic_vector(   0 downto 0);
        signal oVar2S241: std_logic_vector(   0 downto 0);
        signal oVar2S243: std_logic_vector(   0 downto 0);
        signal oVar2S244: std_logic_vector(   0 downto 0);
        signal oVar2S246: std_logic_vector(   0 downto 0);
        signal oVar2S247: std_logic_vector(   0 downto 0);
        signal oVar2S249: std_logic_vector(   0 downto 0);
        signal oVar2S250: std_logic_vector(   0 downto 0);
        signal oVar2S251: std_logic_vector(   0 downto 0);
        signal oVar2S252: std_logic_vector(   0 downto 0);
        signal oVar2S253: std_logic_vector(   0 downto 0);
        signal oVar2S254: std_logic_vector(   0 downto 0);
        signal oVar2S255: std_logic_vector(   0 downto 0);
        signal oVar2S256: std_logic_vector(   0 downto 0);
        signal oVar2S257: std_logic_vector(   0 downto 0);
        signal oVar2S258: std_logic_vector(   0 downto 0);
        signal oVar2S259: std_logic_vector(   0 downto 0);
        signal oVar2S260: std_logic_vector(   0 downto 0);
        signal oVar2S261: std_logic_vector(   0 downto 0);
        signal oVar2S262: std_logic_vector(   0 downto 0);
        signal oVar2S263: std_logic_vector(   0 downto 0);
        signal oVar2S264: std_logic_vector(   0 downto 0);
        signal oVar2S266: std_logic_vector(   0 downto 0);
        signal oVar2S267: std_logic_vector(   0 downto 0);
        signal oVar2S268: std_logic_vector(   0 downto 0);
        signal oVar2S269: std_logic_vector(   0 downto 0);
        signal oVar2S270: std_logic_vector(   0 downto 0);
        signal oVar2S271: std_logic_vector(   0 downto 0);
        signal oVar2S272: std_logic_vector(   0 downto 0);
        signal oVar2S274: std_logic_vector(   0 downto 0);
        signal oVar2S275: std_logic_vector(   0 downto 0);
        signal oVar2S277: std_logic_vector(   0 downto 0);
        signal oVar2S278: std_logic_vector(   0 downto 0);
        signal oVar2S279: std_logic_vector(   0 downto 0);
        signal oVar2S280: std_logic_vector(   0 downto 0);
        signal oVar2S282: std_logic_vector(   0 downto 0);
        signal oVar2S283: std_logic_vector(   0 downto 0);
        signal oVar2S285: std_logic_vector(   0 downto 0);
        signal oVar2S286: std_logic_vector(   0 downto 0);
        signal oVar2S287: std_logic_vector(   0 downto 0);
        signal oVar2S288: std_logic_vector(   0 downto 0);
        signal oVar2S289: std_logic_vector(   0 downto 0);
        signal oVar2S290: std_logic_vector(   0 downto 0);
        signal oVar2S291: std_logic_vector(   0 downto 0);
        signal oVar2S292: std_logic_vector(   0 downto 0);
        signal oVar2S293: std_logic_vector(   0 downto 0);
        signal oVar2S294: std_logic_vector(   0 downto 0);
        signal oVar2S295: std_logic_vector(   0 downto 0);
        signal oVar2S296: std_logic_vector(   0 downto 0);
        signal oVar2S298: std_logic_vector(   0 downto 0);
        signal oVar2S299: std_logic_vector(   0 downto 0);
        signal oVar2S300: std_logic_vector(   0 downto 0);
        signal oVar2S301: std_logic_vector(   0 downto 0);
        signal oVar2S302: std_logic_vector(   0 downto 0);
        signal oVar2S304: std_logic_vector(   0 downto 0);
        signal oVar2S305: std_logic_vector(   0 downto 0);
        signal oVar2S306: std_logic_vector(   0 downto 0);
        signal oVar2S307: std_logic_vector(   0 downto 0);
        signal oVar3S0: std_logic_vector(   0 downto 0);
        signal oVar3S1: std_logic_vector(   0 downto 0);
        signal oVar3S2: std_logic_vector(   0 downto 0);
        signal oVar3S3: std_logic_vector(   0 downto 0);
        signal oVar3S4: std_logic_vector(   0 downto 0);
        signal oVar3S5: std_logic_vector(   0 downto 0);
        signal oVar3S6: std_logic_vector(   0 downto 0);
        signal oVar3S7: std_logic_vector(   0 downto 0);
        signal oVar3S8: std_logic_vector(   0 downto 0);
        signal oVar3S9: std_logic_vector(   0 downto 0);
        signal oVar3S10: std_logic_vector(   0 downto 0);
        signal oVar3S11: std_logic_vector(   0 downto 0);
        signal oVar3S12: std_logic_vector(   0 downto 0);
        signal oVar3S13: std_logic_vector(   0 downto 0);
        signal oVar3S14: std_logic_vector(   0 downto 0);
        signal oVar3S15: std_logic_vector(   0 downto 0);
        signal oVar3S16: std_logic_vector(   0 downto 0);
        signal oVar3S17: std_logic_vector(   0 downto 0);
        signal oVar3S18: std_logic_vector(   0 downto 0);
        signal oVar3S19: std_logic_vector(   0 downto 0);
        signal oVar3S20: std_logic_vector(   0 downto 0);
        signal oVar3S21: std_logic_vector(   0 downto 0);
        signal oVar3S22: std_logic_vector(   0 downto 0);
        signal oVar3S23: std_logic_vector(   0 downto 0);
        signal oVar3S24: std_logic_vector(   0 downto 0);
        signal oVar3S25: std_logic_vector(   0 downto 0);
        signal oVar3S26: std_logic_vector(   0 downto 0);
        signal oVar3S27: std_logic_vector(   0 downto 0);
        signal oVar3S28: std_logic_vector(   0 downto 0);
        signal oVar3S29: std_logic_vector(   0 downto 0);
        signal oVar3S30: std_logic_vector(   0 downto 0);
        signal oVar3S31: std_logic_vector(   0 downto 0);
        signal oVar3S32: std_logic_vector(   0 downto 0);
        signal oVar3S33: std_logic_vector(   0 downto 0);
        signal oVar3S34: std_logic_vector(   0 downto 0);
        signal oVar3S35: std_logic_vector(   0 downto 0);
        signal oVar3S36: std_logic_vector(   0 downto 0);
        signal oVar3S37: std_logic_vector(   0 downto 0);
        signal oVar3S38: std_logic_vector(   0 downto 0);
        signal oVar3S39: std_logic_vector(   0 downto 0);
        signal oVar3S40: std_logic_vector(   0 downto 0);
        signal oVar3S41: std_logic_vector(   0 downto 0);
        signal oVar3S42: std_logic_vector(   0 downto 0);
        signal oVar3S43: std_logic_vector(   0 downto 0);
        signal oVar3S44: std_logic_vector(   0 downto 0);
        signal oVar3S45: std_logic_vector(   0 downto 0);
        signal oVar3S46: std_logic_vector(   0 downto 0);
        signal oVar3S47: std_logic_vector(   0 downto 0);
        signal oVar3S48: std_logic_vector(   0 downto 0);
        signal oVar3S49: std_logic_vector(   0 downto 0);
        signal oVar3S50: std_logic_vector(   0 downto 0);
        signal oVar3S51: std_logic_vector(   0 downto 0);
        signal oVar3S52: std_logic_vector(   0 downto 0);
        signal oVar3S53: std_logic_vector(   0 downto 0);
        signal oVar3S54: std_logic_vector(   0 downto 0);
        signal oVar3S55: std_logic_vector(   0 downto 0);
        signal oVar3S56: std_logic_vector(   0 downto 0);
        signal oVar3S57: std_logic_vector(   0 downto 0);
        signal oVar3S58: std_logic_vector(   0 downto 0);
        signal oVar3S59: std_logic_vector(   0 downto 0);
        signal oVar3S60: std_logic_vector(   0 downto 0);
        signal oVar3S61: std_logic_vector(   0 downto 0);
        signal oVar3S62: std_logic_vector(   0 downto 0);
        signal oVar3S63: std_logic_vector(   0 downto 0);
        signal oVar3S64: std_logic_vector(   0 downto 0);
        signal oVar3S65: std_logic_vector(   0 downto 0);
        signal oVar3S66: std_logic_vector(   0 downto 0);
        signal oVar3S67: std_logic_vector(   0 downto 0);
        signal oVar3S68: std_logic_vector(   0 downto 0);
        signal oVar3S69: std_logic_vector(   0 downto 0);
        signal oVar3S70: std_logic_vector(   0 downto 0);
        signal oVar3S71: std_logic_vector(   0 downto 0);
        signal oVar3S72: std_logic_vector(   0 downto 0);
        signal oVar3S73: std_logic_vector(   0 downto 0);
        signal oVar3S74: std_logic_vector(   0 downto 0);
        signal oVar3S75: std_logic_vector(   0 downto 0);
        signal oVar3S76: std_logic_vector(   0 downto 0);
        signal oVar3S77: std_logic_vector(   0 downto 0);
        signal oVar3S78: std_logic_vector(   0 downto 0);
        signal oVar3S79: std_logic_vector(   0 downto 0);
        signal oVar3S80: std_logic_vector(   0 downto 0);
        signal oVar3S81: std_logic_vector(   0 downto 0);
        signal oVar3S82: std_logic_vector(   0 downto 0);
        signal oVar3S83: std_logic_vector(   0 downto 0);
        signal oVar3S84: std_logic_vector(   0 downto 0);
        signal oVar3S85: std_logic_vector(   0 downto 0);
        signal oVar3S86: std_logic_vector(   0 downto 0);
        signal oVar3S87: std_logic_vector(   0 downto 0);
        signal oVar3S88: std_logic_vector(   0 downto 0);
        signal oVar3S89: std_logic_vector(   0 downto 0);
        signal oVar3S90: std_logic_vector(   0 downto 0);
        signal oVar3S91: std_logic_vector(   0 downto 0);
        signal oVar3S92: std_logic_vector(   0 downto 0);
        signal oVar3S93: std_logic_vector(   0 downto 0);
        signal oVar3S94: std_logic_vector(   0 downto 0);
        signal oVar3S95: std_logic_vector(   0 downto 0);
        signal oVar3S96: std_logic_vector(   0 downto 0);
        signal oVar3S97: std_logic_vector(   0 downto 0);
        signal oVar3S98: std_logic_vector(   0 downto 0);
        signal oVar3S99: std_logic_vector(   0 downto 0);
        signal oVar3S100: std_logic_vector(   0 downto 0);
        signal oVar3S101: std_logic_vector(   0 downto 0);
        signal oVar3S102: std_logic_vector(   0 downto 0);
        signal oVar3S103: std_logic_vector(   0 downto 0);
        signal oVar3S104: std_logic_vector(   0 downto 0);
        signal oVar3S105: std_logic_vector(   0 downto 0);
        signal oVar3S106: std_logic_vector(   0 downto 0);
        signal oVar3S107: std_logic_vector(   0 downto 0);
        signal oVar3S108: std_logic_vector(   0 downto 0);
        signal oVar3S109: std_logic_vector(   0 downto 0);
        signal oVar3S110: std_logic_vector(   0 downto 0);
        signal oVar3S111: std_logic_vector(   0 downto 0);
        signal oVar3S112: std_logic_vector(   0 downto 0);
        signal oVar3S113: std_logic_vector(   0 downto 0);
        signal oVar3S114: std_logic_vector(   0 downto 0);
        signal oVar3S115: std_logic_vector(   0 downto 0);
        signal oVar3S116: std_logic_vector(   0 downto 0);
        signal oVar3S117: std_logic_vector(   0 downto 0);
        signal oVar3S118: std_logic_vector(   0 downto 0);
        signal oVar3S119: std_logic_vector(   0 downto 0);
        signal oVar3S120: std_logic_vector(   0 downto 0);
        signal oVar3S121: std_logic_vector(   0 downto 0);
        signal oVar3S122: std_logic_vector(   0 downto 0);
        signal oVar3S123: std_logic_vector(   0 downto 0);
        signal oVar3S124: std_logic_vector(   0 downto 0);
        signal oVar3S125: std_logic_vector(   0 downto 0);
        signal oVar3S126: std_logic_vector(   0 downto 0);
        signal oVar3S127: std_logic_vector(   0 downto 0);
        signal aVar3S0: std_logic_vector(   15 downto 0);
        signal aVar3S1: std_logic_vector(   15 downto 0);
        signal aVar3S2: std_logic_vector(   15 downto 0);
        signal aVar3S3: std_logic_vector(   15 downto 0);
        signal aVar3S4: std_logic_vector(   15 downto 0);
        signal aVar3S5: std_logic_vector(   15 downto 0);
        signal aVar3S6: std_logic_vector(   15 downto 0);
        signal aVar3S7: std_logic_vector(   15 downto 0);
        signal aVar3S8: std_logic_vector(   15 downto 0);
        signal aVar3S9: std_logic_vector(   15 downto 0);
        signal aVar3S10: std_logic_vector(   15 downto 0);
        signal aVar3S11: std_logic_vector(   15 downto 0);
        signal aVar3S12: std_logic_vector(   15 downto 0);
        signal aVar3S13: std_logic_vector(   15 downto 0);
        signal aVar3S14: std_logic_vector(   15 downto 0);
        signal aVar3S15: std_logic_vector(   15 downto 0);
        signal aVar4S0: std_logic_vector(   15 downto 0);
        signal aVar4S1: std_logic_vector(   15 downto 0);
        signal aVar4S2: std_logic_vector(   15 downto 0);
        signal aVar4S3: std_logic_vector(   15 downto 0);
        signal aVar4S4: std_logic_vector(   15 downto 0);
        signal aVar4S5: std_logic_vector(   15 downto 0);
        signal aVar4S6: std_logic_vector(   15 downto 0);
        signal aVar4S7: std_logic_vector(   15 downto 0);
        signal aVar5S0: std_logic_vector(   15 downto 0);
        signal aVar5S1: std_logic_vector(   15 downto 0);
        signal aVar5S2: std_logic_vector(   15 downto 0);
        signal aVar5S3: std_logic_vector(   15 downto 0);
        signal aVar6S0: std_logic_vector(   15 downto 0);
        signal aVar6S1: std_logic_vector(   15 downto 0);
        signal aVar7S0: std_logic_vector(   15 downto 0);
signal ADDM4K3S1: std_logic_vector(   7 downto 0);
signal ADDM4K3S0: std_logic_vector(   7 downto 0);
signal ADDM4K3S3: std_logic_vector(   7 downto 0);
signal ADDM4K3S2: std_logic_vector(   7 downto 0);
signal ADDM4K3S5: std_logic_vector(   7 downto 0);
signal ADDM4K3S4: std_logic_vector(   7 downto 0);
signal ADDM4K3S7: std_logic_vector(   7 downto 0);
signal ADDM4K3S6: std_logic_vector(   7 downto 0);
signal ADDM4K3S9: std_logic_vector(   7 downto 0);
signal ADDM4K3S8: std_logic_vector(   7 downto 0);
signal ADDM4K3S11: std_logic_vector(   7 downto 0);
signal ADDM4K3S10: std_logic_vector(   7 downto 0);
signal ADDM4K3S13: std_logic_vector(   7 downto 0);
signal ADDM4K3S12: std_logic_vector(   7 downto 0);
signal ADDM4K3S15: std_logic_vector(   7 downto 0);
signal ADDM4K3S14: std_logic_vector(   7 downto 0);
BEGIN
	A (19 downto 0) <= A_DIN_L (19 downto 0);
	B (8 downto 0) <= A_DIN_L (28 downto 20);
	B (17 downto 9) <= B_DIN_L (8 downto 0);
	D (15 downto 0) <= B_DIN_L (24 downto 9);
	E (15 downto 0) <= D_DIN_L (31 downto 16);
	C_DOUT_L (15 downto 0) <= output (15 downto 0);
lookuptable_LV1 : process(c1)
begin
 if c1'event and c1='1' then
        if(E(12)='1' AND B(14)='1' )then
          cVar1S0S0P055P030nsss(0) <='1';
          else
          cVar1S0S0P055P030nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B( 4)='1' )then
          cVar1S1S0P055N030P031nsss(0) <='1';
          else
          cVar1S1S0P055N030P031nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B( 4)='0' AND B(15)='1' )then
          cVar1S2S0P055N030N031P028nsss(0) <='1';
          else
          cVar1S2S0P055N030N031P028nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B( 4)='0' AND B(15)='0' )then
          cVar1S3S0P055N030N031N028(0) <='1';
          else
          cVar1S3S0P055N030N031N028(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B( 4)='0' AND B(15)='0' )then
          cVar1S4S0P055N030N031N028(0) <='1';
          else
          cVar1S4S0P055N030N031N028(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B( 4)='0' AND B(15)='0' )then
          cVar1S5S0P055N030N031N028(0) <='1';
          else
          cVar1S5S0P055N030N031N028(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='1' AND B(13)='1' )then
          cVar1S6S0N055P059P061P032nsss(0) <='1';
          else
          cVar1S6S0N055P059P061P032nsss(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='1' AND B(13)='0' )then
          cVar1S7S0N055P059P061N032(0) <='1';
          else
          cVar1S7S0N055P059P061N032(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='1' AND B(13)='0' )then
          cVar1S8S0N055P059P061N032(0) <='1';
          else
          cVar1S8S0N055P059P061N032(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='1' AND B(13)='0' )then
          cVar1S9S0N055P059P061N032(0) <='1';
          else
          cVar1S9S0N055P059P061N032(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='0' AND E( 3)='1' )then
          cVar1S10S0N055P059N061P058nsss(0) <='1';
          else
          cVar1S10S0N055P059N061P058nsss(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='0' AND E( 3)='0' )then
          cVar1S11S0N055P059N061N058(0) <='1';
          else
          cVar1S11S0N055P059N061N058(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='0' AND E( 3)='0' )then
          cVar1S12S0N055P059N061N058(0) <='1';
          else
          cVar1S12S0N055P059N061N058(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='1' AND D(10)='0' AND E( 3)='0' )then
          cVar1S13S0N055P059N061N058(0) <='1';
          else
          cVar1S13S0N055P059N061N058(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='1' AND B( 5)='1' )then
          cVar1S14S0N055N059P052P029nsss(0) <='1';
          else
          cVar1S14S0N055N059P052P029nsss(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S15S0N055N059P052N029(0) <='1';
          else
          cVar1S15S0N055N059P052N029(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S16S0N055N059P052N029(0) <='1';
          else
          cVar1S16S0N055N059P052N029(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S17S0N055N059P052N029(0) <='1';
          else
          cVar1S17S0N055N059P052N029(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='1' )then
          cVar1S18S0N055N059N052P047(0) <='1';
          else
          cVar1S18S0N055N059N052P047(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='1' )then
          cVar1S19S0N055N059N052P047(0) <='1';
          else
          cVar1S19S0N055N059N052P047(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='1' )then
          cVar1S20S0N055N059N052P047(0) <='1';
          else
          cVar1S20S0N055N059N052P047(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='0' )then
          cVar1S21S0N055N059N052N047(0) <='1';
          else
          cVar1S21S0N055N059N052N047(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='0' )then
          cVar1S22S0N055N059N052N047(0) <='1';
          else
          cVar1S22S0N055N059N052N047(0) <='0';
          end if;
        if(E(12)='0' AND E(11)='0' AND D( 4)='0' AND E(14)='0' )then
          cVar1S23S0N055N059N052N047(0) <='1';
          else
          cVar1S23S0N055N059N052N047(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='1' AND D( 2)='1' )then
          cVar1S0S1P058P033P060nsss(0) <='1';
          else
          cVar1S0S1P058P033P060nsss(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='1' AND D( 2)='0' AND A(10)='0' )then
          cVar1S1S1P058P033N060P018(0) <='1';
          else
          cVar1S1S1P058P033N060P018(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='1' AND D( 2)='0' AND A(10)='0' )then
          cVar1S2S1P058P033N060P018(0) <='1';
          else
          cVar1S2S1P058P033N060P018(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='0' AND B( 4)='1' )then
          cVar1S3S1P058N033P031nsss(0) <='1';
          else
          cVar1S3S1P058N033P031nsss(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='0' AND B( 4)='0' AND B(13)='1' )then
          cVar1S4S1P058N033N031P032nsss(0) <='1';
          else
          cVar1S4S1P058N033N031P032nsss(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S5S1P058N033N031N032(0) <='1';
          else
          cVar1S5S1P058N033N031N032(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S6S1P058N033N031N032(0) <='1';
          else
          cVar1S6S1P058N033N031N032(0) <='0';
          end if;
        if(E( 3)='1' AND B( 3)='0' AND B( 4)='0' AND B(13)='0' )then
          cVar1S7S1P058N033N031N032(0) <='1';
          else
          cVar1S7S1P058N033N031N032(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='1' AND B(15)='1' )then
          cVar1S8S1N058P051P053P028nsss(0) <='1';
          else
          cVar1S8S1N058P051P053P028nsss(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='1' AND B(15)='0' )then
          cVar1S9S1N058P051P053N028(0) <='1';
          else
          cVar1S9S1N058P051P053N028(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='1' AND B(15)='0' )then
          cVar1S10S1N058P051P053N028(0) <='1';
          else
          cVar1S10S1N058P051P053N028(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='1' AND B(15)='0' )then
          cVar1S11S1N058P051P053N028(0) <='1';
          else
          cVar1S11S1N058P051P053N028(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='0' AND B(16)='1' )then
          cVar1S12S1N058P051N053P026nsss(0) <='1';
          else
          cVar1S12S1N058P051N053P026nsss(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='0' AND B(16)='0' )then
          cVar1S13S1N058P051N053N026(0) <='1';
          else
          cVar1S13S1N058P051N053N026(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='0' AND B(16)='0' )then
          cVar1S14S1N058P051N053N026(0) <='1';
          else
          cVar1S14S1N058P051N053N026(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='1' AND D(12)='0' AND B(16)='0' )then
          cVar1S15S1N058P051N053N026(0) <='1';
          else
          cVar1S15S1N058P051N053N026(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='1' AND B( 7)='1' )then
          cVar1S16S1N058N051P046P025nsss(0) <='1';
          else
          cVar1S16S1N058N051P046P025nsss(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S17S1N058N051P046N025(0) <='1';
          else
          cVar1S17S1N058N051P046N025(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S18S1N058N051P046N025(0) <='1';
          else
          cVar1S18S1N058N051P046N025(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='1' AND B( 7)='0' )then
          cVar1S19S1N058N051P046N025(0) <='1';
          else
          cVar1S19S1N058N051P046N025(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='1' )then
          cVar1S20S1N058N051N046P064(0) <='1';
          else
          cVar1S20S1N058N051N046P064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='1' )then
          cVar1S21S1N058N051N046P064(0) <='1';
          else
          cVar1S21S1N058N051N046P064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='1' )then
          cVar1S22S1N058N051N046P064(0) <='1';
          else
          cVar1S22S1N058N051N046P064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='0' )then
          cVar1S23S1N058N051N046N064(0) <='1';
          else
          cVar1S23S1N058N051N046N064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='0' )then
          cVar1S24S1N058N051N046N064(0) <='1';
          else
          cVar1S24S1N058N051N046N064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='0' )then
          cVar1S25S1N058N051N046N064(0) <='1';
          else
          cVar1S25S1N058N051N046N064(0) <='0';
          end if;
        if(E( 3)='0' AND E(13)='0' AND E( 6)='0' AND D( 1)='0' )then
          cVar1S26S1N058N051N046N064(0) <='1';
          else
          cVar1S26S1N058N051N046N064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND E( 1)='1' )then
          cVar1S0S2P068P019P015P066nsss(0) <='1';
          else
          cVar1S0S2P068P019P015P066nsss(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND E( 1)='0' )then
          cVar1S1S2P068P019P015N066(0) <='1';
          else
          cVar1S1S2P068P019P015N066(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='0' )then
          cVar1S2S2P068P019P015P064(0) <='1';
          else
          cVar1S2S2P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='0' )then
          cVar1S3S2P068P019P015P064(0) <='1';
          else
          cVar1S3S2P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='1' )then
          cVar1S4S2P068P019P015P064(0) <='1';
          else
          cVar1S4S2P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='0' AND A(10)='1' )then
          cVar1S5S2P068N019P011P018nsss(0) <='1';
          else
          cVar1S5S2P068N019P011P018nsss(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='0' AND A(10)='0' )then
          cVar1S6S2P068N019P011N018(0) <='1';
          else
          cVar1S6S2P068N019P011N018(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='0' AND A(10)='0' )then
          cVar1S7S2P068N019P011N018(0) <='1';
          else
          cVar1S7S2P068N019P011N018(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='1' AND E( 9)='0' )then
          cVar1S8S2P068N019P011P067(0) <='1';
          else
          cVar1S8S2P068N019P011P067(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='1' AND E( 9)='0' )then
          cVar1S9S2P068N019P011P067(0) <='1';
          else
          cVar1S9S2P068N019P011P067(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A( 4)='1' AND E( 9)='1' )then
          cVar1S10S2P068N019P011P067(0) <='1';
          else
          cVar1S10S2P068N019P011P067(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B(10)='1' )then
          cVar1S11S2N068P040P038nsss(0) <='1';
          else
          cVar1S11S2N068P040P038nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B(10)='0' AND B( 8)='1' )then
          cVar1S12S2N068P040N038P023nsss(0) <='1';
          else
          cVar1S12S2N068P040N038P023nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B(10)='0' AND B( 8)='0' )then
          cVar1S13S2N068P040N038N023(0) <='1';
          else
          cVar1S13S2N068P040N038N023(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B(10)='0' AND B( 8)='0' )then
          cVar1S14S2N068P040N038N023(0) <='1';
          else
          cVar1S14S2N068P040N038N023(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B(10)='0' AND B( 8)='0' )then
          cVar1S15S2N068P040N038N023(0) <='1';
          else
          cVar1S15S2N068P040N038N023(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='1' AND B( 6)='1' )then
          cVar1S16S2N068N040P050P027nsss(0) <='1';
          else
          cVar1S16S2N068N040P050P027nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S17S2N068N040P050N027(0) <='1';
          else
          cVar1S17S2N068N040P050N027(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S18S2N068N040P050N027(0) <='1';
          else
          cVar1S18S2N068N040P050N027(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S19S2N068N040P050N027(0) <='1';
          else
          cVar1S19S2N068N040P050N027(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='1' )then
          cVar1S20S2N068N040N050P046(0) <='1';
          else
          cVar1S20S2N068N040N050P046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='1' )then
          cVar1S21S2N068N040N050P046(0) <='1';
          else
          cVar1S21S2N068N040N050P046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S22S2N068N040N050N046(0) <='1';
          else
          cVar1S22S2N068N040N050N046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S23S2N068N040N050N046(0) <='1';
          else
          cVar1S23S2N068N040N050N046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S24S2N068N040N050N046(0) <='1';
          else
          cVar1S24S2N068N040N050N046(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S0S3P068P019P015P017(0) <='1';
          else
          cVar1S0S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S1S3P068P019P015P017(0) <='1';
          else
          cVar1S1S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S2S3P068P019P015P017(0) <='1';
          else
          cVar1S2S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S3S3P068P019P015P017(0) <='1';
          else
          cVar1S3S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S4S3P068P019P015P017(0) <='1';
          else
          cVar1S4S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S5S3P068P019P015P017(0) <='1';
          else
          cVar1S5S3P068P019P015P017(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='0' )then
          cVar1S6S3P068P019P015P064(0) <='1';
          else
          cVar1S6S3P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='0' )then
          cVar1S7S3P068P019P015P064(0) <='1';
          else
          cVar1S7S3P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='1' AND A( 2)='1' AND D( 1)='1' )then
          cVar1S8S3P068P019P015P064(0) <='1';
          else
          cVar1S8S3P068P019P015P064(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='1' AND A( 9)='0' )then
          cVar1S9S3P068N019P018P001(0) <='1';
          else
          cVar1S9S3P068N019P018P001(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='1' AND A( 9)='0' )then
          cVar1S10S3P068N019P018P001(0) <='1';
          else
          cVar1S10S3P068N019P018P001(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='1' AND A( 9)='0' )then
          cVar1S11S3P068N019P018P001(0) <='1';
          else
          cVar1S11S3P068N019P018P001(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='1' AND A( 9)='0' )then
          cVar1S12S3P068N019P018P001(0) <='1';
          else
          cVar1S12S3P068N019P018P001(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='0' )then
          cVar1S13S3P068N019N018P010(0) <='1';
          else
          cVar1S13S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='0' )then
          cVar1S14S3P068N019N018P010(0) <='1';
          else
          cVar1S14S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='0' )then
          cVar1S15S3P068N019N018P010(0) <='1';
          else
          cVar1S15S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='0' )then
          cVar1S16S3P068N019N018P010(0) <='1';
          else
          cVar1S16S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='1' )then
          cVar1S17S3P068N019N018P010(0) <='1';
          else
          cVar1S17S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='1' AND A( 0)='0' AND A(10)='0' AND A(14)='1' )then
          cVar1S18S3P068N019N018P010(0) <='1';
          else
          cVar1S18S3P068N019N018P010(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S19S3N068P040P021nsss(0) <='1';
          else
          cVar1S19S3N068P040P021nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='1' )then
          cVar1S20S3N068P040N021P020nsss(0) <='1';
          else
          cVar1S20S3N068P040N021P020nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S21S3N068P040N021N020(0) <='1';
          else
          cVar1S21S3N068P040N021N020(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S22S3N068P040N021N020(0) <='1';
          else
          cVar1S22S3N068P040N021N020(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S23S3N068P040N021N020(0) <='1';
          else
          cVar1S23S3N068P040N021N020(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='1' )then
          cVar1S24S3N068N040P050nsss(0) <='1';
          else
          cVar1S24S3N068N040P050nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='1' )then
          cVar1S25S3N068N040N050P046nsss(0) <='1';
          else
          cVar1S25S3N068N040N050P046nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S26S3N068N040N050N046(0) <='1';
          else
          cVar1S26S3N068N040N050N046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S27S3N068N040N050N046(0) <='1';
          else
          cVar1S27S3N068N040N050N046(0) <='0';
          end if;
        if(D( 0)='0' AND D( 7)='0' AND E( 5)='0' AND E( 6)='0' )then
          cVar1S28S3N068N040N050N046(0) <='1';
          else
          cVar1S28S3N068N040N050N046(0) <='0';
          end if;
        if(D( 7)='1' AND B(10)='1' )then
          cVar1S0S4P040P038nsss(0) <='1';
          else
          cVar1S0S4P040P038nsss(0) <='0';
          end if;
        if(D( 7)='1' AND B(10)='0' AND E( 9)='0' AND B( 8)='1' )then
          cVar1S1S4P040N038P067P023nsss(0) <='1';
          else
          cVar1S1S4P040N038P067P023nsss(0) <='0';
          end if;
        if(D( 7)='1' AND B(10)='0' AND E( 9)='0' AND B( 8)='0' )then
          cVar1S2S4P040N038P067N023(0) <='1';
          else
          cVar1S2S4P040N038P067N023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S3S4N040P044P023nsss(0) <='1';
          else
          cVar1S3S4N040P044P023nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND B( 8)='0' AND B(18)='1' )then
          cVar1S4S4N040P044N023P022nsss(0) <='1';
          else
          cVar1S4S4N040P044N023P022nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND B( 8)='0' AND B(18)='0' )then
          cVar1S5S4N040P044N023N022(0) <='1';
          else
          cVar1S5S4N040P044N023N022(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND B( 8)='0' AND B(18)='0' )then
          cVar1S6S4N040P044N023N022(0) <='1';
          else
          cVar1S6S4N040P044N023N022(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND B( 8)='0' AND B(18)='0' )then
          cVar1S7S4N040P044N023N022(0) <='1';
          else
          cVar1S7S4N040P044N023N022(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='1' AND B(17)='1' )then
          cVar1S8S4N040N044P047P024nsss(0) <='1';
          else
          cVar1S8S4N040N044P047P024nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='1' AND B(17)='0' )then
          cVar1S9S4N040N044P047N024(0) <='1';
          else
          cVar1S9S4N040N044P047N024(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='1' AND B(17)='0' )then
          cVar1S10S4N040N044P047N024(0) <='1';
          else
          cVar1S10S4N040N044P047N024(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='1' AND B(17)='0' )then
          cVar1S11S4N040N044P047N024(0) <='1';
          else
          cVar1S11S4N040N044P047N024(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='1' )then
          cVar1S12S4N040N044N047P061(0) <='1';
          else
          cVar1S12S4N040N044N047P061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='1' )then
          cVar1S13S4N040N044N047P061(0) <='1';
          else
          cVar1S13S4N040N044N047P061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='1' )then
          cVar1S14S4N040N044N047P061(0) <='1';
          else
          cVar1S14S4N040N044N047P061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='1' )then
          cVar1S15S4N040N044N047P061(0) <='1';
          else
          cVar1S15S4N040N044N047P061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='0' )then
          cVar1S16S4N040N044N047N061(0) <='1';
          else
          cVar1S16S4N040N044N047N061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='0' )then
          cVar1S17S4N040N044N047N061(0) <='1';
          else
          cVar1S17S4N040N044N047N061(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E(14)='0' AND D(10)='0' )then
          cVar1S18S4N040N044N047N061(0) <='1';
          else
          cVar1S18S4N040N044N047N061(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' )then
          cVar1S0S5P044P023nsss(0) <='1';
          else
          cVar1S0S5P044P023nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='1' )then
          cVar1S1S5P044N023P022nsss(0) <='1';
          else
          cVar1S1S5P044N023P022nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='1' )then
          cVar1S2S5P044N023N022P025nsss(0) <='1';
          else
          cVar1S2S5P044N023N022P025nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='0' )then
          cVar1S3S5P044N023N022N025(0) <='1';
          else
          cVar1S3S5P044N023N022N025(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='0' )then
          cVar1S4S5P044N023N022N025(0) <='1';
          else
          cVar1S4S5P044N023N022N025(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S5S5N044P040P021nsss(0) <='1';
          else
          cVar1S5S5N044P040P021nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='1' )then
          cVar1S6S5N044P040N021P020nsss(0) <='1';
          else
          cVar1S6S5N044P040N021P020nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S7S5N044P040N021N020(0) <='1';
          else
          cVar1S7S5N044P040N021N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S8S5N044P040N021N020(0) <='1';
          else
          cVar1S8S5N044P040N021N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S9S5N044P040N021N020(0) <='1';
          else
          cVar1S9S5N044P040N021N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='1' AND A(16)='1' )then
          cVar1S10S5N044N040P047P006nsss(0) <='1';
          else
          cVar1S10S5N044N040P047P006nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='1' AND A(16)='0' )then
          cVar1S11S5N044N040P047N006(0) <='1';
          else
          cVar1S11S5N044N040P047N006(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='1' AND A(16)='0' )then
          cVar1S12S5N044N040P047N006(0) <='1';
          else
          cVar1S12S5N044N040P047N006(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='1' )then
          cVar1S13S5N044N040N047P056(0) <='1';
          else
          cVar1S13S5N044N040N047P056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='1' )then
          cVar1S14S5N044N040N047P056(0) <='1';
          else
          cVar1S14S5N044N040N047P056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='1' )then
          cVar1S15S5N044N040N047P056(0) <='1';
          else
          cVar1S15S5N044N040N047P056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='1' )then
          cVar1S16S5N044N040N047P056(0) <='1';
          else
          cVar1S16S5N044N040N047P056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='0' )then
          cVar1S17S5N044N040N047N056(0) <='1';
          else
          cVar1S17S5N044N040N047N056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='0' )then
          cVar1S18S5N044N040N047N056(0) <='1';
          else
          cVar1S18S5N044N040N047N056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='0' )then
          cVar1S19S5N044N040N047N056(0) <='1';
          else
          cVar1S19S5N044N040N047N056(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND E(14)='0' AND D( 3)='0' )then
          cVar1S20S5N044N040N047N056(0) <='1';
          else
          cVar1S20S5N044N040N047N056(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' )then
          cVar1S0S6P044P023nsss(0) <='1';
          else
          cVar1S0S6P044P023nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='1' )then
          cVar1S1S6P044N023P004nsss(0) <='1';
          else
          cVar1S1S6P044N023P004nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S2S6P044N023N004P006nsss(0) <='1';
          else
          cVar1S2S6P044N023N004P006nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S3S6P044N023N004N006(0) <='1';
          else
          cVar1S3S6P044N023N004N006(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S4S6P044N023N004N006(0) <='1';
          else
          cVar1S4S6P044N023N004N006(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='1' AND B( 6)='1' )then
          cVar1S5S6N044P015P050P027nsss(0) <='1';
          else
          cVar1S5S6N044P015P050P027nsss(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S6S6N044P015P050N027(0) <='1';
          else
          cVar1S6S6N044P015P050N027(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S7S6N044P015P050N027(0) <='1';
          else
          cVar1S7S6N044P015P050N027(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S8S6N044P015P050N027(0) <='1';
          else
          cVar1S8S6N044P015P050N027(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='0' AND D( 3)='1' )then
          cVar1S9S6N044P015N050P056(0) <='1';
          else
          cVar1S9S6N044P015N050P056(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='0' AND D( 3)='1' )then
          cVar1S10S6N044P015N050P056(0) <='1';
          else
          cVar1S10S6N044P015N050P056(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='0' AND D( 3)='1' )then
          cVar1S11S6N044P015N050P056(0) <='1';
          else
          cVar1S11S6N044P015N050P056(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S12S6N044P015N050N056(0) <='1';
          else
          cVar1S12S6N044P015N050N056(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='0' AND E( 5)='0' AND D( 3)='0' )then
          cVar1S13S6N044P015N050N056(0) <='1';
          else
          cVar1S13S6N044P015N050N056(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='1' AND B( 2)='1' )then
          cVar1S14S6N044P015P062P035(0) <='1';
          else
          cVar1S14S6N044P015P062P035(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='1' AND B( 2)='1' )then
          cVar1S15S6N044P015P062P035(0) <='1';
          else
          cVar1S15S6N044P015P062P035(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='1' AND B( 2)='1' )then
          cVar1S16S6N044P015P062P035(0) <='1';
          else
          cVar1S16S6N044P015P062P035(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='1' AND B( 2)='0' )then
          cVar1S17S6N044P015P062N035(0) <='1';
          else
          cVar1S17S6N044P015P062N035(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='1' AND B( 2)='0' )then
          cVar1S18S6N044P015P062N035(0) <='1';
          else
          cVar1S18S6N044P015P062N035(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='1' )then
          cVar1S19S6N044P015N062P058(0) <='1';
          else
          cVar1S19S6N044P015N062P058(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='1' )then
          cVar1S20S6N044P015N062P058(0) <='1';
          else
          cVar1S20S6N044P015N062P058(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='0' )then
          cVar1S21S6N044P015N062N058(0) <='1';
          else
          cVar1S21S6N044P015N062N058(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='0' )then
          cVar1S22S6N044P015N062N058(0) <='1';
          else
          cVar1S22S6N044P015N062N058(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='0' )then
          cVar1S23S6N044P015N062N058(0) <='1';
          else
          cVar1S23S6N044P015N062N058(0) <='0';
          end if;
        if(D( 6)='0' AND A( 2)='1' AND E( 2)='0' AND E( 3)='0' )then
          cVar1S24S6N044P015N062N058(0) <='1';
          else
          cVar1S24S6N044P015N062N058(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='1' AND D( 5)='1' )then
          cVar1S0S7P050P027P048nsss(0) <='1';
          else
          cVar1S0S7P050P027P048nsss(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='1' AND D( 5)='0' AND A( 5)='1' )then
          cVar1S1S7P050P027N048P009nsss(0) <='1';
          else
          cVar1S1S7P050P027N048P009nsss(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='1' AND D( 5)='0' AND A( 5)='0' )then
          cVar1S2S7P050P027N048N009(0) <='1';
          else
          cVar1S2S7P050P027N048N009(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='1' AND D( 5)='0' AND A( 5)='0' )then
          cVar1S3S7P050P027N048N009(0) <='1';
          else
          cVar1S3S7P050P027N048N009(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='1' AND A(15)='1' )then
          cVar1S4S7P050N027P052P008nsss(0) <='1';
          else
          cVar1S4S7P050N027P052P008nsss(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S5S7P050N027P052N008(0) <='1';
          else
          cVar1S5S7P050N027P052N008(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S6S7P050N027P052N008(0) <='1';
          else
          cVar1S6S7P050N027P052N008(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='1' AND A(15)='0' )then
          cVar1S7S7P050N027P052N008(0) <='1';
          else
          cVar1S7S7P050N027P052N008(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='0' AND D( 5)='1' )then
          cVar1S8S7P050N027N052P048(0) <='1';
          else
          cVar1S8S7P050N027N052P048(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='0' AND D( 5)='1' )then
          cVar1S9S7P050N027N052P048(0) <='1';
          else
          cVar1S9S7P050N027N052P048(0) <='0';
          end if;
        if(E( 5)='1' AND B( 6)='0' AND D( 4)='0' AND D( 5)='0' )then
          cVar1S10S7P050N027N052N048(0) <='1';
          else
          cVar1S10S7P050N027N052N048(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S11S7N050P044P023nsss(0) <='1';
          else
          cVar1S11S7N050P044P023nsss(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='1' AND B( 8)='0' AND A(17)='1' )then
          cVar1S12S7N050P044N023P004nsss(0) <='1';
          else
          cVar1S12S7N050P044N023P004nsss(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='1' AND B( 8)='0' AND A(17)='0' )then
          cVar1S13S7N050P044N023N004(0) <='1';
          else
          cVar1S13S7N050P044N023N004(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='1' AND B( 8)='0' AND A(17)='0' )then
          cVar1S14S7N050P044N023N004(0) <='1';
          else
          cVar1S14S7N050P044N023N004(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='1' AND B( 8)='0' AND A(17)='0' )then
          cVar1S15S7N050P044N023N004(0) <='1';
          else
          cVar1S15S7N050P044N023N004(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='1' AND B( 4)='1' )then
          cVar1S16S7N050N044P056P031(0) <='1';
          else
          cVar1S16S7N050N044P056P031(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='1' AND B( 4)='1' )then
          cVar1S17S7N050N044P056P031(0) <='1';
          else
          cVar1S17S7N050N044P056P031(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='1' AND B( 4)='0' )then
          cVar1S18S7N050N044P056N031(0) <='1';
          else
          cVar1S18S7N050N044P056N031(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='1' AND B( 4)='0' )then
          cVar1S19S7N050N044P056N031(0) <='1';
          else
          cVar1S19S7N050N044P056N031(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='1' )then
          cVar1S20S7N050N044N056P038(0) <='1';
          else
          cVar1S20S7N050N044N056P038(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='1' )then
          cVar1S21S7N050N044N056P038(0) <='1';
          else
          cVar1S21S7N050N044N056P038(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S22S7N050N044N056N038(0) <='1';
          else
          cVar1S22S7N050N044N056N038(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S23S7N050N044N056N038(0) <='1';
          else
          cVar1S23S7N050N044N056N038(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S24S7N050N044N056N038(0) <='1';
          else
          cVar1S24S7N050N044N056N038(0) <='0';
          end if;
        if(E( 5)='0' AND D( 6)='0' AND D( 3)='0' AND B(10)='0' )then
          cVar1S25S7N050N044N056N038(0) <='1';
          else
          cVar1S25S7N050N044N056N038(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S0S8P044P023P005nsss(0) <='1';
          else
          cVar1S0S8P044P023P005nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S1S8P044P023N005P004nsss(0) <='1';
          else
          cVar1S1S8P044P023N005P004nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S2S8P044P023N005N004(0) <='1';
          else
          cVar1S2S8P044P023N005N004(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='1' )then
          cVar1S3S8P044N023P004nsss(0) <='1';
          else
          cVar1S3S8P044N023P004nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S4S8P044N023N004P006nsss(0) <='1';
          else
          cVar1S4S8P044N023N004P006nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S5S8P044N023N004N006(0) <='1';
          else
          cVar1S5S8P044N023N004N006(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S6S8P044N023N004N006(0) <='1';
          else
          cVar1S6S8P044N023N004N006(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S7S8P044N023N004N006(0) <='1';
          else
          cVar1S7S8P044N023N004N006(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='1' AND A( 5)='1' )then
          cVar1S8S8N044P050P027P009nsss(0) <='1';
          else
          cVar1S8S8N044P050P027P009nsss(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S9S8N044P050P027N009(0) <='1';
          else
          cVar1S9S8N044P050P027N009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S10S8N044P050P027N009(0) <='1';
          else
          cVar1S10S8N044P050P027N009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S11S8N044P050P027N009(0) <='1';
          else
          cVar1S11S8N044P050P027N009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='0' AND B(16)='1' )then
          cVar1S12S8N044P050N027P026(0) <='1';
          else
          cVar1S12S8N044P050N027P026(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='0' AND B(16)='1' )then
          cVar1S13S8N044P050N027P026(0) <='1';
          else
          cVar1S13S8N044P050N027P026(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='0' AND B(16)='1' )then
          cVar1S14S8N044P050N027P026(0) <='1';
          else
          cVar1S14S8N044P050N027P026(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='0' AND B(16)='0' )then
          cVar1S15S8N044P050N027N026(0) <='1';
          else
          cVar1S15S8N044P050N027N026(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='1' AND B( 6)='0' AND B(16)='0' )then
          cVar1S16S8N044P050N027N026(0) <='1';
          else
          cVar1S16S8N044P050N027N026(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='1' )then
          cVar1S17S8N044N050P014P051(0) <='1';
          else
          cVar1S17S8N044N050P014P051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='1' )then
          cVar1S18S8N044N050P014P051(0) <='1';
          else
          cVar1S18S8N044N050P014P051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='1' )then
          cVar1S19S8N044N050P014P051(0) <='1';
          else
          cVar1S19S8N044N050P014P051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='0' )then
          cVar1S20S8N044N050P014N051(0) <='1';
          else
          cVar1S20S8N044N050P014N051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='0' )then
          cVar1S21S8N044N050P014N051(0) <='1';
          else
          cVar1S21S8N044N050P014N051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='0' AND E(13)='0' )then
          cVar1S22S8N044N050P014N051(0) <='1';
          else
          cVar1S22S8N044N050P014N051(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='1' )then
          cVar1S23S8N044N050P014P032(0) <='1';
          else
          cVar1S23S8N044N050P014P032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='1' )then
          cVar1S24S8N044N050P014P032(0) <='1';
          else
          cVar1S24S8N044N050P014P032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='1' )then
          cVar1S25S8N044N050P014P032(0) <='1';
          else
          cVar1S25S8N044N050P014P032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='0' )then
          cVar1S26S8N044N050P014N032(0) <='1';
          else
          cVar1S26S8N044N050P014N032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='0' )then
          cVar1S27S8N044N050P014N032(0) <='1';
          else
          cVar1S27S8N044N050P014N032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 5)='0' AND A(12)='1' AND B(13)='0' )then
          cVar1S28S8N044N050P014N032(0) <='1';
          else
          cVar1S28S8N044N050P014N032(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='1' AND E(12)='0' )then
          cVar1S0S9P051P028P055nsss(0) <='1';
          else
          cVar1S0S9P051P028P055nsss(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='1' AND E(12)='1' AND D(11)='1' )then
          cVar1S1S9P051P028P055P057nsss(0) <='1';
          else
          cVar1S1S9P051P028P055P057nsss(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='1' )then
          cVar1S2S9P051N028P029nsss(0) <='1';
          else
          cVar1S2S9P051N028P029nsss(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='0' AND B(16)='1' )then
          cVar1S3S9P051N028N029P026(0) <='1';
          else
          cVar1S3S9P051N028N029P026(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='0' AND B(16)='1' )then
          cVar1S4S9P051N028N029P026(0) <='1';
          else
          cVar1S4S9P051N028N029P026(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='0' AND B(16)='1' )then
          cVar1S5S9P051N028N029P026(0) <='1';
          else
          cVar1S5S9P051N028N029P026(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='0' AND B(16)='0' )then
          cVar1S6S9P051N028N029N026(0) <='1';
          else
          cVar1S6S9P051N028N029N026(0) <='0';
          end if;
        if(E(13)='1' AND B(15)='0' AND B( 5)='0' AND B(16)='0' )then
          cVar1S7S9P051N028N029N026(0) <='1';
          else
          cVar1S7S9P051N028N029N026(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='1' AND E(15)='1' AND E( 2)='0' )then
          cVar1S8S9N051P022P043P062nsss(0) <='1';
          else
          cVar1S8S9N051P022P043P062nsss(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar1S9S9N051P022N043P004nsss(0) <='1';
          else
          cVar1S9S9N051P022N043P004nsss(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='1' AND E(15)='0' AND A(17)='0' )then
          cVar1S10S9N051P022N043N004(0) <='1';
          else
          cVar1S10S9N051P022N043N004(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S11S9N051N022P044P023nsss(0) <='1';
          else
          cVar1S11S9N051N022P044P023nsss(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S12S9N051N022P044N023(0) <='1';
          else
          cVar1S12S9N051N022P044N023(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S13S9N051N022P044N023(0) <='1';
          else
          cVar1S13S9N051N022P044N023(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S14S9N051N022P044N023(0) <='1';
          else
          cVar1S14S9N051N022P044N023(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S15S9N051N022N044P050(0) <='1';
          else
          cVar1S15S9N051N022N044P050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S16S9N051N022N044P050(0) <='1';
          else
          cVar1S16S9N051N022N044P050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S17S9N051N022N044P050(0) <='1';
          else
          cVar1S17S9N051N022N044P050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S18S9N051N022N044N050(0) <='1';
          else
          cVar1S18S9N051N022N044N050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S19S9N051N022N044N050(0) <='1';
          else
          cVar1S19S9N051N022N044N050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S20S9N051N022N044N050(0) <='1';
          else
          cVar1S20S9N051N022N044N050(0) <='0';
          end if;
        if(E(13)='0' AND B(18)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S21S9N051N022N044N050(0) <='1';
          else
          cVar1S21S9N051N022N044N050(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='1' AND E(10)='0' )then
          cVar1S0S10P017P037P051P063(0) <='1';
          else
          cVar1S0S10P017P037P051P063(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='1' AND E(10)='0' )then
          cVar1S1S10P017P037P051P063(0) <='1';
          else
          cVar1S1S10P017P037P051P063(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='1' AND E(10)='0' )then
          cVar1S2S10P017P037P051P063(0) <='1';
          else
          cVar1S2S10P017P037P051P063(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='1' )then
          cVar1S3S10P017P037N051P048(0) <='1';
          else
          cVar1S3S10P017P037N051P048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='1' )then
          cVar1S4S10P017P037N051P048(0) <='1';
          else
          cVar1S4S10P017P037N051P048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='1' )then
          cVar1S5S10P017P037N051P048(0) <='1';
          else
          cVar1S5S10P017P037N051P048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='0' )then
          cVar1S6S10P017P037N051N048(0) <='1';
          else
          cVar1S6S10P017P037N051N048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='0' )then
          cVar1S7S10P017P037N051N048(0) <='1';
          else
          cVar1S7S10P017P037N051N048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='0' AND E(13)='0' AND D( 5)='0' )then
          cVar1S8S10P017P037N051N048(0) <='1';
          else
          cVar1S8S10P017P037N051N048(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='1' AND D( 1)='0' )then
          cVar1S9S10P017P037P019P064(0) <='1';
          else
          cVar1S9S10P017P037P019P064(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='1' AND D( 1)='0' )then
          cVar1S10S10P017P037P019P064(0) <='1';
          else
          cVar1S10S10P017P037P019P064(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='1' AND D( 1)='0' )then
          cVar1S11S10P017P037P019P064(0) <='1';
          else
          cVar1S11S10P017P037P019P064(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='1' AND D( 1)='1' )then
          cVar1S12S10P017P037P019P064(0) <='1';
          else
          cVar1S12S10P017P037P019P064(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='1' AND D( 1)='1' )then
          cVar1S13S10P017P037P019P064(0) <='1';
          else
          cVar1S13S10P017P037P019P064(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='0' AND E(10)='0' )then
          cVar1S14S10P017P037N019P063(0) <='1';
          else
          cVar1S14S10P017P037N019P063(0) <='0';
          end if;
        if(A( 1)='0' AND B( 1)='1' AND A( 0)='0' AND E(10)='1' )then
          cVar1S15S10P017P037N019P063(0) <='1';
          else
          cVar1S15S10P017P037N019P063(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND D( 0)='0' )then
          cVar1S16S10P017P064P019P068(0) <='1';
          else
          cVar1S16S10P017P064P019P068(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND D( 0)='0' )then
          cVar1S17S10P017P064P019P068(0) <='1';
          else
          cVar1S17S10P017P064P019P068(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S18S10P017P064P019P068(0) <='1';
          else
          cVar1S18S10P017P064P019P068(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND A( 2)='1' )then
          cVar1S19S10P017P064P019P015(0) <='1';
          else
          cVar1S19S10P017P064P019P015(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND A( 2)='1' )then
          cVar1S20S10P017P064P019P015(0) <='1';
          else
          cVar1S20S10P017P064P019P015(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND A( 2)='1' )then
          cVar1S21S10P017P064P019P015(0) <='1';
          else
          cVar1S21S10P017P064P019P015(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND A( 2)='0' )then
          cVar1S22S10P017P064P019N015(0) <='1';
          else
          cVar1S22S10P017P064P019N015(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='1' AND D( 9)='0' )then
          cVar1S23S10P017N064P015P065(0) <='1';
          else
          cVar1S23S10P017N064P015P065(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='1' AND D( 9)='0' )then
          cVar1S24S10P017N064P015P065(0) <='1';
          else
          cVar1S24S10P017N064P015P065(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='1' AND D( 9)='0' )then
          cVar1S25S10P017N064P015P065(0) <='1';
          else
          cVar1S25S10P017N064P015P065(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='1' AND D( 9)='1' )then
          cVar1S26S10P017N064P015P065(0) <='1';
          else
          cVar1S26S10P017N064P015P065(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='1' )then
          cVar1S27S10P017N064N015P037(0) <='1';
          else
          cVar1S27S10P017N064N015P037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='1' )then
          cVar1S28S10P017N064N015P037(0) <='1';
          else
          cVar1S28S10P017N064N015P037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='1' )then
          cVar1S29S10P017N064N015P037(0) <='1';
          else
          cVar1S29S10P017N064N015P037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='1' )then
          cVar1S30S10P017N064N015P037(0) <='1';
          else
          cVar1S30S10P017N064N015P037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='0' )then
          cVar1S31S10P017N064N015N037(0) <='1';
          else
          cVar1S31S10P017N064N015N037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='0' )then
          cVar1S32S10P017N064N015N037(0) <='1';
          else
          cVar1S32S10P017N064N015N037(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND A( 2)='0' AND B( 1)='0' )then
          cVar1S33S10P017N064N015N037(0) <='1';
          else
          cVar1S33S10P017N064N015N037(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S11P048P025P007nsss(0) <='1';
          else
          cVar1S0S11P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='1' )then
          cVar1S1S11P048P025N007P006nsss(0) <='1';
          else
          cVar1S1S11P048P025N007P006nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S2S11P048P025N007N006(0) <='1';
          else
          cVar1S2S11P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S3S11P048P025N007N006(0) <='1';
          else
          cVar1S3S11P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S4S11P048P025N007N006(0) <='1';
          else
          cVar1S4S11P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='0' )then
          cVar1S5S11P048N025P027P011(0) <='1';
          else
          cVar1S5S11P048N025P027P011(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='0' )then
          cVar1S6S11P048N025P027P011(0) <='1';
          else
          cVar1S6S11P048N025P027P011(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='0' )then
          cVar1S7S11P048N025P027P011(0) <='1';
          else
          cVar1S7S11P048N025P027P011(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='1' )then
          cVar1S8S11P048N025P027P011(0) <='1';
          else
          cVar1S8S11P048N025P027P011(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S9S11P048N025N027P007(0) <='1';
          else
          cVar1S9S11P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S10S11P048N025N027P007(0) <='1';
          else
          cVar1S10S11P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S11S11P048N025N027P007(0) <='1';
          else
          cVar1S11S11P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S12S11P048N025N027P007(0) <='1';
          else
          cVar1S12S11P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND B(15)='1' AND E(12)='0' )then
          cVar1S13S11N048P051P028P055nsss(0) <='1';
          else
          cVar1S13S11N048P051P028P055nsss(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND B(15)='0' AND B( 5)='1' )then
          cVar1S14S11N048P051N028P029nsss(0) <='1';
          else
          cVar1S14S11N048P051N028P029nsss(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND B(15)='0' AND B( 5)='0' )then
          cVar1S15S11N048P051N028N029(0) <='1';
          else
          cVar1S15S11N048P051N028N029(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND B(15)='0' AND B( 5)='0' )then
          cVar1S16S11N048P051N028N029(0) <='1';
          else
          cVar1S16S11N048P051N028N029(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND B(15)='0' AND B( 5)='0' )then
          cVar1S17S11N048P051N028N029(0) <='1';
          else
          cVar1S17S11N048P051N028N029(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='1' AND E(15)='1' )then
          cVar1S18S11N048N051P022P043(0) <='1';
          else
          cVar1S18S11N048N051P022P043(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S19S11N048N051P022N043(0) <='1';
          else
          cVar1S19S11N048N051P022N043(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S20S11N048N051P022N043(0) <='1';
          else
          cVar1S20S11N048N051P022N043(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S21S11N048N051P022N043(0) <='1';
          else
          cVar1S21S11N048N051P022N043(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='1' )then
          cVar1S22S11N048N051N022P023(0) <='1';
          else
          cVar1S22S11N048N051N022P023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='1' )then
          cVar1S23S11N048N051N022P023(0) <='1';
          else
          cVar1S23S11N048N051N022P023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='1' )then
          cVar1S24S11N048N051N022P023(0) <='1';
          else
          cVar1S24S11N048N051N022P023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='0' )then
          cVar1S25S11N048N051N022N023(0) <='1';
          else
          cVar1S25S11N048N051N022N023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='0' )then
          cVar1S26S11N048N051N022N023(0) <='1';
          else
          cVar1S26S11N048N051N022N023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='0' )then
          cVar1S27S11N048N051N022N023(0) <='1';
          else
          cVar1S27S11N048N051N022N023(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(18)='0' AND B( 8)='0' )then
          cVar1S28S11N048N051N022N023(0) <='1';
          else
          cVar1S28S11N048N051N022N023(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S12P048P025P007nsss(0) <='1';
          else
          cVar1S0S12P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='1' )then
          cVar1S1S12P048P025N007P006nsss(0) <='1';
          else
          cVar1S1S12P048P025N007P006nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S2S12P048P025N007N006(0) <='1';
          else
          cVar1S2S12P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S3S12P048P025N007N006(0) <='1';
          else
          cVar1S3S12P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(16)='0' )then
          cVar1S4S12P048P025N007N006(0) <='1';
          else
          cVar1S4S12P048P025N007N006(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND D( 4)='0' )then
          cVar1S5S12P048N025P027P052nsss(0) <='1';
          else
          cVar1S5S12P048N025P027P052nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 9)='0' )then
          cVar1S6S12P048N025N027P067(0) <='1';
          else
          cVar1S6S12P048N025N027P067(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 9)='0' )then
          cVar1S7S12P048N025N027P067(0) <='1';
          else
          cVar1S7S12P048N025N027P067(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 9)='0' )then
          cVar1S8S12P048N025N027P067(0) <='1';
          else
          cVar1S8S12P048N025N027P067(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='1' AND A( 3)='0' )then
          cVar1S9S12N048P001P051P013(0) <='1';
          else
          cVar1S9S12N048P001P051P013(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='1' AND A( 3)='0' )then
          cVar1S10S12N048P001P051P013(0) <='1';
          else
          cVar1S10S12N048P001P051P013(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='1' AND A( 3)='0' )then
          cVar1S11S12N048P001P051P013(0) <='1';
          else
          cVar1S11S12N048P001P051P013(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='1' AND A( 3)='1' )then
          cVar1S12S12N048P001P051P013(0) <='1';
          else
          cVar1S12S12N048P001P051P013(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='1' AND A( 3)='1' )then
          cVar1S13S12N048P001P051P013(0) <='1';
          else
          cVar1S13S12N048P001P051P013(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='0' AND A(15)='0' )then
          cVar1S14S12N048P001N051P008(0) <='1';
          else
          cVar1S14S12N048P001N051P008(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='0' AND A(15)='0' )then
          cVar1S15S12N048P001N051P008(0) <='1';
          else
          cVar1S15S12N048P001N051P008(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='0' AND A(15)='1' )then
          cVar1S16S12N048P001N051P008(0) <='1';
          else
          cVar1S16S12N048P001N051P008(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='0' AND A(15)='1' )then
          cVar1S17S12N048P001N051P008(0) <='1';
          else
          cVar1S17S12N048P001N051P008(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='0' AND E(13)='0' AND A(15)='1' )then
          cVar1S18S12N048P001N051P008(0) <='1';
          else
          cVar1S18S12N048P001N051P008(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='1' AND D(15)='1' )then
          cVar1S19S12N048P001P041nsss(0) <='1';
          else
          cVar1S19S12N048P001P041nsss(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='1' AND D(15)='0' AND A( 1)='1' )then
          cVar1S20S12N048P001N041P017(0) <='1';
          else
          cVar1S20S12N048P001N041P017(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='1' AND D(15)='0' AND A( 1)='1' )then
          cVar1S21S12N048P001N041P017(0) <='1';
          else
          cVar1S21S12N048P001N041P017(0) <='0';
          end if;
        if(D( 5)='0' AND A( 9)='1' AND D(15)='0' AND A( 1)='0' )then
          cVar1S22S12N048P001N041N017(0) <='1';
          else
          cVar1S22S12N048P001N041N017(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S13P048P025P007nsss(0) <='1';
          else
          cVar1S0S13P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(11)='0' )then
          cVar1S1S13P048P025N007P016nsss(0) <='1';
          else
          cVar1S1S13P048P025N007P016nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='0' )then
          cVar1S2S13P048N025P027P011nsss(0) <='1';
          else
          cVar1S2S13P048N025P027P011nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 4)='1' )then
          cVar1S3S13P048N025P027P011(0) <='1';
          else
          cVar1S3S13P048N025P027P011(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S4S13P048N025N027P007(0) <='1';
          else
          cVar1S4S13P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S5S13P048N025N027P007(0) <='1';
          else
          cVar1S5S13P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S6S13P048N025N027P007(0) <='1';
          else
          cVar1S6S13P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar1S7S13P048N025N027P007(0) <='1';
          else
          cVar1S7S13P048N025N027P007(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar1S8S13N048P051P008P013(0) <='1';
          else
          cVar1S8S13N048P051P008P013(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar1S9S13N048P051P008P013(0) <='1';
          else
          cVar1S9S13N048P051P008P013(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='1' )then
          cVar1S10S13N048P051N008P028(0) <='1';
          else
          cVar1S10S13N048P051N008P028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='1' )then
          cVar1S11S13N048P051N008P028(0) <='1';
          else
          cVar1S11S13N048P051N008P028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='1' )then
          cVar1S12S13N048P051N008P028(0) <='1';
          else
          cVar1S12S13N048P051N008P028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='1' )then
          cVar1S13S13N048P051N008P028(0) <='1';
          else
          cVar1S13S13N048P051N008P028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='0' )then
          cVar1S14S13N048P051N008N028(0) <='1';
          else
          cVar1S14S13N048P051N008N028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='0' )then
          cVar1S15S13N048P051N008N028(0) <='1';
          else
          cVar1S15S13N048P051N008N028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='1' AND A(15)='0' AND B(15)='0' )then
          cVar1S16S13N048P051N008N028(0) <='1';
          else
          cVar1S16S13N048P051N008N028(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='1' AND B( 9)='1' )then
          cVar1S17S13N048N051P038P021nsss(0) <='1';
          else
          cVar1S17S13N048N051P038P021nsss(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='1' AND B( 9)='0' )then
          cVar1S18S13N048N051P038N021(0) <='1';
          else
          cVar1S18S13N048N051P038N021(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='1' AND B( 9)='0' )then
          cVar1S19S13N048N051P038N021(0) <='1';
          else
          cVar1S19S13N048N051P038N021(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='1' AND B( 9)='0' )then
          cVar1S20S13N048N051P038N021(0) <='1';
          else
          cVar1S20S13N048N051P038N021(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='1' )then
          cVar1S21S13N048N051N038P061(0) <='1';
          else
          cVar1S21S13N048N051N038P061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='1' )then
          cVar1S22S13N048N051N038P061(0) <='1';
          else
          cVar1S22S13N048N051N038P061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='1' )then
          cVar1S23S13N048N051N038P061(0) <='1';
          else
          cVar1S23S13N048N051N038P061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='0' )then
          cVar1S24S13N048N051N038N061(0) <='1';
          else
          cVar1S24S13N048N051N038N061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='0' )then
          cVar1S25S13N048N051N038N061(0) <='1';
          else
          cVar1S25S13N048N051N038N061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='0' )then
          cVar1S26S13N048N051N038N061(0) <='1';
          else
          cVar1S26S13N048N051N038N061(0) <='0';
          end if;
        if(D( 5)='0' AND E(13)='0' AND B(10)='0' AND D(10)='0' )then
          cVar1S27S13N048N051N038N061(0) <='1';
          else
          cVar1S27S13N048N051N038N061(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S0S14P017P048P025nsss(0) <='1';
          else
          cVar1S0S14P017P048P025nsss(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S1S14P017P048N025P027(0) <='1';
          else
          cVar1S1S14P017P048N025P027(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S2S14P017P048N025P027(0) <='1';
          else
          cVar1S2S14P017P048N025P027(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S3S14P017P048N025P027(0) <='1';
          else
          cVar1S3S14P017P048N025P027(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S4S14P017P048N025N027(0) <='1';
          else
          cVar1S4S14P017P048N025N027(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S5S14P017P048N025N027(0) <='1';
          else
          cVar1S5S14P017P048N025N027(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S6S14P017N048P044P023nsss(0) <='1';
          else
          cVar1S6S14P017N048P044P023nsss(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S7S14P017N048P044N023(0) <='1';
          else
          cVar1S7S14P017N048P044N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S8S14P017N048P044N023(0) <='1';
          else
          cVar1S8S14P017N048P044N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S9S14P017N048P044N023(0) <='1';
          else
          cVar1S9S14P017N048P044N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S10S14P017N048P044N023(0) <='1';
          else
          cVar1S10S14P017N048P044N023(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='0' AND B(10)='1' )then
          cVar1S11S14P017N048N044P038(0) <='1';
          else
          cVar1S11S14P017N048N044P038(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='0' AND B(10)='1' )then
          cVar1S12S14P017N048N044P038(0) <='1';
          else
          cVar1S12S14P017N048N044P038(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='0' AND B(10)='1' )then
          cVar1S13S14P017N048N044P038(0) <='1';
          else
          cVar1S13S14P017N048N044P038(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='0' AND B(10)='0' )then
          cVar1S14S14P017N048N044N038(0) <='1';
          else
          cVar1S14S14P017N048N044N038(0) <='0';
          end if;
        if(A( 1)='0' AND D( 5)='0' AND D( 6)='0' AND B(10)='0' )then
          cVar1S15S14P017N048N044N038(0) <='1';
          else
          cVar1S15S14P017N048N044N038(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND A( 5)='0' )then
          cVar1S16S14P017P064P019P009(0) <='1';
          else
          cVar1S16S14P017P064P019P009(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND A( 5)='0' )then
          cVar1S17S14P017P064P019P009(0) <='1';
          else
          cVar1S17S14P017P064P019P009(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='0' AND A( 5)='0' )then
          cVar1S18S14P017P064P019P009(0) <='1';
          else
          cVar1S18S14P017P064P019P009(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND E( 5)='1' )then
          cVar1S19S14P017P064P019P050nsss(0) <='1';
          else
          cVar1S19S14P017P064P019P050nsss(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND E( 5)='0' )then
          cVar1S20S14P017P064P019N050(0) <='1';
          else
          cVar1S20S14P017P064P019N050(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND A( 0)='1' AND E( 5)='0' )then
          cVar1S21S14P017P064P019N050(0) <='1';
          else
          cVar1S21S14P017P064P019N050(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='1' AND A( 8)='0' )then
          cVar1S22S14P017N064P061P003(0) <='1';
          else
          cVar1S22S14P017N064P061P003(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='1' AND A( 8)='0' )then
          cVar1S23S14P017N064P061P003(0) <='1';
          else
          cVar1S23S14P017N064P061P003(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='1' AND A( 8)='0' )then
          cVar1S24S14P017N064P061P003(0) <='1';
          else
          cVar1S24S14P017N064P061P003(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='1' AND A( 8)='0' )then
          cVar1S25S14P017N064P061P003(0) <='1';
          else
          cVar1S25S14P017N064P061P003(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S26S14P017N064N061P051(0) <='1';
          else
          cVar1S26S14P017N064N061P051(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S27S14P017N064N061P051(0) <='1';
          else
          cVar1S27S14P017N064N061P051(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='0' AND E(13)='1' )then
          cVar1S28S14P017N064N061P051(0) <='1';
          else
          cVar1S28S14P017N064N061P051(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='0' AND E(13)='0' )then
          cVar1S29S14P017N064N061N051(0) <='1';
          else
          cVar1S29S14P017N064N061N051(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND D(10)='0' AND E(13)='0' )then
          cVar1S30S14P017N064N061N051(0) <='1';
          else
          cVar1S30S14P017N064N061N051(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S0S15P044P023P005nsss(0) <='1';
          else
          cVar1S0S15P044P023P005nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S1S15P044P023N005P004nsss(0) <='1';
          else
          cVar1S1S15P044P023N005P004nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S2S15P044P023N005N004(0) <='1';
          else
          cVar1S2S15P044P023N005N004(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S3S15P044P023N005N004(0) <='1';
          else
          cVar1S3S15P044P023N005N004(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='1' AND A( 2)='0' )then
          cVar1S4S15P044N023P022P015nsss(0) <='1';
          else
          cVar1S4S15P044N023P022P015nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='1' )then
          cVar1S5S15P044N023N022P025(0) <='1';
          else
          cVar1S5S15P044N023N022P025(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='1' )then
          cVar1S6S15P044N023N022P025(0) <='1';
          else
          cVar1S6S15P044N023N022P025(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='1' )then
          cVar1S7S15P044N023N022P025(0) <='1';
          else
          cVar1S7S15P044N023N022P025(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='0' )then
          cVar1S8S15P044N023N022N025(0) <='1';
          else
          cVar1S8S15P044N023N022N025(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND B(18)='0' AND B( 7)='0' )then
          cVar1S9S15P044N023N022N025(0) <='1';
          else
          cVar1S9S15P044N023N022N025(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S10S15N044P048P025P007nsss(0) <='1';
          else
          cVar1S10S15N044P048P025P007nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S11S15N044P048P025N007(0) <='1';
          else
          cVar1S11S15N044P048P025N007(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S12S15N044P048P025N007(0) <='1';
          else
          cVar1S12S15N044P048P025N007(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S13S15N044P048P025N007(0) <='1';
          else
          cVar1S13S15N044P048P025N007(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S14S15N044P048N025P027(0) <='1';
          else
          cVar1S14S15N044P048N025P027(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S15S15N044P048N025P027(0) <='1';
          else
          cVar1S15S15N044P048N025P027(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S16S15N044P048N025N027(0) <='1';
          else
          cVar1S16S15N044P048N025N027(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S17S15N044P048N025N027(0) <='1';
          else
          cVar1S17S15N044P048N025N027(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S18S15N044P048N025N027(0) <='1';
          else
          cVar1S18S15N044P048N025N027(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='1' )then
          cVar1S19S15N044N048P007P040(0) <='1';
          else
          cVar1S19S15N044N048P007P040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='1' )then
          cVar1S20S15N044N048P007P040(0) <='1';
          else
          cVar1S20S15N044N048P007P040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='1' )then
          cVar1S21S15N044N048P007P040(0) <='1';
          else
          cVar1S21S15N044N048P007P040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='0' )then
          cVar1S22S15N044N048P007N040(0) <='1';
          else
          cVar1S22S15N044N048P007N040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='0' )then
          cVar1S23S15N044N048P007N040(0) <='1';
          else
          cVar1S23S15N044N048P007N040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='0' AND D( 7)='0' )then
          cVar1S24S15N044N048P007N040(0) <='1';
          else
          cVar1S24S15N044N048P007N040(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='1' AND E(15)='1' )then
          cVar1S25S15N044N048P007P043(0) <='1';
          else
          cVar1S25S15N044N048P007P043(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='1' AND E(15)='1' )then
          cVar1S26S15N044N048P007P043(0) <='1';
          else
          cVar1S26S15N044N048P007P043(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='1' AND E(15)='1' )then
          cVar1S27S15N044N048P007P043(0) <='1';
          else
          cVar1S27S15N044N048P007P043(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='1' AND E(15)='0' )then
          cVar1S28S15N044N048P007N043(0) <='1';
          else
          cVar1S28S15N044N048P007N043(0) <='0';
          end if;
        if(D( 6)='0' AND D( 5)='0' AND A( 6)='1' AND E(15)='0' )then
          cVar1S29S15N044N048P007N043(0) <='1';
          else
          cVar1S29S15N044N048P007N043(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='1' AND B( 7)='1' AND E( 5)='0' )then
          cVar1S0S16P067P048P025P050nsss(0) <='1';
          else
          cVar1S0S16P067P048P025P050nsss(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S1S16P067P048N025P027nsss(0) <='1';
          else
          cVar1S1S16P067P048N025P027nsss(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S2S16P067P048N025N027(0) <='1';
          else
          cVar1S2S16P067P048N025N027(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S3S16P067P048N025N027(0) <='1';
          else
          cVar1S3S16P067P048N025N027(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S4S16P067P048N025N027(0) <='1';
          else
          cVar1S4S16P067P048N025N027(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S5S16P067N048P051P008(0) <='1';
          else
          cVar1S5S16P067N048P051P008(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S6S16P067N048P051P008(0) <='1';
          else
          cVar1S6S16P067N048P051P008(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S7S16P067N048P051P008(0) <='1';
          else
          cVar1S7S16P067N048P051P008(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S8S16P067N048P051N008(0) <='1';
          else
          cVar1S8S16P067N048P051N008(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S9S16P067N048P051N008(0) <='1';
          else
          cVar1S9S16P067N048P051N008(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='1' )then
          cVar1S10S16P067N048N051P022(0) <='1';
          else
          cVar1S10S16P067N048N051P022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='1' )then
          cVar1S11S16P067N048N051P022(0) <='1';
          else
          cVar1S11S16P067N048N051P022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='1' )then
          cVar1S12S16P067N048N051P022(0) <='1';
          else
          cVar1S12S16P067N048N051P022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='0' )then
          cVar1S13S16P067N048N051N022(0) <='1';
          else
          cVar1S13S16P067N048N051N022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='0' )then
          cVar1S14S16P067N048N051N022(0) <='1';
          else
          cVar1S14S16P067N048N051N022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='0' )then
          cVar1S15S16P067N048N051N022(0) <='1';
          else
          cVar1S15S16P067N048N051N022(0) <='0';
          end if;
        if(E( 9)='0' AND D( 5)='0' AND E(13)='0' AND B(18)='0' )then
          cVar1S16S16P067N048N051N022(0) <='1';
          else
          cVar1S16S16P067N048N051N022(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(14)='0' )then
          cVar1S17S16P067P069P018P010(0) <='1';
          else
          cVar1S17S16P067P069P018P010(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(14)='0' )then
          cVar1S18S16P067P069P018P010(0) <='1';
          else
          cVar1S18S16P067P069P018P010(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(14)='0' )then
          cVar1S19S16P067P069P018P010(0) <='1';
          else
          cVar1S19S16P067P069P018P010(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(14)='1' )then
          cVar1S20S16P067P069P018P010(0) <='1';
          else
          cVar1S20S16P067P069P018P010(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar1S21S16P067P069N018P019(0) <='1';
          else
          cVar1S21S16P067P069N018P019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar1S22S16P067P069N018P019(0) <='1';
          else
          cVar1S22S16P067P069N018P019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar1S23S16P067P069N018P019(0) <='1';
          else
          cVar1S23S16P067P069N018P019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S24S16P067P069N018N019(0) <='1';
          else
          cVar1S24S16P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S25S16P067P069N018N019(0) <='1';
          else
          cVar1S25S16P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S26S16P067P069N018N019(0) <='1';
          else
          cVar1S26S16P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 4)='1' )then
          cVar1S27S16P067N069P052nsss(0) <='1';
          else
          cVar1S27S16P067N069P052nsss(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 4)='0' AND D( 9)='1' )then
          cVar1S28S16P067N069N052P065(0) <='1';
          else
          cVar1S28S16P067N069N052P065(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 4)='0' AND D( 9)='1' )then
          cVar1S29S16P067N069N052P065(0) <='1';
          else
          cVar1S29S16P067N069N052P065(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 4)='0' AND D( 9)='0' )then
          cVar1S30S16P067N069N052N065(0) <='1';
          else
          cVar1S30S16P067N069N052N065(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND E( 2)='0' )then
          cVar1S0S17P022P043P062nsss(0) <='1';
          else
          cVar1S0S17P022P043P062nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND D( 8)='0' AND A(17)='1' )then
          cVar1S1S17P022N043P069P004nsss(0) <='1';
          else
          cVar1S1S17P022N043P069P004nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND D( 8)='0' AND A(17)='0' )then
          cVar1S2S17P022N043P069N004(0) <='1';
          else
          cVar1S2S17P022N043P069N004(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND D( 8)='0' AND A(17)='0' )then
          cVar1S3S17P022N043P069N004(0) <='1';
          else
          cVar1S3S17P022N043P069N004(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S4S17N022P048P025P007nsss(0) <='1';
          else
          cVar1S4S17N022P048P025P007nsss(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S5S17N022P048P025N007(0) <='1';
          else
          cVar1S5S17N022P048P025N007(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S6S17N022P048P025N007(0) <='1';
          else
          cVar1S6S17N022P048P025N007(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S7S17N022P048P025N007(0) <='1';
          else
          cVar1S7S17N022P048P025N007(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S8S17N022P048N025P027(0) <='1';
          else
          cVar1S8S17N022P048N025P027(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S9S17N022P048N025N027(0) <='1';
          else
          cVar1S9S17N022P048N025N027(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S10S17N022P048N025N027(0) <='1';
          else
          cVar1S10S17N022P048N025N027(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S11S17N022P048N025N027(0) <='1';
          else
          cVar1S11S17N022P048N025N027(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S12S17N022N048P051P008(0) <='1';
          else
          cVar1S12S17N022N048P051P008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S13S17N022N048P051P008(0) <='1';
          else
          cVar1S13S17N022N048P051P008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S14S17N022N048P051P008(0) <='1';
          else
          cVar1S14S17N022N048P051P008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S15S17N022N048P051N008(0) <='1';
          else
          cVar1S15S17N022N048P051N008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S16S17N022N048P051N008(0) <='1';
          else
          cVar1S16S17N022N048P051N008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S17S17N022N048P051N008(0) <='1';
          else
          cVar1S17S17N022N048P051N008(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='1' )then
          cVar1S18S17N022N048N051P038(0) <='1';
          else
          cVar1S18S17N022N048N051P038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='1' )then
          cVar1S19S17N022N048N051P038(0) <='1';
          else
          cVar1S19S17N022N048N051P038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='1' )then
          cVar1S20S17N022N048N051P038(0) <='1';
          else
          cVar1S20S17N022N048N051P038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='0' )then
          cVar1S21S17N022N048N051N038(0) <='1';
          else
          cVar1S21S17N022N048N051N038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='0' )then
          cVar1S22S17N022N048N051N038(0) <='1';
          else
          cVar1S22S17N022N048N051N038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='0' )then
          cVar1S23S17N022N048N051N038(0) <='1';
          else
          cVar1S23S17N022N048N051N038(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND E(13)='0' AND B(10)='0' )then
          cVar1S24S17N022N048N051N038(0) <='1';
          else
          cVar1S24S17N022N048N051N038(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' )then
          cVar1S0S18P041P020nsss(0) <='1';
          else
          cVar1S0S18P041P020nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='1' AND B( 0)='1' )then
          cVar1S1S18P041N020P021P039nsss(0) <='1';
          else
          cVar1S1S18P041N020P021P039nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='1' )then
          cVar1S2S18P041N020N021P022(0) <='1';
          else
          cVar1S2S18P041N020N021P022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='1' )then
          cVar1S3S18P041N020N021P022(0) <='1';
          else
          cVar1S3S18P041N020N021P022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='0' )then
          cVar1S4S18P041N020N021N022(0) <='1';
          else
          cVar1S4S18P041N020N021N022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='0' )then
          cVar1S5S18P041N020N021N022(0) <='1';
          else
          cVar1S5S18P041N020N021N022(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S6S18N041P039P020P044(0) <='1';
          else
          cVar1S6S18N041P039P020P044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S7S18N041P039P020P044(0) <='1';
          else
          cVar1S7S18N041P039P020P044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S8S18N041P039P020P044(0) <='1';
          else
          cVar1S8S18N041P039P020P044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S9S18N041P039P020N044(0) <='1';
          else
          cVar1S9S18N041P039P020N044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S10S18N041P039P020N044(0) <='1';
          else
          cVar1S10S18N041P039P020N044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S11S18N041P039P020N044(0) <='1';
          else
          cVar1S11S18N041P039P020N044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S12S18N041P039P020N044(0) <='1';
          else
          cVar1S12S18N041P039P020N044(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='1' AND D( 7)='1' )then
          cVar1S13S18N041P039P020P040(0) <='1';
          else
          cVar1S13S18N041P039P020P040(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='1' AND D( 7)='0' )then
          cVar1S14S18N041P039P020N040(0) <='1';
          else
          cVar1S14S18N041P039P020N040(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND B(19)='1' AND D( 7)='0' )then
          cVar1S15S18N041P039P020N040(0) <='1';
          else
          cVar1S15S18N041P039P020N040(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND A( 7)='1' )then
          cVar1S16S18N041P039P005nsss(0) <='1';
          else
          cVar1S16S18N041P039P005nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND A( 7)='0' AND B(19)='1' )then
          cVar1S17S18N041P039N005P020nsss(0) <='1';
          else
          cVar1S17S18N041P039N005P020nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND A( 7)='0' AND B(19)='0' )then
          cVar1S18S18N041P039N005N020(0) <='1';
          else
          cVar1S18S18N041P039N005N020(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' )then
          cVar1S0S19P041P020nsss(0) <='1';
          else
          cVar1S0S19P041P020nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='1' AND A( 8)='1' )then
          cVar1S1S19P041N020P021P003nsss(0) <='1';
          else
          cVar1S1S19P041N020P021P003nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='1' AND A( 8)='0' )then
          cVar1S2S19P041N020P021N003(0) <='1';
          else
          cVar1S2S19P041N020P021N003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='1' )then
          cVar1S3S19P041N020N021P022(0) <='1';
          else
          cVar1S3S19P041N020N021P022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='1' )then
          cVar1S4S19P041N020N021P022(0) <='1';
          else
          cVar1S4S19P041N020N021P022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='0' )then
          cVar1S5S19P041N020N021N022(0) <='1';
          else
          cVar1S5S19P041N020N021N022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='0' )then
          cVar1S6S19P041N020N021N022(0) <='1';
          else
          cVar1S6S19P041N020N021N022(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND B(18)='0' )then
          cVar1S7S19P041N020N021N022(0) <='1';
          else
          cVar1S7S19P041N020N021N022(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S8S19N041P039P044P023(0) <='1';
          else
          cVar1S8S19N041P039P044P023(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S9S19N041P039P044P023(0) <='1';
          else
          cVar1S9S19N041P039P044P023(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S10S19N041P039P044P023(0) <='1';
          else
          cVar1S10S19N041P039P044P023(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S11S19N041P039P044N023psss(0) <='1';
          else
          cVar1S11S19N041P039P044N023psss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S12S19N041P039N044P050(0) <='1';
          else
          cVar1S12S19N041P039N044P050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S13S19N041P039N044P050(0) <='1';
          else
          cVar1S13S19N041P039N044P050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S14S19N041P039N044P050(0) <='1';
          else
          cVar1S14S19N041P039N044P050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='1' )then
          cVar1S15S19N041P039N044P050(0) <='1';
          else
          cVar1S15S19N041P039N044P050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S16S19N041P039N044N050(0) <='1';
          else
          cVar1S16S19N041P039N044N050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S17S19N041P039N044N050(0) <='1';
          else
          cVar1S17S19N041P039N044N050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND D( 6)='0' AND E( 5)='0' )then
          cVar1S18S19N041P039N044N050(0) <='1';
          else
          cVar1S18S19N041P039N044N050(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND A( 7)='1' )then
          cVar1S19S19N041P039P005nsss(0) <='1';
          else
          cVar1S19S19N041P039P005nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND A( 7)='0' AND D( 1)='0' )then
          cVar1S20S19N041P039N005N064(0) <='1';
          else
          cVar1S20S19N041P039N005N064(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S0S20P011P029P048P025(0) <='1';
          else
          cVar1S0S20P011P029P048P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S1S20P011P029P048P025(0) <='1';
          else
          cVar1S1S20P011P029P048P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S2S20P011P029P048P025(0) <='1';
          else
          cVar1S2S20P011P029P048P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='1' AND B( 7)='0' )then
          cVar1S3S20P011P029P048N025psss(0) <='1';
          else
          cVar1S3S20P011P029P048N025psss(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='1' )then
          cVar1S4S20P011P029N048P041(0) <='1';
          else
          cVar1S4S20P011P029N048P041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='1' )then
          cVar1S5S20P011P029N048P041(0) <='1';
          else
          cVar1S5S20P011P029N048P041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='1' )then
          cVar1S6S20P011P029N048P041(0) <='1';
          else
          cVar1S6S20P011P029N048P041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='0' )then
          cVar1S7S20P011P029N048N041(0) <='1';
          else
          cVar1S7S20P011P029N048N041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='0' )then
          cVar1S8S20P011P029N048N041(0) <='1';
          else
          cVar1S8S20P011P029N048N041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='0' )then
          cVar1S9S20P011P029N048N041(0) <='1';
          else
          cVar1S9S20P011P029N048N041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND D( 5)='0' AND D(15)='0' )then
          cVar1S10S20P011P029N048N041(0) <='1';
          else
          cVar1S10S20P011P029N048N041(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A(14)='1' AND D( 4)='1' )then
          cVar1S11S20P011P029P010P052nsss(0) <='1';
          else
          cVar1S11S20P011P029P010P052nsss(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A(14)='1' AND D( 4)='0' )then
          cVar1S12S20P011P029P010N052(0) <='1';
          else
          cVar1S12S20P011P029P010N052(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A(14)='0' AND A( 5)='1' )then
          cVar1S13S20P011P029N010P009(0) <='1';
          else
          cVar1S13S20P011P029N010P009(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A(14)='0' AND A( 5)='1' )then
          cVar1S14S20P011P029N010P009(0) <='1';
          else
          cVar1S14S20P011P029N010P009(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A(14)='0' AND A( 5)='0' )then
          cVar1S15S20P011P029N010N009(0) <='1';
          else
          cVar1S15S20P011P029N010N009(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND D( 2)='0' AND A(12)='0' )then
          cVar1S16S20P011P029P060P014(0) <='1';
          else
          cVar1S16S20P011P029P060P014(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND D( 2)='0' AND A(12)='0' )then
          cVar1S17S20P011P029P060P014(0) <='1';
          else
          cVar1S17S20P011P029P060P014(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND D( 2)='0' AND A(12)='1' )then
          cVar1S18S20P011P029P060P014(0) <='1';
          else
          cVar1S18S20P011P029P060P014(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND D( 2)='0' AND A(12)='1' )then
          cVar1S19S20P011P029P060P014(0) <='1';
          else
          cVar1S19S20P011P029P060P014(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='1' AND B( 3)='0' )then
          cVar1S20S20P011N029P015P033(0) <='1';
          else
          cVar1S20S20P011N029P015P033(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='1' AND B( 3)='0' )then
          cVar1S21S20P011N029P015P033(0) <='1';
          else
          cVar1S21S20P011N029P015P033(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='1' AND B( 3)='0' )then
          cVar1S22S20P011N029P015P033(0) <='1';
          else
          cVar1S22S20P011N029P015P033(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='1' AND B( 3)='1' )then
          cVar1S23S20P011N029P015P033(0) <='1';
          else
          cVar1S23S20P011N029P015P033(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S24S20P011N029N015P017(0) <='1';
          else
          cVar1S24S20P011N029N015P017(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S25S20P011N029N015P017(0) <='1';
          else
          cVar1S25S20P011N029N015P017(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='0' AND A( 1)='1' )then
          cVar1S26S20P011N029N015P017(0) <='1';
          else
          cVar1S26S20P011N029N015P017(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S27S20P011N029N015N017(0) <='1';
          else
          cVar1S27S20P011N029N015N017(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND A( 2)='0' AND A( 1)='0' )then
          cVar1S28S20P011N029N015N017(0) <='1';
          else
          cVar1S28S20P011N029N015N017(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' )then
          cVar1S0S21P041P020nsss(0) <='1';
          else
          cVar1S0S21P041P020nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='1' AND A( 8)='1' )then
          cVar1S1S21P041N020P021P003nsss(0) <='1';
          else
          cVar1S1S21P041N020P021P003nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='1' AND A( 8)='0' )then
          cVar1S2S21P041N020P021N003(0) <='1';
          else
          cVar1S2S21P041N020P021N003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND A(17)='1' )then
          cVar1S3S21P041N020N021P004nsss(0) <='1';
          else
          cVar1S3S21P041N020N021P004nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND A(17)='0' )then
          cVar1S4S21P041N020N021N004(0) <='1';
          else
          cVar1S4S21P041N020N021N004(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND A(17)='0' )then
          cVar1S5S21P041N020N021N004(0) <='1';
          else
          cVar1S5S21P041N020N021N004(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND B( 9)='0' AND A(17)='0' )then
          cVar1S6S21P041N020N021N004(0) <='1';
          else
          cVar1S6S21P041N020N021N004(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='1' )then
          cVar1S7S21N041P039P000P048(0) <='1';
          else
          cVar1S7S21N041P039P000P048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='1' )then
          cVar1S8S21N041P039P000P048(0) <='1';
          else
          cVar1S8S21N041P039P000P048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='1' )then
          cVar1S9S21N041P039P000P048(0) <='1';
          else
          cVar1S9S21N041P039P000P048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='0' )then
          cVar1S10S21N041P039P000N048(0) <='1';
          else
          cVar1S10S21N041P039P000N048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='0' )then
          cVar1S11S21N041P039P000N048(0) <='1';
          else
          cVar1S11S21N041P039P000N048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='0' AND D( 5)='0' )then
          cVar1S12S21N041P039P000N048(0) <='1';
          else
          cVar1S12S21N041P039P000N048(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='1' AND D( 7)='1' )then
          cVar1S13S21N041P039P000P040nsss(0) <='1';
          else
          cVar1S13S21N041P039P000P040nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='1' AND D( 7)='0' )then
          cVar1S14S21N041P039P000N040(0) <='1';
          else
          cVar1S14S21N041P039P000N040(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND A(19)='1' AND D( 7)='0' )then
          cVar1S15S21N041P039P000N040(0) <='1';
          else
          cVar1S15S21N041P039P000N040(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND E(13)='1' )then
          cVar1S16S21N041P039P051nsss(0) <='1';
          else
          cVar1S16S21N041P039P051nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND E(13)='0' AND B(19)='1' )then
          cVar1S17S21N041P039N051P020nsss(0) <='1';
          else
          cVar1S17S21N041P039N051P020nsss(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='1' AND B( 0)='1' )then
          cVar1S0S22P000P041P020P039nsss(0) <='1';
          else
          cVar1S0S22P000P041P020P039nsss(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S1S22P000P041N020P005(0) <='1';
          else
          cVar1S1S22P000P041N020P005(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S2S22P000P041N020P005(0) <='1';
          else
          cVar1S2S22P000P041N020P005(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S3S22P000P041N020N005(0) <='1';
          else
          cVar1S3S22P000P041N020N005(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S4S22P000P041N020N005(0) <='1';
          else
          cVar1S4S22P000P041N020N005(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S5S22P000P041N020N005(0) <='1';
          else
          cVar1S5S22P000P041N020N005(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='0' )then
          cVar1S6S22P000N041P039P012(0) <='1';
          else
          cVar1S6S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='0' )then
          cVar1S7S22P000N041P039P012(0) <='1';
          else
          cVar1S7S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='0' )then
          cVar1S8S22P000N041P039P012(0) <='1';
          else
          cVar1S8S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='1' )then
          cVar1S9S22P000N041P039P012(0) <='1';
          else
          cVar1S9S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='1' )then
          cVar1S10S22P000N041P039P012(0) <='1';
          else
          cVar1S10S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='0' AND A(13)='1' )then
          cVar1S11S22P000N041P039P012(0) <='1';
          else
          cVar1S11S22P000N041P039P012(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='1' )then
          cVar1S12S22P000N041P039P049nsss(0) <='1';
          else
          cVar1S12S22P000N041P039P049nsss(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='0' )then
          cVar1S13S22P000N041P039N049(0) <='1';
          else
          cVar1S13S22P000N041P039N049(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='0' )then
          cVar1S14S22P000N041P039N049(0) <='1';
          else
          cVar1S14S22P000N041P039N049(0) <='0';
          end if;
        if(A(19)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='0' )then
          cVar1S15S22P000N041P039N049(0) <='1';
          else
          cVar1S15S22P000N041P039N049(0) <='0';
          end if;
        if(A(19)='1' AND D( 7)='1' )then
          cVar1S16S22P000P040nsss(0) <='1';
          else
          cVar1S16S22P000P040nsss(0) <='0';
          end if;
        if(A(19)='1' AND D( 7)='0' AND E(11)='0' AND D(15)='1' )then
          cVar1S17S22P000N040P059P041nsss(0) <='1';
          else
          cVar1S17S22P000N040P059P041nsss(0) <='0';
          end if;
        if(A(19)='1' AND D( 7)='0' AND E(11)='0' AND D(15)='0' )then
          cVar1S18S22P000N040P059N041(0) <='1';
          else
          cVar1S18S22P000N040P059N041(0) <='0';
          end if;
        if(A(19)='1' AND D( 7)='0' AND E(11)='0' AND D(15)='0' )then
          cVar1S19S22P000N040P059N041(0) <='1';
          else
          cVar1S19S22P000N040P059N041(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A(14)='0' )then
          cVar1S0S23P041P020P010nsss(0) <='1';
          else
          cVar1S0S23P041P020P010nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='1' )then
          cVar1S1S23P041N020P005P021nsss(0) <='1';
          else
          cVar1S1S23P041N020P005P021nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='0' )then
          cVar1S2S23P041N020P005N021(0) <='1';
          else
          cVar1S2S23P041N020P005N021(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='0' )then
          cVar1S3S23P041N020P005N021(0) <='1';
          else
          cVar1S3S23P041N020P005N021(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='1' )then
          cVar1S4S23P041N020N005P003(0) <='1';
          else
          cVar1S4S23P041N020N005P003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S5S23P041N020N005N003(0) <='1';
          else
          cVar1S5S23P041N020N005N003(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='0' AND D( 3)='0' )then
          cVar1S6S23N041P055P061P056(0) <='1';
          else
          cVar1S6S23N041P055P061P056(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='0' AND D( 3)='0' )then
          cVar1S7S23N041P055P061P056(0) <='1';
          else
          cVar1S7S23N041P055P061P056(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='0' AND D( 3)='0' )then
          cVar1S8S23N041P055P061P056(0) <='1';
          else
          cVar1S8S23N041P055P061P056(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='0' AND D( 3)='1' )then
          cVar1S9S23N041P055P061P056(0) <='1';
          else
          cVar1S9S23N041P055P061P056(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='1' AND E( 4)='1' )then
          cVar1S10S23N041P055P061P054nsss(0) <='1';
          else
          cVar1S10S23N041P055P061P054nsss(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='1' AND D(10)='1' AND E( 4)='0' )then
          cVar1S11S23N041P055P061N054(0) <='1';
          else
          cVar1S11S23N041P055P061N054(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='0' AND B( 0)='0' )then
          cVar1S12S23N041N055P010P039(0) <='1';
          else
          cVar1S12S23N041N055P010P039(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='0' AND B( 0)='0' )then
          cVar1S13S23N041N055P010P039(0) <='1';
          else
          cVar1S13S23N041N055P010P039(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='0' AND B( 0)='0' )then
          cVar1S14S23N041N055P010P039(0) <='1';
          else
          cVar1S14S23N041N055P010P039(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='0' AND B( 0)='0' )then
          cVar1S15S23N041N055P010P039(0) <='1';
          else
          cVar1S15S23N041N055P010P039(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='0' AND B( 0)='1' )then
          cVar1S16S23N041N055P010P039(0) <='1';
          else
          cVar1S16S23N041N055P010P039(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='1' AND B(15)='1' )then
          cVar1S17S23N041N055P010P028(0) <='1';
          else
          cVar1S17S23N041N055P010P028(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='1' AND B(15)='0' )then
          cVar1S18S23N041N055P010N028(0) <='1';
          else
          cVar1S18S23N041N055P010N028(0) <='0';
          end if;
        if(D(15)='0' AND E(12)='0' AND A(14)='1' AND B(15)='0' )then
          cVar1S19S23N041N055P010N028(0) <='1';
          else
          cVar1S19S23N041N055P010N028(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND B( 0)='1' )then
          cVar1S0S24P041P020P039nsss(0) <='1';
          else
          cVar1S0S24P041P020P039nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='1' )then
          cVar1S1S24P041N020P005P021nsss(0) <='1';
          else
          cVar1S1S24P041N020P005P021nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='0' )then
          cVar1S2S24P041N020P005N021(0) <='1';
          else
          cVar1S2S24P041N020P005N021(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='0' )then
          cVar1S3S24P041N020P005N021(0) <='1';
          else
          cVar1S3S24P041N020P005N021(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='1' )then
          cVar1S4S24P041N020N005P003(0) <='1';
          else
          cVar1S4S24P041N020N005P003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S5S24P041N020N005N003(0) <='1';
          else
          cVar1S5S24P041N020N005N003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S6S24P041N020N005N003(0) <='1';
          else
          cVar1S6S24P041N020N005N003(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S7S24N041P039P058P033(0) <='1';
          else
          cVar1S7S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S8S24N041P039P058P033(0) <='1';
          else
          cVar1S8S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S9S24N041P039P058P033(0) <='1';
          else
          cVar1S9S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S10S24N041P039P058P033(0) <='1';
          else
          cVar1S10S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='1' )then
          cVar1S11S24N041P039P058P033(0) <='1';
          else
          cVar1S11S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='1' )then
          cVar1S12S24N041P039P058P033(0) <='1';
          else
          cVar1S12S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='0' AND B( 3)='1' )then
          cVar1S13S24N041P039P058P033(0) <='1';
          else
          cVar1S13S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='1' AND B( 3)='1' )then
          cVar1S14S24N041P039P058P033(0) <='1';
          else
          cVar1S14S24N041P039P058P033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S15S24N041P039P058N033(0) <='1';
          else
          cVar1S15S24N041P039P058N033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S16S24N041P039P058N033(0) <='1';
          else
          cVar1S16S24N041P039P058N033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S17S24N041P039P058N033(0) <='1';
          else
          cVar1S17S24N041P039P058N033(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND E(13)='1' )then
          cVar1S18S24N041P039P051nsss(0) <='1';
          else
          cVar1S18S24N041P039P051nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND E(13)='0' AND D( 1)='1' )then
          cVar1S19S24N041P039N051P064nsss(0) <='1';
          else
          cVar1S19S24N041P039N051P064nsss(0) <='0';
          end if;
        if(D(15)='0' AND B( 0)='1' AND E(13)='0' AND D( 1)='0' )then
          cVar1S20S24N041P039N051N064(0) <='1';
          else
          cVar1S20S24N041P039N051N064(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' )then
          cVar1S0S25P041P020nsss(0) <='1';
          else
          cVar1S0S25P041P020nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='1' )then
          cVar1S1S25P041N020P005P021nsss(0) <='1';
          else
          cVar1S1S25P041N020P005P021nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='1' AND B( 9)='0' )then
          cVar1S2S25P041N020P005N021(0) <='1';
          else
          cVar1S2S25P041N020P005N021(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='1' )then
          cVar1S3S25P041N020N005P003(0) <='1';
          else
          cVar1S3S25P041N020N005P003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S4S25P041N020N005N003(0) <='1';
          else
          cVar1S4S25P041N020N005N003(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S5S25P041N020N005N003(0) <='1';
          else
          cVar1S5S25P041N020N005N003(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='1' AND D( 3)='1' )then
          cVar1S6S25N041P013P031P056(0) <='1';
          else
          cVar1S6S25N041P013P031P056(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='1' AND D( 3)='1' )then
          cVar1S7S25N041P013P031P056(0) <='1';
          else
          cVar1S7S25N041P013P031P056(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='1' AND D( 3)='0' )then
          cVar1S8S25N041P013P031N056(0) <='1';
          else
          cVar1S8S25N041P013P031N056(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='1' AND D( 3)='0' )then
          cVar1S9S25N041P013P031N056(0) <='1';
          else
          cVar1S9S25N041P013P031N056(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='0' AND A( 2)='1' )then
          cVar1S10S25N041P013N031P015(0) <='1';
          else
          cVar1S10S25N041P013N031P015(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='0' AND A( 2)='1' )then
          cVar1S11S25N041P013N031P015(0) <='1';
          else
          cVar1S11S25N041P013N031P015(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='0' AND A( 2)='1' )then
          cVar1S12S25N041P013N031P015(0) <='1';
          else
          cVar1S12S25N041P013N031P015(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='0' AND A( 2)='0' )then
          cVar1S13S25N041P013N031N015(0) <='1';
          else
          cVar1S13S25N041P013N031N015(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='1' AND B( 4)='0' AND A( 2)='0' )then
          cVar1S14S25N041P013N031N015(0) <='1';
          else
          cVar1S14S25N041P013N031N015(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='0' AND D( 6)='1' )then
          cVar1S15S25N041N013P031P044(0) <='1';
          else
          cVar1S15S25N041N013P031P044(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='0' AND D( 6)='1' )then
          cVar1S16S25N041N013P031P044(0) <='1';
          else
          cVar1S16S25N041N013P031P044(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='0' AND D( 6)='0' )then
          cVar1S17S25N041N013P031N044(0) <='1';
          else
          cVar1S17S25N041N013P031N044(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='0' AND D( 6)='0' )then
          cVar1S18S25N041N013P031N044(0) <='1';
          else
          cVar1S18S25N041N013P031N044(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='0' AND D( 6)='0' )then
          cVar1S19S25N041N013P031N044(0) <='1';
          else
          cVar1S19S25N041N013P031N044(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='1' AND A( 4)='1' )then
          cVar1S20S25N041N013P031P011(0) <='1';
          else
          cVar1S20S25N041N013P031P011(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='1' AND A( 4)='1' )then
          cVar1S21S25N041N013P031P011(0) <='1';
          else
          cVar1S21S25N041N013P031P011(0) <='0';
          end if;
        if(D(15)='0' AND A( 3)='0' AND B( 4)='1' AND A( 4)='0' )then
          cVar1S22S25N041N013P031N011(0) <='1';
          else
          cVar1S22S25N041N013P031N011(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='1' AND B(19)='1' AND A(11)='0' )then
          cVar1S0S26P068P041P020P016nsss(0) <='1';
          else
          cVar1S0S26P068P041P020P016nsss(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S1S26P068P041N020P005(0) <='1';
          else
          cVar1S1S26P068P041N020P005(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S2S26P068P041N020P005(0) <='1';
          else
          cVar1S2S26P068P041N020P005(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S3S26P068P041N020N005(0) <='1';
          else
          cVar1S3S26P068P041N020N005(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S4S26P068P041N020N005(0) <='1';
          else
          cVar1S4S26P068P041N020N005(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S5S26P068N041P024P006(0) <='1';
          else
          cVar1S5S26P068N041P024P006(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S6S26P068N041P024P006(0) <='1';
          else
          cVar1S6S26P068N041P024P006(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S7S26P068N041P024P006(0) <='1';
          else
          cVar1S7S26P068N041P024P006(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='1' AND A(16)='0' )then
          cVar1S8S26P068N041P024N006(0) <='1';
          else
          cVar1S8S26P068N041P024N006(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='1' AND A(16)='0' )then
          cVar1S9S26P068N041P024N006(0) <='1';
          else
          cVar1S9S26P068N041P024N006(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='1' )then
          cVar1S10S26P068N041N024P023(0) <='1';
          else
          cVar1S10S26P068N041N024P023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='1' )then
          cVar1S11S26P068N041N024P023(0) <='1';
          else
          cVar1S11S26P068N041N024P023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='1' )then
          cVar1S12S26P068N041N024P023(0) <='1';
          else
          cVar1S12S26P068N041N024P023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='1' )then
          cVar1S13S26P068N041N024P023(0) <='1';
          else
          cVar1S13S26P068N041N024P023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='0' )then
          cVar1S14S26P068N041N024N023(0) <='1';
          else
          cVar1S14S26P068N041N024N023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='0' )then
          cVar1S15S26P068N041N024N023(0) <='1';
          else
          cVar1S15S26P068N041N024N023(0) <='0';
          end if;
        if(D( 0)='0' AND D(15)='0' AND B(17)='0' AND B( 8)='0' )then
          cVar1S16S26P068N041N024N023(0) <='1';
          else
          cVar1S16S26P068N041N024N023(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='1' AND D(10)='0' )then
          cVar1S17S26P068P065P019P061(0) <='1';
          else
          cVar1S17S26P068P065P019P061(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='1' AND D(10)='0' )then
          cVar1S18S26P068P065P019P061(0) <='1';
          else
          cVar1S18S26P068P065P019P061(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='1' )then
          cVar1S19S26P068P065N019P037(0) <='1';
          else
          cVar1S19S26P068P065N019P037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='1' )then
          cVar1S20S26P068P065N019P037(0) <='1';
          else
          cVar1S20S26P068P065N019P037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='1' )then
          cVar1S21S26P068P065N019P037(0) <='1';
          else
          cVar1S21S26P068P065N019P037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='0' )then
          cVar1S22S26P068P065N019N037(0) <='1';
          else
          cVar1S22S26P068P065N019N037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='0' )then
          cVar1S23S26P068P065N019N037(0) <='1';
          else
          cVar1S23S26P068P065N019N037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='0' AND A( 0)='0' AND B( 1)='0' )then
          cVar1S24S26P068P065N019N037(0) <='1';
          else
          cVar1S24S26P068P065N019N037(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='1' AND B(11)='0' )then
          cVar1S25S26P068P065P069P036(0) <='1';
          else
          cVar1S25S26P068P065P069P036(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='1' AND B(11)='0' )then
          cVar1S26S26P068P065P069P036(0) <='1';
          else
          cVar1S26S26P068P065P069P036(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='1' AND B(11)='1' )then
          cVar1S27S26P068P065P069P036(0) <='1';
          else
          cVar1S27S26P068P065P069P036(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='0' AND A(11)='1' )then
          cVar1S28S26P068P065N069P016(0) <='1';
          else
          cVar1S28S26P068P065N069P016(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='0' AND A(11)='1' )then
          cVar1S29S26P068P065N069P016(0) <='1';
          else
          cVar1S29S26P068P065N069P016(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='0' AND A(11)='0' )then
          cVar1S30S26P068P065N069N016(0) <='1';
          else
          cVar1S30S26P068P065N069N016(0) <='0';
          end if;
        if(D( 0)='1' AND D( 9)='1' AND D( 8)='0' AND A(11)='0' )then
          cVar1S31S26P068P065N069N016(0) <='1';
          else
          cVar1S31S26P068P065N069N016(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S0S27P041P020P003nsss(0) <='1';
          else
          cVar1S0S27P041P020P003nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='1' )then
          cVar1S1S27P041P020N003P002nsss(0) <='1';
          else
          cVar1S1S27P041P020N003P002nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='0' )then
          cVar1S2S27P041P020N003N002(0) <='1';
          else
          cVar1S2S27P041P020N003N002(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='0' )then
          cVar1S3S27P041P020N003N002(0) <='1';
          else
          cVar1S3S27P041P020N003N002(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND D( 0)='0' AND A( 7)='1' )then
          cVar1S4S27P041N020P068P005(0) <='1';
          else
          cVar1S4S27P041N020P068P005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND D( 0)='0' AND A( 7)='1' )then
          cVar1S5S27P041N020P068P005(0) <='1';
          else
          cVar1S5S27P041N020P068P005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND D( 0)='0' AND A( 7)='0' )then
          cVar1S6S27P041N020P068N005(0) <='1';
          else
          cVar1S6S27P041N020P068N005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND D( 0)='1' AND B( 0)='0' )then
          cVar1S7S27P041N020P068P039(0) <='1';
          else
          cVar1S7S27P041N020P068P039(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='1' AND E(14)='1' )then
          cVar1S8S27N041P024P006P047nsss(0) <='1';
          else
          cVar1S8S27N041P024P006P047nsss(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='1' AND E(14)='0' )then
          cVar1S9S27N041P024P006N047(0) <='1';
          else
          cVar1S9S27N041P024P006N047(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='1' AND E(14)='0' )then
          cVar1S10S27N041P024P006N047(0) <='1';
          else
          cVar1S10S27N041P024P006N047(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='1' AND E(14)='0' )then
          cVar1S11S27N041P024P006N047(0) <='1';
          else
          cVar1S11S27N041P024P006N047(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='0' AND D(13)='1' )then
          cVar1S12S27N041P024N006P049(0) <='1';
          else
          cVar1S12S27N041P024N006P049(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='0' AND D(13)='1' )then
          cVar1S13S27N041P024N006P049(0) <='1';
          else
          cVar1S13S27N041P024N006P049(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='0' AND D(13)='0' )then
          cVar1S14S27N041P024N006N049(0) <='1';
          else
          cVar1S14S27N041P024N006N049(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='1' AND A(16)='0' AND D(13)='0' )then
          cVar1S15S27N041P024N006N049(0) <='1';
          else
          cVar1S15S27N041P024N006N049(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S16S27N041N024P023P005(0) <='1';
          else
          cVar1S16S27N041N024P023P005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S17S27N041N024P023P005(0) <='1';
          else
          cVar1S17S27N041N024P023P005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S18S27N041N024P023N005(0) <='1';
          else
          cVar1S18S27N041N024P023N005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S19S27N041N024P023N005(0) <='1';
          else
          cVar1S19S27N041N024P023N005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S20S27N041N024P023N005(0) <='1';
          else
          cVar1S20S27N041N024P023N005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S21S27N041N024P023N005(0) <='1';
          else
          cVar1S21S27N041N024P023N005(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='1' )then
          cVar1S22S27N041N024N023P050(0) <='1';
          else
          cVar1S22S27N041N024N023P050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='1' )then
          cVar1S23S27N041N024N023P050(0) <='1';
          else
          cVar1S23S27N041N024N023P050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='1' )then
          cVar1S24S27N041N024N023P050(0) <='1';
          else
          cVar1S24S27N041N024N023P050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='1' )then
          cVar1S25S27N041N024N023P050(0) <='1';
          else
          cVar1S25S27N041N024N023P050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='0' )then
          cVar1S26S27N041N024N023N050(0) <='1';
          else
          cVar1S26S27N041N024N023N050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='0' )then
          cVar1S27S27N041N024N023N050(0) <='1';
          else
          cVar1S27S27N041N024N023N050(0) <='0';
          end if;
        if(D(15)='0' AND B(17)='0' AND B( 8)='0' AND E( 5)='0' )then
          cVar1S28S27N041N024N023N050(0) <='1';
          else
          cVar1S28S27N041N024N023N050(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='1' )then
          cVar1S0S28P024P006P047nsss(0) <='1';
          else
          cVar1S0S28P024P006P047nsss(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='1' )then
          cVar1S1S28P024P006N047P045nsss(0) <='1';
          else
          cVar1S1S28P024P006N047P045nsss(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='0' )then
          cVar1S2S28P024P006N047N045(0) <='1';
          else
          cVar1S2S28P024P006N047N045(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='0' )then
          cVar1S3S28P024P006N047N045(0) <='1';
          else
          cVar1S3S28P024P006N047N045(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND B(12)='0' )then
          cVar1S4S28P024N006P068P034(0) <='1';
          else
          cVar1S4S28P024N006P068P034(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND B(12)='0' )then
          cVar1S5S28P024N006P068P034(0) <='1';
          else
          cVar1S5S28P024N006P068P034(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND B(12)='1' )then
          cVar1S6S28P024N006P068P034(0) <='1';
          else
          cVar1S6S28P024N006P068P034(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='1' AND E(14)='1' )then
          cVar1S7S28P024N006P068P047nsss(0) <='1';
          else
          cVar1S7S28P024N006P068P047nsss(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S8S28N024P040P002nsss(0) <='1';
          else
          cVar1S8S28N024P040P002nsss(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S9S28N024P040N002P004nsss(0) <='1';
          else
          cVar1S9S28N024P040N002P004nsss(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S10S28N024P040N002N004(0) <='1';
          else
          cVar1S10S28N024P040N002N004(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S11S28N024P040N002N004(0) <='1';
          else
          cVar1S11S28N024P040N002N004(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S12S28N024N040P044P023(0) <='1';
          else
          cVar1S12S28N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S13S28N024N040P044P023(0) <='1';
          else
          cVar1S13S28N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S14S28N024N040P044P023(0) <='1';
          else
          cVar1S14S28N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S15S28N024N040P044N023(0) <='1';
          else
          cVar1S15S28N024N040P044N023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S16S28N024N040P044N023(0) <='1';
          else
          cVar1S16S28N024N040P044N023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S17S28N024N040P044N023(0) <='1';
          else
          cVar1S17S28N024N040P044N023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND E( 7)='0' )then
          cVar1S18S28N024N040N044P042(0) <='1';
          else
          cVar1S18S28N024N040N044P042(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND E( 7)='0' )then
          cVar1S19S28N024N040N044P042(0) <='1';
          else
          cVar1S19S28N024N040N044P042(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND E( 7)='0' )then
          cVar1S20S28N024N040N044P042(0) <='1';
          else
          cVar1S20S28N024N040N044P042(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND E( 7)='1' )then
          cVar1S21S28N024N040N044P042(0) <='1';
          else
          cVar1S21S28N024N040N044P042(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND E( 7)='1' )then
          cVar1S22S28N024N040N044P042(0) <='1';
          else
          cVar1S22S28N024N040N044P042(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='1' )then
          cVar1S0S29P024P006P047nsss(0) <='1';
          else
          cVar1S0S29P024P006P047nsss(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='1' )then
          cVar1S1S29P024P006N047P045nsss(0) <='1';
          else
          cVar1S1S29P024P006N047P045nsss(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='0' )then
          cVar1S2S29P024P006N047N045(0) <='1';
          else
          cVar1S2S29P024P006N047N045(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='1' AND E(14)='0' AND D(14)='0' )then
          cVar1S3S29P024P006N047N045(0) <='1';
          else
          cVar1S3S29P024P006N047N045(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND A( 6)='1' )then
          cVar1S4S29P024N006P068P007(0) <='1';
          else
          cVar1S4S29P024N006P068P007(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND A( 6)='1' )then
          cVar1S5S29P024N006P068P007(0) <='1';
          else
          cVar1S5S29P024N006P068P007(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='0' AND A( 6)='0' )then
          cVar1S6S29P024N006P068N007(0) <='1';
          else
          cVar1S6S29P024N006P068N007(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='1' AND A(13)='1' )then
          cVar1S7S29P024N006P068P012nsss(0) <='1';
          else
          cVar1S7S29P024N006P068P012nsss(0) <='0';
          end if;
        if(B(17)='1' AND A(16)='0' AND D( 0)='1' AND A(13)='0' )then
          cVar1S8S29P024N006P068N012(0) <='1';
          else
          cVar1S8S29P024N006P068N012(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S9S29N024P040P002nsss(0) <='1';
          else
          cVar1S9S29N024P040P002nsss(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S10S29N024P040N002P034(0) <='1';
          else
          cVar1S10S29N024P040N002P034(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S11S29N024P040N002P034(0) <='1';
          else
          cVar1S11S29N024P040N002P034(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S12S29N024P040N002P034(0) <='1';
          else
          cVar1S12S29N024P040N002P034(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S13S29N024P040N002P034(0) <='1';
          else
          cVar1S13S29N024P040N002P034(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S14S29N024N040P044P023(0) <='1';
          else
          cVar1S14S29N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S15S29N024N040P044P023(0) <='1';
          else
          cVar1S15S29N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S16S29N024N040P044P023(0) <='1';
          else
          cVar1S16S29N024N040P044P023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S17S29N024N040P044N023(0) <='1';
          else
          cVar1S17S29N024N040P044N023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S18S29N024N040P044N023(0) <='1';
          else
          cVar1S18S29N024N040P044N023(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND D(15)='1' )then
          cVar1S19S29N024N040N044P041(0) <='1';
          else
          cVar1S19S29N024N040N044P041(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND D(15)='1' )then
          cVar1S20S29N024N040N044P041(0) <='1';
          else
          cVar1S20S29N024N040N044P041(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND D(15)='1' )then
          cVar1S21S29N024N040N044P041(0) <='1';
          else
          cVar1S21S29N024N040N044P041(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND D(15)='1' )then
          cVar1S22S29N024N040N044P041(0) <='1';
          else
          cVar1S22S29N024N040N044P041(0) <='0';
          end if;
        if(B(17)='0' AND D( 7)='0' AND D( 6)='0' AND D(15)='0' )then
          cVar1S23S29N024N040N044N041(0) <='1';
          else
          cVar1S23S29N024N040N044N041(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S0S30P067P018P048P025nsss(0) <='1';
          else
          cVar1S0S30P067P018P048P025nsss(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='1' AND B( 7)='0' )then
          cVar1S1S30P067P018P048N025(0) <='1';
          else
          cVar1S1S30P067P018P048N025(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='1' AND B( 7)='0' )then
          cVar1S2S30P067P018P048N025(0) <='1';
          else
          cVar1S2S30P067P018P048N025(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='1' AND B( 7)='0' )then
          cVar1S3S30P067P018P048N025(0) <='1';
          else
          cVar1S3S30P067P018P048N025(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='1' )then
          cVar1S4S30P067P018N048P014(0) <='1';
          else
          cVar1S4S30P067P018N048P014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='1' )then
          cVar1S5S30P067P018N048P014(0) <='1';
          else
          cVar1S5S30P067P018N048P014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='1' )then
          cVar1S6S30P067P018N048P014(0) <='1';
          else
          cVar1S6S30P067P018N048P014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='1' )then
          cVar1S7S30P067P018N048P014(0) <='1';
          else
          cVar1S7S30P067P018N048P014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='0' )then
          cVar1S8S30P067P018N048N014(0) <='1';
          else
          cVar1S8S30P067P018N048N014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='0' AND D( 5)='0' AND A(12)='0' )then
          cVar1S9S30P067P018N048N014(0) <='1';
          else
          cVar1S9S30P067P018N048N014(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S10S30P067P018P060P011(0) <='1';
          else
          cVar1S10S30P067P018P060P011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S11S30P067P018P060P011(0) <='1';
          else
          cVar1S11S30P067P018P060P011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='1' )then
          cVar1S12S30P067P018P060P011(0) <='1';
          else
          cVar1S12S30P067P018P060P011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S13S30P067P018P060N011(0) <='1';
          else
          cVar1S13S30P067P018P060N011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S14S30P067P018P060N011(0) <='1';
          else
          cVar1S14S30P067P018P060N011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='0' AND A( 4)='0' )then
          cVar1S15S30P067P018P060N011(0) <='1';
          else
          cVar1S15S30P067P018P060N011(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='1' AND A( 3)='1' )then
          cVar1S16S30P067P018P060P013(0) <='1';
          else
          cVar1S16S30P067P018P060P013(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='1' AND A( 3)='1' )then
          cVar1S17S30P067P018P060P013(0) <='1';
          else
          cVar1S17S30P067P018P060P013(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='1' AND A( 3)='0' )then
          cVar1S18S30P067P018P060N013(0) <='1';
          else
          cVar1S18S30P067P018P060N013(0) <='0';
          end if;
        if(E( 9)='0' AND A(10)='1' AND D( 2)='1' AND A( 3)='0' )then
          cVar1S19S30P067P018P060N013(0) <='1';
          else
          cVar1S19S30P067P018P060N013(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(11)='0' )then
          cVar1S20S30P067P069P018P016(0) <='1';
          else
          cVar1S20S30P067P069P018P016(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(11)='0' )then
          cVar1S21S30P067P069P018P016(0) <='1';
          else
          cVar1S21S30P067P069P018P016(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(11)='0' )then
          cVar1S22S30P067P069P018P016(0) <='1';
          else
          cVar1S22S30P067P069P018P016(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='1' AND A(11)='1' )then
          cVar1S23S30P067P069P018P016(0) <='1';
          else
          cVar1S23S30P067P069P018P016(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar1S24S30P067P069N018P019(0) <='1';
          else
          cVar1S24S30P067P069N018P019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='1' )then
          cVar1S25S30P067P069N018P019(0) <='1';
          else
          cVar1S25S30P067P069N018P019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S26S30P067P069N018N019(0) <='1';
          else
          cVar1S26S30P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S27S30P067P069N018N019(0) <='1';
          else
          cVar1S27S30P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='1' AND A(10)='0' AND A( 0)='0' )then
          cVar1S28S30P067P069N018N019(0) <='1';
          else
          cVar1S28S30P067P069N018N019(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 9)='1' AND E(10)='0' )then
          cVar1S29S30P067N069P065P063nsss(0) <='1';
          else
          cVar1S29S30P067N069P065P063nsss(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 9)='1' AND E(10)='1' )then
          cVar1S30S30P067N069P065P063(0) <='1';
          else
          cVar1S30S30P067N069P065P063(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 9)='0' AND D( 4)='1' )then
          cVar1S31S30P067N069N065P052nsss(0) <='1';
          else
          cVar1S31S30P067N069N065P052nsss(0) <='0';
          end if;
        if(E( 9)='1' AND D( 8)='0' AND D( 9)='0' AND D( 4)='0' )then
          cVar1S32S30P067N069N065N052(0) <='1';
          else
          cVar1S32S30P067N069N065N052(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='0' )then
          cVar1S0S31P018P060P054P062(0) <='1';
          else
          cVar1S0S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='0' )then
          cVar1S1S31P018P060P054P062(0) <='1';
          else
          cVar1S1S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='0' )then
          cVar1S2S31P018P060P054P062(0) <='1';
          else
          cVar1S2S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='1' )then
          cVar1S3S31P018P060P054P062(0) <='1';
          else
          cVar1S3S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='1' )then
          cVar1S4S31P018P060P054P062(0) <='1';
          else
          cVar1S4S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='0' AND E( 2)='1' )then
          cVar1S5S31P018P060P054P062(0) <='1';
          else
          cVar1S5S31P018P060P054P062(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='1' AND A( 4)='1' )then
          cVar1S6S31P018P060P054P011(0) <='1';
          else
          cVar1S6S31P018P060P054P011(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='0' AND E( 4)='1' AND A( 4)='0' )then
          cVar1S7S31P018P060P054N011(0) <='1';
          else
          cVar1S7S31P018P060P054N011(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='1' AND B( 5)='0' AND E( 5)='1' )then
          cVar1S8S31P018P060P029P050nsss(0) <='1';
          else
          cVar1S8S31P018P060P029P050nsss(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='1' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S9S31P018P060P029N050(0) <='1';
          else
          cVar1S9S31P018P060P029N050(0) <='0';
          end if;
        if(A(10)='1' AND D( 2)='1' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S10S31P018P060P029N050(0) <='1';
          else
          cVar1S10S31P018P060P029N050(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S11S31N018P048P025P007nsss(0) <='1';
          else
          cVar1S11S31N018P048P025P007nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S12S31N018P048P025N007(0) <='1';
          else
          cVar1S12S31N018P048P025N007(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S13S31N018P048P025N007(0) <='1';
          else
          cVar1S13S31N018P048P025N007(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B(11)='0' )then
          cVar1S14S31N018P048N025P036nsss(0) <='1';
          else
          cVar1S14S31N018P048N025P036nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='1' AND B(12)='1' )then
          cVar1S15S31N018N048P014P034(0) <='1';
          else
          cVar1S15S31N018N048P014P034(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='1' AND B(12)='0' )then
          cVar1S16S31N018N048P014N034(0) <='1';
          else
          cVar1S16S31N018N048P014N034(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='1' AND B(12)='0' )then
          cVar1S17S31N018N048P014N034(0) <='1';
          else
          cVar1S17S31N018N048P014N034(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='1' AND B(12)='0' )then
          cVar1S18S31N018N048P014N034(0) <='1';
          else
          cVar1S18S31N018N048P014N034(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='1' )then
          cVar1S19S31N018N048N014P030(0) <='1';
          else
          cVar1S19S31N018N048N014P030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='1' )then
          cVar1S20S31N018N048N014P030(0) <='1';
          else
          cVar1S20S31N018N048N014P030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='1' )then
          cVar1S21S31N018N048N014P030(0) <='1';
          else
          cVar1S21S31N018N048N014P030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='1' )then
          cVar1S22S31N018N048N014P030(0) <='1';
          else
          cVar1S22S31N018N048N014P030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='0' )then
          cVar1S23S31N018N048N014N030(0) <='1';
          else
          cVar1S23S31N018N048N014N030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='0' )then
          cVar1S24S31N018N048N014N030(0) <='1';
          else
          cVar1S24S31N018N048N014N030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='0' )then
          cVar1S25S31N018N048N014N030(0) <='1';
          else
          cVar1S25S31N018N048N014N030(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(12)='0' AND B(14)='0' )then
          cVar1S26S31N018N048N014N030(0) <='1';
          else
          cVar1S26S31N018N048N014N030(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S0S32P015P018P040P021nsss(0) <='1';
          else
          cVar1S0S32P015P018P040P021nsss(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S1S32P015P018P040N021(0) <='1';
          else
          cVar1S1S32P015P018P040N021(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S2S32P015P018P040N021(0) <='1';
          else
          cVar1S2S32P015P018P040N021(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S3S32P015P018P040N021(0) <='1';
          else
          cVar1S3S32P015P018P040N021(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='1' )then
          cVar1S4S32P015P018N040P063(0) <='1';
          else
          cVar1S4S32P015P018N040P063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='1' )then
          cVar1S5S32P015P018N040P063(0) <='1';
          else
          cVar1S5S32P015P018N040P063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='1' )then
          cVar1S6S32P015P018N040P063(0) <='1';
          else
          cVar1S6S32P015P018N040P063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='1' )then
          cVar1S7S32P015P018N040P063(0) <='1';
          else
          cVar1S7S32P015P018N040P063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='0' )then
          cVar1S8S32P015P018N040N063(0) <='1';
          else
          cVar1S8S32P015P018N040N063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='0' )then
          cVar1S9S32P015P018N040N063(0) <='1';
          else
          cVar1S9S32P015P018N040N063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='0' )then
          cVar1S10S32P015P018N040N063(0) <='1';
          else
          cVar1S10S32P015P018N040N063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='0' AND D( 7)='0' AND E(10)='0' )then
          cVar1S11S32P015P018N040N063(0) <='1';
          else
          cVar1S11S32P015P018N040N063(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='0' )then
          cVar1S12S32P015P018P004P062(0) <='1';
          else
          cVar1S12S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='0' )then
          cVar1S13S32P015P018P004P062(0) <='1';
          else
          cVar1S13S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='0' )then
          cVar1S14S32P015P018P004P062(0) <='1';
          else
          cVar1S14S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='0' )then
          cVar1S15S32P015P018P004P062(0) <='1';
          else
          cVar1S15S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='1' )then
          cVar1S16S32P015P018P004P062(0) <='1';
          else
          cVar1S16S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='0' AND E( 2)='1' )then
          cVar1S17S32P015P018P004P062(0) <='1';
          else
          cVar1S17S32P015P018P004P062(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='1' AND D(15)='1' )then
          cVar1S18S32P015P018P004P041nsss(0) <='1';
          else
          cVar1S18S32P015P018P004P041nsss(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='1' AND D(15)='0' )then
          cVar1S19S32P015P018P004N041(0) <='1';
          else
          cVar1S19S32P015P018P004N041(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='1' AND D(15)='0' )then
          cVar1S20S32P015P018P004N041(0) <='1';
          else
          cVar1S20S32P015P018P004N041(0) <='0';
          end if;
        if(A( 2)='0' AND A(10)='1' AND A(17)='1' AND D(15)='0' )then
          cVar1S21S32P015P018P004N041(0) <='1';
          else
          cVar1S21S32P015P018P004N041(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='1' AND E(10)='0' )then
          cVar1S22S32P015P017P060P063(0) <='1';
          else
          cVar1S22S32P015P017P060P063(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='1' AND E(10)='0' )then
          cVar1S23S32P015P017P060P063(0) <='1';
          else
          cVar1S23S32P015P017P060P063(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='1' AND E(10)='0' )then
          cVar1S24S32P015P017P060P063(0) <='1';
          else
          cVar1S24S32P015P017P060P063(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='1' AND E(10)='0' )then
          cVar1S25S32P015P017P060P063(0) <='1';
          else
          cVar1S25S32P015P017P060P063(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='1' )then
          cVar1S26S32P015P017N060P018(0) <='1';
          else
          cVar1S26S32P015P017N060P018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='1' )then
          cVar1S27S32P015P017N060P018(0) <='1';
          else
          cVar1S27S32P015P017N060P018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='0' )then
          cVar1S28S32P015P017N060N018(0) <='1';
          else
          cVar1S28S32P015P017N060N018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='0' )then
          cVar1S29S32P015P017N060N018(0) <='1';
          else
          cVar1S29S32P015P017N060N018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='0' )then
          cVar1S30S32P015P017N060N018(0) <='1';
          else
          cVar1S30S32P015P017N060N018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND D( 2)='0' AND A(10)='0' )then
          cVar1S31S32P015P017N060N018(0) <='1';
          else
          cVar1S31S32P015P017N060N018(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(15)='1' AND E( 1)='0' )then
          cVar1S32S32P015P017P008P066nsss(0) <='1';
          else
          cVar1S32S32P015P017P008P066nsss(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(15)='1' AND E( 1)='1' )then
          cVar1S33S32P015P017P008P066(0) <='1';
          else
          cVar1S33S32P015P017P008P066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(15)='0' AND D( 3)='0' )then
          cVar1S34S32P015P017N008P056(0) <='1';
          else
          cVar1S34S32P015P017N008P056(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(15)='0' AND D( 3)='0' )then
          cVar1S35S32P015P017N008P056(0) <='1';
          else
          cVar1S35S32P015P017N008P056(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND A(15)='0' AND D( 3)='1' )then
          cVar1S36S32P015P017N008P056(0) <='1';
          else
          cVar1S36S32P015P017N008P056(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='0' AND E(11)='0' )then
          cVar1S0S33P016P063P056P059(0) <='1';
          else
          cVar1S0S33P016P063P056P059(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='0' AND E(11)='0' )then
          cVar1S1S33P016P063P056P059(0) <='1';
          else
          cVar1S1S33P016P063P056P059(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='0' AND E(11)='0' )then
          cVar1S2S33P016P063P056P059(0) <='1';
          else
          cVar1S2S33P016P063P056P059(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='0' AND E(11)='0' )then
          cVar1S3S33P016P063P056P059(0) <='1';
          else
          cVar1S3S33P016P063P056P059(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='0' AND E(11)='1' )then
          cVar1S4S33P016P063P056P059(0) <='1';
          else
          cVar1S4S33P016P063P056P059(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND D( 3)='1' AND E( 2)='0' )then
          cVar1S5S33P016P063P056P062(0) <='1';
          else
          cVar1S5S33P016P063P056P062(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='1' )then
          cVar1S6S33P016N063P059P014(0) <='1';
          else
          cVar1S6S33P016N063P059P014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='1' )then
          cVar1S7S33P016N063P059P014(0) <='1';
          else
          cVar1S7S33P016N063P059P014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='1' )then
          cVar1S8S33P016N063P059P014(0) <='1';
          else
          cVar1S8S33P016N063P059P014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='0' )then
          cVar1S9S33P016N063P059N014(0) <='1';
          else
          cVar1S9S33P016N063P059N014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='0' )then
          cVar1S10S33P016N063P059N014(0) <='1';
          else
          cVar1S10S33P016N063P059N014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='0' AND A(12)='0' )then
          cVar1S11S33P016N063P059N014(0) <='1';
          else
          cVar1S11S33P016N063P059N014(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='1' AND B(13)='1' )then
          cVar1S12S33P016N063P059P032(0) <='1';
          else
          cVar1S12S33P016N063P059P032(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='1' AND B(13)='1' )then
          cVar1S13S33P016N063P059P032(0) <='1';
          else
          cVar1S13S33P016N063P059P032(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='1' AND B(13)='0' )then
          cVar1S14S33P016N063P059N032(0) <='1';
          else
          cVar1S14S33P016N063P059N032(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND E(11)='1' AND B(13)='0' )then
          cVar1S15S33P016N063P059N032(0) <='1';
          else
          cVar1S15S33P016N063P059N032(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S16S33N016P034P040P021(0) <='1';
          else
          cVar1S16S33N016P034P040P021(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S17S33N016P034P040P021(0) <='1';
          else
          cVar1S17S33N016P034P040P021(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S18S33N016P034P040P021(0) <='1';
          else
          cVar1S18S33N016P034P040P021(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S19S33N016P034P040N021(0) <='1';
          else
          cVar1S19S33N016P034P040N021(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S20S33N016P034P040N021(0) <='1';
          else
          cVar1S20S33N016P034P040N021(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S21S33N016P034N040P044(0) <='1';
          else
          cVar1S21S33N016P034N040P044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S22S33N016P034N040P044(0) <='1';
          else
          cVar1S22S33N016P034N040P044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S23S33N016P034N040P044(0) <='1';
          else
          cVar1S23S33N016P034N040P044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S24S33N016P034N040N044(0) <='1';
          else
          cVar1S24S33N016P034N040N044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S25S33N016P034N040N044(0) <='1';
          else
          cVar1S25S33N016P034N040N044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S26S33N016P034N040N044(0) <='1';
          else
          cVar1S26S33N016P034N040N044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S27S33N016P034N040N044(0) <='1';
          else
          cVar1S27S33N016P034N040N044(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='1' AND A(12)='1' AND D(12)='0' )then
          cVar1S28S33N016P034P014P053(0) <='1';
          else
          cVar1S28S33N016P034P014P053(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='1' AND A(12)='1' AND D(12)='0' )then
          cVar1S29S33N016P034P014P053(0) <='1';
          else
          cVar1S29S33N016P034P014P053(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='1' AND A(12)='1' AND D(12)='0' )then
          cVar1S30S33N016P034P014P053(0) <='1';
          else
          cVar1S30S33N016P034P014P053(0) <='0';
          end if;
        if(A(11)='0' AND B(12)='1' AND A(12)='0' AND A( 1)='1' )then
          cVar1S31S33N016P034N014P017(0) <='1';
          else
          cVar1S31S33N016P034N014P017(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='1' )then
          cVar1S0S34P067P062P008P049(0) <='1';
          else
          cVar1S0S34P067P062P008P049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='1' )then
          cVar1S1S34P067P062P008P049(0) <='1';
          else
          cVar1S1S34P067P062P008P049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='0' )then
          cVar1S2S34P067P062P008N049(0) <='1';
          else
          cVar1S2S34P067P062P008N049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='0' )then
          cVar1S3S34P067P062P008N049(0) <='1';
          else
          cVar1S3S34P067P062P008N049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='0' )then
          cVar1S4S34P067P062P008N049(0) <='1';
          else
          cVar1S4S34P067P062P008N049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='1' AND D(13)='0' )then
          cVar1S5S34P067P062P008N049(0) <='1';
          else
          cVar1S5S34P067P062P008N049(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='0' )then
          cVar1S6S34P067P062N008P035(0) <='1';
          else
          cVar1S6S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='0' )then
          cVar1S7S34P067P062N008P035(0) <='1';
          else
          cVar1S7S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='0' )then
          cVar1S8S34P067P062N008P035(0) <='1';
          else
          cVar1S8S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='0' )then
          cVar1S9S34P067P062N008P035(0) <='1';
          else
          cVar1S9S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='1' )then
          cVar1S10S34P067P062N008P035(0) <='1';
          else
          cVar1S10S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='1' )then
          cVar1S11S34P067P062N008P035(0) <='1';
          else
          cVar1S11S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='1' )then
          cVar1S12S34P067P062N008P035(0) <='1';
          else
          cVar1S12S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='0' AND A(15)='0' AND B( 2)='1' )then
          cVar1S13S34P067P062N008P035(0) <='1';
          else
          cVar1S13S34P067P062N008P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='1' )then
          cVar1S14S34P067P062P055P035(0) <='1';
          else
          cVar1S14S34P067P062P055P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='1' )then
          cVar1S15S34P067P062P055P035(0) <='1';
          else
          cVar1S15S34P067P062P055P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='1' )then
          cVar1S16S34P067P062P055P035(0) <='1';
          else
          cVar1S16S34P067P062P055P035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S17S34P067P062P055N035(0) <='1';
          else
          cVar1S17S34P067P062P055N035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S18S34P067P062P055N035(0) <='1';
          else
          cVar1S18S34P067P062P055N035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='0' AND B( 2)='0' )then
          cVar1S19S34P067P062P055N035(0) <='1';
          else
          cVar1S19S34P067P062P055N035(0) <='0';
          end if;
        if(E( 9)='0' AND E( 2)='1' AND E(12)='1' AND D( 0)='1' )then
          cVar1S20S34P067P062P055P068nsss(0) <='1';
          else
          cVar1S20S34P067P062P055P068nsss(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='0' AND D( 8)='1' AND B( 4)='0' )then
          cVar1S21S34P067P010P069P031(0) <='1';
          else
          cVar1S21S34P067P010P069P031(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='0' AND D( 8)='1' AND B( 4)='0' )then
          cVar1S22S34P067P010P069P031(0) <='1';
          else
          cVar1S22S34P067P010P069P031(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='0' AND D( 8)='1' AND B( 4)='0' )then
          cVar1S23S34P067P010P069P031(0) <='1';
          else
          cVar1S23S34P067P010P069P031(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='0' AND D( 8)='1' AND B( 4)='1' )then
          cVar1S24S34P067P010P069P031(0) <='1';
          else
          cVar1S24S34P067P010P069P031(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='0' AND D( 8)='0' AND D( 4)='1' )then
          cVar1S25S34P067P010N069P052nsss(0) <='1';
          else
          cVar1S25S34P067P010N069P052nsss(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='1' AND A( 2)='1' AND B(11)='0' )then
          cVar1S26S34P067P010P015P036(0) <='1';
          else
          cVar1S26S34P067P010P015P036(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='1' AND A( 2)='1' AND B(11)='1' )then
          cVar1S27S34P067P010P015P036(0) <='1';
          else
          cVar1S27S34P067P010P015P036(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='1' AND A( 2)='0' AND E( 5)='1' )then
          cVar1S28S34P067P010N015P050nsss(0) <='1';
          else
          cVar1S28S34P067P010N015P050nsss(0) <='0';
          end if;
        if(E( 9)='1' AND A(14)='1' AND A( 2)='0' AND E( 5)='0' )then
          cVar1S29S34P067P010N015N050(0) <='1';
          else
          cVar1S29S34P067P010N015N050(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S0S35P058P035P013P066(0) <='1';
          else
          cVar1S0S35P058P035P013P066(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S1S35P058P035P013P066(0) <='1';
          else
          cVar1S1S35P058P035P013P066(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='1' AND E( 1)='0' )then
          cVar1S2S35P058P035P013P066(0) <='1';
          else
          cVar1S2S35P058P035P013P066(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='1' AND E( 1)='1' )then
          cVar1S3S35P058P035P013P066(0) <='1';
          else
          cVar1S3S35P058P035P013P066(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='0' AND A(17)='0' )then
          cVar1S4S35P058P035N013P004(0) <='1';
          else
          cVar1S4S35P058P035N013P004(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='0' AND A(17)='0' )then
          cVar1S5S35P058P035N013P004(0) <='1';
          else
          cVar1S5S35P058P035N013P004(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='0' AND A( 3)='0' AND A(17)='0' )then
          cVar1S6S35P058P035N013P004(0) <='1';
          else
          cVar1S6S35P058P035N013P004(0) <='0';
          end if;
        if(E( 3)='1' AND B( 2)='1' AND D( 2)='1' AND B(12)='0' )then
          cVar1S7S35P058P035P060P034(0) <='1';
          else
          cVar1S7S35P058P035P060P034(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='1' AND B( 4)='0' )then
          cVar1S8S35N058P030P012P031(0) <='1';
          else
          cVar1S8S35N058P030P012P031(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='1' AND B( 4)='0' )then
          cVar1S9S35N058P030P012P031(0) <='1';
          else
          cVar1S9S35N058P030P012P031(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='1' AND B( 4)='0' )then
          cVar1S10S35N058P030P012P031(0) <='1';
          else
          cVar1S10S35N058P030P012P031(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='0' AND A(14)='1' )then
          cVar1S11S35N058P030N012P010(0) <='1';
          else
          cVar1S11S35N058P030N012P010(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='0' AND A(14)='1' )then
          cVar1S12S35N058P030N012P010(0) <='1';
          else
          cVar1S12S35N058P030N012P010(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='1' AND A(13)='0' AND A(14)='0' )then
          cVar1S13S35N058P030N012N010(0) <='1';
          else
          cVar1S13S35N058P030N012N010(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S14S35N058N030P024P006(0) <='1';
          else
          cVar1S14S35N058N030P024P006(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S15S35N058N030P024P006(0) <='1';
          else
          cVar1S15S35N058N030P024P006(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='1' AND A(16)='1' )then
          cVar1S16S35N058N030P024P006(0) <='1';
          else
          cVar1S16S35N058N030P024P006(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='1' AND A(16)='0' )then
          cVar1S17S35N058N030P024N006(0) <='1';
          else
          cVar1S17S35N058N030P024N006(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='1' AND A(16)='0' )then
          cVar1S18S35N058N030P024N006(0) <='1';
          else
          cVar1S18S35N058N030P024N006(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='1' )then
          cVar1S19S35N058N030N024P037(0) <='1';
          else
          cVar1S19S35N058N030N024P037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='1' )then
          cVar1S20S35N058N030N024P037(0) <='1';
          else
          cVar1S20S35N058N030N024P037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='1' )then
          cVar1S21S35N058N030N024P037(0) <='1';
          else
          cVar1S21S35N058N030N024P037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='0' )then
          cVar1S22S35N058N030N024N037(0) <='1';
          else
          cVar1S22S35N058N030N024N037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='0' )then
          cVar1S23S35N058N030N024N037(0) <='1';
          else
          cVar1S23S35N058N030N024N037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='0' )then
          cVar1S24S35N058N030N024N037(0) <='1';
          else
          cVar1S24S35N058N030N024N037(0) <='0';
          end if;
        if(E( 3)='0' AND B(14)='0' AND B(17)='0' AND B( 1)='0' )then
          cVar1S25S35N058N030N024N037(0) <='1';
          else
          cVar1S25S35N058N030N024N037(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='1' AND B( 7)='1' AND E( 9)='0' )then
          cVar1S0S36P037P048P025P067nsss(0) <='1';
          else
          cVar1S0S36P037P048P025P067nsss(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='1' AND B( 7)='0' AND A( 5)='1' )then
          cVar1S1S36P037P048N025P009(0) <='1';
          else
          cVar1S1S36P037P048N025P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='1' AND B( 7)='0' AND A( 5)='1' )then
          cVar1S2S36P037P048N025P009(0) <='1';
          else
          cVar1S2S36P037P048N025P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='1' AND B( 7)='0' AND A( 5)='0' )then
          cVar1S3S36P037P048N025N009(0) <='1';
          else
          cVar1S3S36P037P048N025N009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='1' AND B( 7)='0' AND A( 5)='0' )then
          cVar1S4S36P037P048N025N009(0) <='1';
          else
          cVar1S4S36P037P048N025N009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S5S36P037N048P046P009(0) <='1';
          else
          cVar1S5S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S6S36P037N048P046P009(0) <='1';
          else
          cVar1S6S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S7S36P037N048P046P009(0) <='1';
          else
          cVar1S7S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='1' )then
          cVar1S8S36P037N048P046P009(0) <='1';
          else
          cVar1S8S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='1' )then
          cVar1S9S36P037N048P046P009(0) <='1';
          else
          cVar1S9S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='0' AND A( 5)='1' )then
          cVar1S10S36P037N048P046P009(0) <='1';
          else
          cVar1S10S36P037N048P046P009(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='1' AND D( 6)='1' )then
          cVar1S11S36P037N048P046P044(0) <='1';
          else
          cVar1S11S36P037N048P046P044(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='1' AND D( 6)='1' )then
          cVar1S12S36P037N048P046P044(0) <='1';
          else
          cVar1S12S36P037N048P046P044(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='1' AND D( 6)='1' )then
          cVar1S13S36P037N048P046P044(0) <='1';
          else
          cVar1S13S36P037N048P046P044(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='1' AND D( 6)='1' )then
          cVar1S14S36P037N048P046P044(0) <='1';
          else
          cVar1S14S36P037N048P046P044(0) <='0';
          end if;
        if(B( 1)='0' AND D( 5)='0' AND E( 6)='1' AND D( 6)='0' )then
          cVar1S15S36P037N048P046N044(0) <='1';
          else
          cVar1S15S36P037N048P046N044(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='0' AND B( 2)='1' )then
          cVar1S16S36P037P059P005P035(0) <='1';
          else
          cVar1S16S36P037P059P005P035(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='0' AND B( 2)='1' )then
          cVar1S17S36P037P059P005P035(0) <='1';
          else
          cVar1S17S36P037P059P005P035(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='0' AND B( 2)='0' )then
          cVar1S18S36P037P059P005N035(0) <='1';
          else
          cVar1S18S36P037P059P005N035(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='0' AND B( 2)='0' )then
          cVar1S19S36P037P059P005N035(0) <='1';
          else
          cVar1S19S36P037P059P005N035(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='0' AND B( 2)='0' )then
          cVar1S20S36P037P059P005N035(0) <='1';
          else
          cVar1S20S36P037P059P005N035(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='0' AND A( 7)='1' AND E(10)='0' )then
          cVar1S21S36P037P059P005P063(0) <='1';
          else
          cVar1S21S36P037P059P005P063(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='1' AND A(15)='1' )then
          cVar1S22S36P037P059P008nsss(0) <='1';
          else
          cVar1S22S36P037P059P008nsss(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='1' AND A(15)='0' AND D( 2)='1' )then
          cVar1S23S36P037P059N008P060(0) <='1';
          else
          cVar1S23S36P037P059N008P060(0) <='0';
          end if;
        if(B( 1)='1' AND E(11)='1' AND A(15)='0' AND D( 2)='0' )then
          cVar1S24S36P037P059N008N060(0) <='1';
          else
          cVar1S24S36P037P059N008N060(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S37P048P025P007nsss(0) <='1';
          else
          cVar1S0S37P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='1' )then
          cVar1S1S37P048P025N007P004nsss(0) <='1';
          else
          cVar1S1S37P048P025N007P004nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S2S37P048P025N007N004(0) <='1';
          else
          cVar1S2S37P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S3S37P048P025N007N004(0) <='1';
          else
          cVar1S3S37P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S4S37P048P025N007N004(0) <='1';
          else
          cVar1S4S37P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='0' AND A( 1)='0' )then
          cVar1S5S37P048N025P037P017nsss(0) <='1';
          else
          cVar1S5S37P048N025P037P017nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='0' AND A( 1)='1' )then
          cVar1S6S37P048N025P037P017(0) <='1';
          else
          cVar1S6S37P048N025P037P017(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='0' AND A( 1)='1' )then
          cVar1S7S37P048N025P037P017(0) <='1';
          else
          cVar1S7S37P048N025P037P017(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='0' AND A( 1)='1' )then
          cVar1S8S37P048N025P037P017(0) <='1';
          else
          cVar1S8S37P048N025P037P017(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='1' AND A(16)='1' )then
          cVar1S9S37P048N025P037P006nsss(0) <='1';
          else
          cVar1S9S37P048N025P037P006nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 1)='1' AND A(16)='0' )then
          cVar1S10S37P048N025P037N006(0) <='1';
          else
          cVar1S10S37P048N025P037N006(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='1' )then
          cVar1S11S37N048P044P004nsss(0) <='1';
          else
          cVar1S11S37N048P044P004nsss(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='1' )then
          cVar1S12S37N048P044N004P005(0) <='1';
          else
          cVar1S12S37N048P044N004P005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='1' )then
          cVar1S13S37N048P044N004P005(0) <='1';
          else
          cVar1S13S37N048P044N004P005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S14S37N048P044N004N005(0) <='1';
          else
          cVar1S14S37N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S15S37N048P044N004N005(0) <='1';
          else
          cVar1S15S37N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S16S37N048P044N004N005(0) <='1';
          else
          cVar1S16S37N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S17S37N048P044N004N005(0) <='1';
          else
          cVar1S17S37N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S18S37N048N044P046P025(0) <='1';
          else
          cVar1S18S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S19S37N048N044P046P025(0) <='1';
          else
          cVar1S19S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='0' )then
          cVar1S20S37N048N044P046P025(0) <='1';
          else
          cVar1S20S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='1' )then
          cVar1S21S37N048N044P046P025(0) <='1';
          else
          cVar1S21S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='1' )then
          cVar1S22S37N048N044P046P025(0) <='1';
          else
          cVar1S22S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND B( 7)='1' )then
          cVar1S23S37N048N044P046P025(0) <='1';
          else
          cVar1S23S37N048N044P046P025(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S24S37N048N044P046P027(0) <='1';
          else
          cVar1S24S37N048N044P046P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S38P048P025P007nsss(0) <='1';
          else
          cVar1S0S38P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='1' )then
          cVar1S1S38P048P025N007P004nsss(0) <='1';
          else
          cVar1S1S38P048P025N007P004nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S2S38P048P025N007N004(0) <='1';
          else
          cVar1S2S38P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S3S38P048P025N007N004(0) <='1';
          else
          cVar1S3S38P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S4S38P048P025N007N004(0) <='1';
          else
          cVar1S4S38P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='1' )then
          cVar1S5S38P048N025P052P027(0) <='1';
          else
          cVar1S5S38P048N025P052P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='1' )then
          cVar1S6S38P048N025P052P027(0) <='1';
          else
          cVar1S6S38P048N025P052P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='1' )then
          cVar1S7S38P048N025P052P027(0) <='1';
          else
          cVar1S7S38P048N025P052P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='0' )then
          cVar1S8S38P048N025P052N027(0) <='1';
          else
          cVar1S8S38P048N025P052N027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='0' )then
          cVar1S9S38P048N025P052N027(0) <='1';
          else
          cVar1S9S38P048N025P052N027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND B( 6)='0' )then
          cVar1S10S38P048N025P052N027(0) <='1';
          else
          cVar1S10S38P048N025P052N027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='1' AND E( 6)='1' )then
          cVar1S11S38P048N025P052P046nsss(0) <='1';
          else
          cVar1S11S38P048N025P052P046nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='1' AND E( 6)='0' )then
          cVar1S12S38P048N025P052N046(0) <='1';
          else
          cVar1S12S38P048N025P052N046(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='1' )then
          cVar1S13S38N048P025P046P018(0) <='1';
          else
          cVar1S13S38N048P025P046P018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='1' )then
          cVar1S14S38N048P025P046P018(0) <='1';
          else
          cVar1S14S38N048P025P046P018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='1' )then
          cVar1S15S38N048P025P046P018(0) <='1';
          else
          cVar1S15S38N048P025P046P018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='0' )then
          cVar1S16S38N048P025P046N018(0) <='1';
          else
          cVar1S16S38N048P025P046N018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='0' )then
          cVar1S17S38N048P025P046N018(0) <='1';
          else
          cVar1S17S38N048P025P046N018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='0' )then
          cVar1S18S38N048P025P046N018(0) <='1';
          else
          cVar1S18S38N048P025P046N018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='0' AND A(10)='0' )then
          cVar1S19S38N048P025P046N018(0) <='1';
          else
          cVar1S19S38N048P025P046N018(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S20S38N048P025P046P027(0) <='1';
          else
          cVar1S20S38N048P025P046P027(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S21S38N048P025P046P027(0) <='1';
          else
          cVar1S21S38N048P025P046P027(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S22S38N048P025P046P027(0) <='1';
          else
          cVar1S22S38N048P025P046P027(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='1' AND A( 6)='1' AND A( 5)='0' )then
          cVar1S23S38N048P025P007P009(0) <='1';
          else
          cVar1S23S38N048P025P007P009(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='1' AND A( 6)='1' AND A( 5)='0' )then
          cVar1S24S38N048P025P007P009(0) <='1';
          else
          cVar1S24S38N048P025P007P009(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='1' AND A( 6)='1' AND A( 5)='0' )then
          cVar1S25S38N048P025P007P009(0) <='1';
          else
          cVar1S25S38N048P025P007P009(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='1' AND A( 6)='0' AND D( 6)='1' )then
          cVar1S26S38N048P025N007P044(0) <='1';
          else
          cVar1S26S38N048P025N007P044(0) <='0';
          end if;
        if(D( 5)='0' AND B( 7)='1' AND A( 6)='0' AND D( 6)='0' )then
          cVar1S27S38N048P025N007N044(0) <='1';
          else
          cVar1S27S38N048P025N007N044(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S39P048P025P007nsss(0) <='1';
          else
          cVar1S0S39P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='1' )then
          cVar1S1S39P048P025N007P004nsss(0) <='1';
          else
          cVar1S1S39P048P025N007P004nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S2S39P048P025N007N004(0) <='1';
          else
          cVar1S2S39P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S3S39P048P025N007N004(0) <='1';
          else
          cVar1S3S39P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S4S39P048P025N007N004(0) <='1';
          else
          cVar1S4S39P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 6)='1' )then
          cVar1S5S39P048N025P027P007nsss(0) <='1';
          else
          cVar1S5S39P048N025P027P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 6)='0' )then
          cVar1S6S39P048N025P027N007(0) <='1';
          else
          cVar1S6S39P048N025P027N007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 6)='0' )then
          cVar1S7S39P048N025P027N007(0) <='1';
          else
          cVar1S7S39P048N025P027N007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='1' AND A( 6)='0' )then
          cVar1S8S39P048N025P027N007(0) <='1';
          else
          cVar1S8S39P048N025P027N007(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 3)='1' )then
          cVar1S9S39P048N025N027P058nsss(0) <='1';
          else
          cVar1S9S39P048N025N027P058nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 3)='0' )then
          cVar1S10S39P048N025N027N058(0) <='1';
          else
          cVar1S10S39P048N025N027N058(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 3)='0' )then
          cVar1S11S39P048N025N027N058(0) <='1';
          else
          cVar1S11S39P048N025N027N058(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND B( 6)='0' AND E( 3)='0' )then
          cVar1S12S39P048N025N027N058(0) <='1';
          else
          cVar1S12S39P048N025N027N058(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='1' )then
          cVar1S13S39N048P044P004nsss(0) <='1';
          else
          cVar1S13S39N048P044P004nsss(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='1' )then
          cVar1S14S39N048P044N004P005(0) <='1';
          else
          cVar1S14S39N048P044N004P005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='1' )then
          cVar1S15S39N048P044N004P005(0) <='1';
          else
          cVar1S15S39N048P044N004P005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S16S39N048P044N004N005(0) <='1';
          else
          cVar1S16S39N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S17S39N048P044N004N005(0) <='1';
          else
          cVar1S17S39N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S18S39N048P044N004N005(0) <='1';
          else
          cVar1S18S39N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='1' AND A(17)='0' AND A( 7)='0' )then
          cVar1S19S39N048P044N004N005(0) <='1';
          else
          cVar1S19S39N048P044N004N005(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='1' )then
          cVar1S20S39N048N044P046P052(0) <='1';
          else
          cVar1S20S39N048N044P046P052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='1' )then
          cVar1S21S39N048N044P046P052(0) <='1';
          else
          cVar1S21S39N048N044P046P052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='1' )then
          cVar1S22S39N048N044P046P052(0) <='1';
          else
          cVar1S22S39N048N044P046P052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='1' )then
          cVar1S23S39N048N044P046P052(0) <='1';
          else
          cVar1S23S39N048N044P046P052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='0' )then
          cVar1S24S39N048N044P046N052(0) <='1';
          else
          cVar1S24S39N048N044P046N052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='0' )then
          cVar1S25S39N048N044P046N052(0) <='1';
          else
          cVar1S25S39N048N044P046N052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='0' AND D( 4)='0' )then
          cVar1S26S39N048N044P046N052(0) <='1';
          else
          cVar1S26S39N048N044P046N052(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S27S39N048N044P046P027(0) <='1';
          else
          cVar1S27S39N048N044P046P027(0) <='0';
          end if;
        if(D( 5)='0' AND D( 6)='0' AND E( 6)='1' AND B( 6)='0' )then
          cVar1S28S39N048N044P046P027(0) <='1';
          else
          cVar1S28S39N048N044P046P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S0S40P018P048P025nsss(0) <='1';
          else
          cVar1S0S40P018P048P025nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S1S40P018P048N025P027(0) <='1';
          else
          cVar1S1S40P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S2S40P018P048N025P027(0) <='1';
          else
          cVar1S2S40P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S3S40P018P048N025P027(0) <='1';
          else
          cVar1S3S40P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S4S40P018P048N025N027(0) <='1';
          else
          cVar1S4S40P018P048N025N027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S5S40P018P048N025N027(0) <='1';
          else
          cVar1S5S40P018P048N025N027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='1' )then
          cVar1S6S40P018N048P010P032(0) <='1';
          else
          cVar1S6S40P018N048P010P032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='1' )then
          cVar1S7S40P018N048P010P032(0) <='1';
          else
          cVar1S7S40P018N048P010P032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='1' )then
          cVar1S8S40P018N048P010P032(0) <='1';
          else
          cVar1S8S40P018N048P010P032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='1' )then
          cVar1S9S40P018N048P010P032(0) <='1';
          else
          cVar1S9S40P018N048P010P032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='0' )then
          cVar1S10S40P018N048P010N032(0) <='1';
          else
          cVar1S10S40P018N048P010N032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='0' )then
          cVar1S11S40P018N048P010N032(0) <='1';
          else
          cVar1S11S40P018N048P010N032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='0' )then
          cVar1S12S40P018N048P010N032(0) <='1';
          else
          cVar1S12S40P018N048P010N032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='0' AND B(13)='0' )then
          cVar1S13S40P018N048P010N032(0) <='1';
          else
          cVar1S13S40P018N048P010N032(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='1' )then
          cVar1S14S40P018N048P010P028(0) <='1';
          else
          cVar1S14S40P018N048P010P028(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='1' )then
          cVar1S15S40P018N048P010P028(0) <='1';
          else
          cVar1S15S40P018N048P010P028(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='1' )then
          cVar1S16S40P018N048P010P028(0) <='1';
          else
          cVar1S16S40P018N048P010P028(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='0' )then
          cVar1S17S40P018N048P010N028(0) <='1';
          else
          cVar1S17S40P018N048P010N028(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='0' )then
          cVar1S18S40P018N048P010N028(0) <='1';
          else
          cVar1S18S40P018N048P010N028(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND A(14)='1' AND B(15)='0' )then
          cVar1S19S40P018N048P010N028(0) <='1';
          else
          cVar1S19S40P018N048P010N028(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='1' AND D( 0)='0' )then
          cVar1S20S40P018P069P009P068(0) <='1';
          else
          cVar1S20S40P018P069P009P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='1' AND D( 0)='1' )then
          cVar1S21S40P018P069P009P068(0) <='1';
          else
          cVar1S21S40P018P069P009P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='1' AND D( 0)='1' )then
          cVar1S22S40P018P069P009P068(0) <='1';
          else
          cVar1S22S40P018P069P009P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='1' )then
          cVar1S23S40P018P069N009P003(0) <='1';
          else
          cVar1S23S40P018P069N009P003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='1' )then
          cVar1S24S40P018P069N009P003(0) <='1';
          else
          cVar1S24S40P018P069N009P003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='0' )then
          cVar1S25S40P018P069N009N003(0) <='1';
          else
          cVar1S25S40P018P069N009N003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='0' )then
          cVar1S26S40P018P069N009N003(0) <='1';
          else
          cVar1S26S40P018P069N009N003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='0' )then
          cVar1S27S40P018P069N009N003(0) <='1';
          else
          cVar1S27S40P018P069N009N003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND A( 5)='0' AND A( 8)='0' )then
          cVar1S28S40P018P069N009N003(0) <='1';
          else
          cVar1S28S40P018P069N009N003(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND D( 4)='1' AND B( 5)='0' )then
          cVar1S29S40P018P069P052P029nsss(0) <='1';
          else
          cVar1S29S40P018P069P052P029nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S41P048P025P007nsss(0) <='1';
          else
          cVar1S0S41P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='1' )then
          cVar1S1S41P048P025N007P004nsss(0) <='1';
          else
          cVar1S1S41P048P025N007P004nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S2S41P048P025N007N004(0) <='1';
          else
          cVar1S2S41P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S3S41P048P025N007N004(0) <='1';
          else
          cVar1S3S41P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S4S41P048P025N007N004(0) <='1';
          else
          cVar1S4S41P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND D( 9)='0' )then
          cVar1S5S41P048N025P052P065(0) <='1';
          else
          cVar1S5S41P048N025P052P065(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND D( 9)='0' )then
          cVar1S6S41P048N025P052P065(0) <='1';
          else
          cVar1S6S41P048N025P052P065(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND D( 9)='0' )then
          cVar1S7S41P048N025P052P065(0) <='1';
          else
          cVar1S7S41P048N025P052P065(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='0' AND D( 9)='1' )then
          cVar1S8S41P048N025P052P065(0) <='1';
          else
          cVar1S8S41P048N025P052P065(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='1' AND A( 2)='1' )then
          cVar1S9S41P048N025P052P015nsss(0) <='1';
          else
          cVar1S9S41P048N025P052P015nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='1' AND A( 2)='0' )then
          cVar1S10S41P048N025P052N015(0) <='1';
          else
          cVar1S10S41P048N025P052N015(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND D( 4)='1' AND A( 2)='0' )then
          cVar1S11S41P048N025P052N015(0) <='1';
          else
          cVar1S11S41P048N025P052N015(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='0' )then
          cVar1S12S41N048P018P059P045(0) <='1';
          else
          cVar1S12S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='0' )then
          cVar1S13S41N048P018P059P045(0) <='1';
          else
          cVar1S13S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='0' )then
          cVar1S14S41N048P018P059P045(0) <='1';
          else
          cVar1S14S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='1' )then
          cVar1S15S41N048P018P059P045(0) <='1';
          else
          cVar1S15S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='1' )then
          cVar1S16S41N048P018P059P045(0) <='1';
          else
          cVar1S16S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='0' AND D(14)='1' )then
          cVar1S17S41N048P018P059P045(0) <='1';
          else
          cVar1S17S41N048P018P059P045(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='1' AND E( 5)='1' )then
          cVar1S18S41N048P018P059P050nsss(0) <='1';
          else
          cVar1S18S41N048P018P059P050nsss(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='1' AND E( 5)='0' )then
          cVar1S19S41N048P018P059N050(0) <='1';
          else
          cVar1S19S41N048P018P059N050(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='1' AND E(11)='1' AND E( 5)='0' )then
          cVar1S20S41N048P018P059N050(0) <='1';
          else
          cVar1S20S41N048P018P059N050(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='1' AND B(15)='0' )then
          cVar1S21S41N048N018P032P028(0) <='1';
          else
          cVar1S21S41N048N018P032P028(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='1' AND B(15)='0' )then
          cVar1S22S41N048N018P032P028(0) <='1';
          else
          cVar1S22S41N048N018P032P028(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='1' AND B(15)='0' )then
          cVar1S23S41N048N018P032P028(0) <='1';
          else
          cVar1S23S41N048N018P032P028(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='1' )then
          cVar1S24S41N048N018N032P056(0) <='1';
          else
          cVar1S24S41N048N018N032P056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='1' )then
          cVar1S25S41N048N018N032P056(0) <='1';
          else
          cVar1S25S41N048N018N032P056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='1' )then
          cVar1S26S41N048N018N032P056(0) <='1';
          else
          cVar1S26S41N048N018N032P056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='1' )then
          cVar1S27S41N048N018N032P056(0) <='1';
          else
          cVar1S27S41N048N018N032P056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='0' )then
          cVar1S28S41N048N018N032N056(0) <='1';
          else
          cVar1S28S41N048N018N032N056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='0' )then
          cVar1S29S41N048N018N032N056(0) <='1';
          else
          cVar1S29S41N048N018N032N056(0) <='0';
          end if;
        if(D( 5)='0' AND A(10)='0' AND B(13)='0' AND D( 3)='0' )then
          cVar1S30S41N048N018N032N056(0) <='1';
          else
          cVar1S30S41N048N018N032N056(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='1' )then
          cVar1S0S42P018P048P025nsss(0) <='1';
          else
          cVar1S0S42P018P048P025nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S1S42P018P048N025P027(0) <='1';
          else
          cVar1S1S42P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S2S42P018P048N025P027(0) <='1';
          else
          cVar1S2S42P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='1' )then
          cVar1S3S42P018P048N025P027(0) <='1';
          else
          cVar1S3S42P018P048N025P027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S4S42P018P048N025N027(0) <='1';
          else
          cVar1S4S42P018P048N025N027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S5S42P018P048N025N027(0) <='1';
          else
          cVar1S5S42P018P048N025N027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='1' AND B( 7)='0' AND B( 6)='0' )then
          cVar1S6S42P018P048N025N027(0) <='1';
          else
          cVar1S6S42P018P048N025N027(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='1' AND A(18)='1' )then
          cVar1S7S42P018N048P038P002nsss(0) <='1';
          else
          cVar1S7S42P018N048P038P002nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='1' AND A(18)='0' )then
          cVar1S8S42P018N048P038N002(0) <='1';
          else
          cVar1S8S42P018N048P038N002(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='1' AND A(18)='0' )then
          cVar1S9S42P018N048P038N002(0) <='1';
          else
          cVar1S9S42P018N048P038N002(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='0' AND A(19)='0' )then
          cVar1S10S42P018N048N038P000(0) <='1';
          else
          cVar1S10S42P018N048N038P000(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='0' AND A(19)='0' )then
          cVar1S11S42P018N048N038P000(0) <='1';
          else
          cVar1S11S42P018N048N038P000(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='0' AND A(19)='0' )then
          cVar1S12S42P018N048N038P000(0) <='1';
          else
          cVar1S12S42P018N048N038P000(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='0' AND A(19)='0' )then
          cVar1S13S42P018N048N038P000(0) <='1';
          else
          cVar1S13S42P018N048N038P000(0) <='0';
          end if;
        if(A(10)='0' AND D( 5)='0' AND B(10)='0' AND A(19)='1' )then
          cVar1S14S42P018N048N038P000(0) <='1';
          else
          cVar1S14S42P018N048N038P000(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='1' AND A( 4)='0' AND A(15)='0' )then
          cVar1S15S42P018P048P011P008(0) <='1';
          else
          cVar1S15S42P018P048P011P008(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='1' AND A( 4)='0' AND A(15)='0' )then
          cVar1S16S42P018P048P011P008(0) <='1';
          else
          cVar1S16S42P018P048P011P008(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='1' AND A( 4)='0' AND A(15)='0' )then
          cVar1S17S42P018P048P011P008(0) <='1';
          else
          cVar1S17S42P018P048P011P008(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='1' AND A( 4)='0' AND A(15)='1' )then
          cVar1S18S42P018P048P011P008(0) <='1';
          else
          cVar1S18S42P018P048P011P008(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='1' AND A( 4)='1' AND A( 3)='0' )then
          cVar1S19S42P018P048P011P013(0) <='1';
          else
          cVar1S19S42P018P048P011P013(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='1' AND B( 8)='1' )then
          cVar1S20S42P018N048P044P023nsss(0) <='1';
          else
          cVar1S20S42P018N048P044P023nsss(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S21S42P018N048P044N023(0) <='1';
          else
          cVar1S21S42P018N048P044N023(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='1' AND B( 8)='0' )then
          cVar1S22S42P018N048P044N023(0) <='1';
          else
          cVar1S22S42P018N048P044N023(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='0' AND A(17)='0' )then
          cVar1S23S42P018N048N044P004(0) <='1';
          else
          cVar1S23S42P018N048N044P004(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='0' AND A(17)='0' )then
          cVar1S24S42P018N048N044P004(0) <='1';
          else
          cVar1S24S42P018N048N044P004(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='0' AND A(17)='1' )then
          cVar1S25S42P018N048N044P004(0) <='1';
          else
          cVar1S25S42P018N048N044P004(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='0' AND A(17)='1' )then
          cVar1S26S42P018N048N044P004(0) <='1';
          else
          cVar1S26S42P018N048N044P004(0) <='0';
          end if;
        if(A(10)='1' AND D( 5)='0' AND D( 6)='0' AND A(17)='1' )then
          cVar1S27S42P018N048N044P004(0) <='1';
          else
          cVar1S27S42P018N048N044P004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S0S43P048P025P007nsss(0) <='1';
          else
          cVar1S0S43P048P025P007nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='1' )then
          cVar1S1S43P048P025N007P004nsss(0) <='1';
          else
          cVar1S1S43P048P025N007P004nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S2S43P048P025N007N004(0) <='1';
          else
          cVar1S2S43P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S3S43P048P025N007N004(0) <='1';
          else
          cVar1S3S43P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='1' AND A( 6)='0' AND A(17)='0' )then
          cVar1S4S43P048P025N007N004(0) <='1';
          else
          cVar1S4S43P048P025N007N004(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='1' AND E( 3)='1' )then
          cVar1S5S43P048N025P062P058nsss(0) <='1';
          else
          cVar1S5S43P048N025P062P058nsss(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='1' AND E( 3)='0' )then
          cVar1S6S43P048N025P062N058(0) <='1';
          else
          cVar1S6S43P048N025P062N058(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S7S43P048N025N062P027(0) <='1';
          else
          cVar1S7S43P048N025N062P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S8S43P048N025N062P027(0) <='1';
          else
          cVar1S8S43P048N025N062P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S9S43P048N025N062P027(0) <='1';
          else
          cVar1S9S43P048N025N062P027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S10S43P048N025N062N027(0) <='1';
          else
          cVar1S10S43P048N025N062N027(0) <='0';
          end if;
        if(D( 5)='1' AND B( 7)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S11S43P048N025N062N027(0) <='1';
          else
          cVar1S11S43P048N025N062N027(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='1' AND E(15)='1' AND A(13)='0' )then
          cVar1S12S43N048P022P043P012(0) <='1';
          else
          cVar1S12S43N048P022P043P012(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar1S13S43N048P022N043P004(0) <='1';
          else
          cVar1S13S43N048P022N043P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='1' AND E(15)='0' AND A(17)='0' )then
          cVar1S14S43N048P022N043N004(0) <='1';
          else
          cVar1S14S43N048P022N043N004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='1' AND B( 9)='1' )then
          cVar1S15S43N048N022P038P021(0) <='1';
          else
          cVar1S15S43N048N022P038P021(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='1' AND B( 9)='1' )then
          cVar1S16S43N048N022P038P021(0) <='1';
          else
          cVar1S16S43N048N022P038P021(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='1' AND B( 9)='0' )then
          cVar1S17S43N048N022P038N021(0) <='1';
          else
          cVar1S17S43N048N022P038N021(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='1' AND B( 9)='0' )then
          cVar1S18S43N048N022P038N021(0) <='1';
          else
          cVar1S18S43N048N022P038N021(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='0' )then
          cVar1S19S43N048N022N038P004(0) <='1';
          else
          cVar1S19S43N048N022N038P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='0' )then
          cVar1S20S43N048N022N038P004(0) <='1';
          else
          cVar1S20S43N048N022N038P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='0' )then
          cVar1S21S43N048N022N038P004(0) <='1';
          else
          cVar1S21S43N048N022N038P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='1' )then
          cVar1S22S43N048N022N038P004(0) <='1';
          else
          cVar1S22S43N048N022N038P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='1' )then
          cVar1S23S43N048N022N038P004(0) <='1';
          else
          cVar1S23S43N048N022N038P004(0) <='0';
          end if;
        if(D( 5)='0' AND B(18)='0' AND B(10)='0' AND A(17)='1' )then
          cVar1S24S43N048N022N038P004(0) <='1';
          else
          cVar1S24S43N048N022N038P004(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND B( 1)='0' AND A(14)='0' )then
          cVar1S0S44P022P043P037P010nsss(0) <='1';
          else
          cVar1S0S44P022P043P037P010nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND B( 1)='1' AND A(17)='1' )then
          cVar1S1S44P022P043P037P004nsss(0) <='1';
          else
          cVar1S1S44P022P043P037P004nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar1S2S44P022N043P004nsss(0) <='1';
          else
          cVar1S2S44P022N043P004nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND E(14)='0' )then
          cVar1S3S44P022N043N004P047(0) <='1';
          else
          cVar1S3S44P022N043N004P047(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='0' )then
          cVar1S4S44N022P004P043P045(0) <='1';
          else
          cVar1S4S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='0' )then
          cVar1S5S44N022P004P043P045(0) <='1';
          else
          cVar1S5S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='0' )then
          cVar1S6S44N022P004P043P045(0) <='1';
          else
          cVar1S6S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='1' )then
          cVar1S7S44N022P004P043P045(0) <='1';
          else
          cVar1S7S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='1' )then
          cVar1S8S44N022P004P043P045(0) <='1';
          else
          cVar1S8S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='1' )then
          cVar1S9S44N022P004P043P045(0) <='1';
          else
          cVar1S9S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='0' AND D(14)='1' )then
          cVar1S10S44N022P004P043P045(0) <='1';
          else
          cVar1S10S44N022P004P043P045(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='1' AND B( 8)='1' )then
          cVar1S11S44N022P004P043P023(0) <='1';
          else
          cVar1S11S44N022P004P043P023(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='1' AND B( 8)='1' )then
          cVar1S12S44N022P004P043P023(0) <='1';
          else
          cVar1S12S44N022P004P043P023(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='1' AND B( 8)='0' )then
          cVar1S13S44N022P004P043N023(0) <='1';
          else
          cVar1S13S44N022P004P043N023(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='1' AND B( 8)='0' )then
          cVar1S14S44N022P004P043N023(0) <='1';
          else
          cVar1S14S44N022P004P043N023(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='0' AND E(15)='1' AND B( 8)='0' )then
          cVar1S15S44N022P004P043N023(0) <='1';
          else
          cVar1S15S44N022P004P043N023(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='1' )then
          cVar1S16S44N022P004P040nsss(0) <='1';
          else
          cVar1S16S44N022P004P040nsss(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='0' AND A( 1)='1' )then
          cVar1S17S44N022P004N040P017(0) <='1';
          else
          cVar1S17S44N022P004N040P017(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='0' AND A( 1)='1' )then
          cVar1S18S44N022P004N040P017(0) <='1';
          else
          cVar1S18S44N022P004N040P017(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='0' AND A( 1)='0' )then
          cVar1S19S44N022P004N040N017(0) <='1';
          else
          cVar1S19S44N022P004N040N017(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='0' AND A( 1)='0' )then
          cVar1S20S44N022P004N040N017(0) <='1';
          else
          cVar1S20S44N022P004N040N017(0) <='0';
          end if;
        if(B(18)='0' AND A(17)='1' AND D( 7)='0' AND A( 1)='0' )then
          cVar1S21S44N022P004N040N017(0) <='1';
          else
          cVar1S21S44N022P004N040N017(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='1' )then
          cVar1S0S45P022P043P019nsss(0) <='1';
          else
          cVar1S0S45P022P043P019nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='0' AND A(13)='0' )then
          cVar1S1S45P022P043N019P012(0) <='1';
          else
          cVar1S1S45P022P043N019P012(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='1' AND E( 7)='1' )then
          cVar1S2S45P022N043P004P042nsss(0) <='1';
          else
          cVar1S2S45P022N043P004P042nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar1S3S45P022N043N004P007nsss(0) <='1';
          else
          cVar1S3S45P022N043N004P007nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND A( 6)='0' )then
          cVar1S4S45P022N043N004N007(0) <='1';
          else
          cVar1S4S45P022N043N004N007(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND A( 6)='0' )then
          cVar1S5S45P022N043N004N007(0) <='1';
          else
          cVar1S5S45P022N043N004N007(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND A( 6)='0' )then
          cVar1S6S45P022N043N004N007(0) <='1';
          else
          cVar1S6S45P022N043N004N007(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='1' )then
          cVar1S7S45N022P047P006nsss(0) <='1';
          else
          cVar1S7S45N022P047P006nsss(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='1' )then
          cVar1S8S45N022P047N006P008(0) <='1';
          else
          cVar1S8S45N022P047N006P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='1' )then
          cVar1S9S45N022P047N006P008(0) <='1';
          else
          cVar1S9S45N022P047N006P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='1' )then
          cVar1S10S45N022P047N006P008(0) <='1';
          else
          cVar1S10S45N022P047N006P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='0' )then
          cVar1S11S45N022P047N006N008(0) <='1';
          else
          cVar1S11S45N022P047N006N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='0' )then
          cVar1S12S45N022P047N006N008(0) <='1';
          else
          cVar1S12S45N022P047N006N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='1' AND A(16)='0' AND A(15)='0' )then
          cVar1S13S45N022P047N006N008(0) <='1';
          else
          cVar1S13S45N022P047N006N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S14S45N022N047P051P008(0) <='1';
          else
          cVar1S14S45N022N047P051P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S15S45N022N047P051P008(0) <='1';
          else
          cVar1S15S45N022N047P051P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='1' )then
          cVar1S16S45N022N047P051P008(0) <='1';
          else
          cVar1S16S45N022N047P051P008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S17S45N022N047P051N008(0) <='1';
          else
          cVar1S17S45N022N047P051N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S18S45N022N047P051N008(0) <='1';
          else
          cVar1S18S45N022N047P051N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='1' AND A(15)='0' )then
          cVar1S19S45N022N047P051N008(0) <='1';
          else
          cVar1S19S45N022N047P051N008(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='0' AND D(13)='0' )then
          cVar1S20S45N022N047N051P049(0) <='1';
          else
          cVar1S20S45N022N047N051P049(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='0' AND D(13)='0' )then
          cVar1S21S45N022N047N051P049(0) <='1';
          else
          cVar1S21S45N022N047N051P049(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='0' AND D(13)='0' )then
          cVar1S22S45N022N047N051P049(0) <='1';
          else
          cVar1S22S45N022N047N051P049(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='0' AND D(13)='1' )then
          cVar1S23S45N022N047N051P049(0) <='1';
          else
          cVar1S23S45N022N047N051P049(0) <='0';
          end if;
        if(B(18)='0' AND E(14)='0' AND E(13)='0' AND D(13)='1' )then
          cVar1S24S45N022N047N051P049(0) <='1';
          else
          cVar1S24S45N022N047N051P049(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='1' )then
          cVar1S0S46P022P043P019nsss(0) <='1';
          else
          cVar1S0S46P022P043P019nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='0' AND B( 1)='0' )then
          cVar1S1S46P022P043N019P037nsss(0) <='1';
          else
          cVar1S1S46P022P043N019P037nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar1S2S46P022N043P004nsss(0) <='1';
          else
          cVar1S2S46P022N043P004nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND E(14)='0' )then
          cVar1S3S46P022N043N004P047(0) <='1';
          else
          cVar1S3S46P022N043N004P047(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND E(14)='0' )then
          cVar1S4S46P022N043N004P047(0) <='1';
          else
          cVar1S4S46P022N043N004P047(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='1' AND E( 5)='0' )then
          cVar1S5S46N022P048P025P050(0) <='1';
          else
          cVar1S5S46N022P048P025P050(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND E(15)='0' )then
          cVar1S6S46N022P048N025P043(0) <='1';
          else
          cVar1S6S46N022P048N025P043(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND E(15)='0' )then
          cVar1S7S46N022P048N025P043(0) <='1';
          else
          cVar1S7S46N022P048N025P043(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='1' AND B( 7)='0' AND E(15)='0' )then
          cVar1S8S46N022P048N025P043(0) <='1';
          else
          cVar1S8S46N022P048N025P043(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='1' AND D( 9)='0' )then
          cVar1S9S46N022N048P037P065(0) <='1';
          else
          cVar1S9S46N022N048P037P065(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='1' AND D( 9)='0' )then
          cVar1S10S46N022N048P037P065(0) <='1';
          else
          cVar1S10S46N022N048P037P065(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='1' AND D( 9)='0' )then
          cVar1S11S46N022N048P037P065(0) <='1';
          else
          cVar1S11S46N022N048P037P065(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='1' AND D( 9)='1' )then
          cVar1S12S46N022N048P037P065(0) <='1';
          else
          cVar1S12S46N022N048P037P065(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='1' AND D( 9)='1' )then
          cVar1S13S46N022N048P037P065(0) <='1';
          else
          cVar1S13S46N022N048P037P065(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='1' )then
          cVar1S14S46N022N048N037P023(0) <='1';
          else
          cVar1S14S46N022N048N037P023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='1' )then
          cVar1S15S46N022N048N037P023(0) <='1';
          else
          cVar1S15S46N022N048N037P023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='1' )then
          cVar1S16S46N022N048N037P023(0) <='1';
          else
          cVar1S16S46N022N048N037P023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='0' )then
          cVar1S17S46N022N048N037N023(0) <='1';
          else
          cVar1S17S46N022N048N037N023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='0' )then
          cVar1S18S46N022N048N037N023(0) <='1';
          else
          cVar1S18S46N022N048N037N023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='0' )then
          cVar1S19S46N022N048N037N023(0) <='1';
          else
          cVar1S19S46N022N048N037N023(0) <='0';
          end if;
        if(B(18)='0' AND D( 5)='0' AND B( 1)='0' AND B( 8)='0' )then
          cVar1S20S46N022N048N037N023(0) <='1';
          else
          cVar1S20S46N022N048N037N023(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='1' )then
          cVar1S0S47P022P043P019nsss(0) <='1';
          else
          cVar1S0S47P022P043P019nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='0' AND A( 3)='0' )then
          cVar1S1S47P022P043N019P013(0) <='1';
          else
          cVar1S1S47P022P043N019P013(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='0' AND A( 3)='0' )then
          cVar1S2S47P022P043N019P013(0) <='1';
          else
          cVar1S2S47P022P043N019P013(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' AND A( 0)='0' AND A( 3)='0' )then
          cVar1S3S47P022P043N019P013(0) <='1';
          else
          cVar1S3S47P022P043N019P013(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='1' AND E( 7)='1' )then
          cVar1S4S47P022N043P004P042nsss(0) <='1';
          else
          cVar1S4S47P022N043P004P042nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND E(14)='0' )then
          cVar1S5S47P022N043N004P047(0) <='1';
          else
          cVar1S5S47P022N043N004P047(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND A(17)='0' AND E(14)='0' )then
          cVar1S6S47P022N043N004P047(0) <='1';
          else
          cVar1S6S47P022N043N004P047(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S7S47N022P023P005P068(0) <='1';
          else
          cVar1S7S47N022P023P005P068(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S8S47N022P023P005P068(0) <='1';
          else
          cVar1S8S47N022P023P005P068(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='1' AND A( 7)='0' AND B(12)='0' )then
          cVar1S9S47N022P023N005P034(0) <='1';
          else
          cVar1S9S47N022P023N005P034(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='1' AND A( 7)='0' AND B(12)='0' )then
          cVar1S10S47N022P023N005P034(0) <='1';
          else
          cVar1S10S47N022P023N005P034(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='1' AND A( 7)='0' AND B(12)='0' )then
          cVar1S11S47N022P023N005P034(0) <='1';
          else
          cVar1S11S47N022P023N005P034(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='1' )then
          cVar1S12S47N022N023P043P048(0) <='1';
          else
          cVar1S12S47N022N023P043P048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='1' )then
          cVar1S13S47N022N023P043P048(0) <='1';
          else
          cVar1S13S47N022N023P043P048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='1' )then
          cVar1S14S47N022N023P043P048(0) <='1';
          else
          cVar1S14S47N022N023P043P048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='0' )then
          cVar1S15S47N022N023P043N048(0) <='1';
          else
          cVar1S15S47N022N023P043N048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='0' )then
          cVar1S16S47N022N023P043N048(0) <='1';
          else
          cVar1S16S47N022N023P043N048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='0' )then
          cVar1S17S47N022N023P043N048(0) <='1';
          else
          cVar1S17S47N022N023P043N048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='0' AND D( 5)='0' )then
          cVar1S18S47N022N023P043N048(0) <='1';
          else
          cVar1S18S47N022N023P043N048(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='1' AND A(16)='1' )then
          cVar1S19S47N022N023P043P006nsss(0) <='1';
          else
          cVar1S19S47N022N023P043P006nsss(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='1' AND A(16)='0' )then
          cVar1S20S47N022N023P043N006(0) <='1';
          else
          cVar1S20S47N022N023P043N006(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='1' AND A(16)='0' )then
          cVar1S21S47N022N023P043N006(0) <='1';
          else
          cVar1S21S47N022N023P043N006(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='1' AND A(16)='0' )then
          cVar1S22S47N022N023P043N006(0) <='1';
          else
          cVar1S22S47N022N023P043N006(0) <='0';
          end if;
        if(B(18)='0' AND B( 8)='0' AND E(15)='1' AND A(16)='0' )then
          cVar1S23S47N022N023P043N006(0) <='1';
          else
          cVar1S23S47N022N023P043N006(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='1' )then
          cVar1S0S48P016P065P034P059(0) <='1';
          else
          cVar1S0S48P016P065P034P059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='1' )then
          cVar1S1S48P016P065P034P059(0) <='1';
          else
          cVar1S1S48P016P065P034P059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S2S48P016P065P034N059(0) <='1';
          else
          cVar1S2S48P016P065P034N059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S3S48P016P065P034N059(0) <='1';
          else
          cVar1S3S48P016P065P034N059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S4S48P016P065P034N059(0) <='1';
          else
          cVar1S4S48P016P065P034N059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='0' AND E(11)='0' )then
          cVar1S5S48P016P065P034N059(0) <='1';
          else
          cVar1S5S48P016P065P034N059(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S6S48P016P065P034P014(0) <='1';
          else
          cVar1S6S48P016P065P034P014(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S7S48P016P065P034P014(0) <='1';
          else
          cVar1S7S48P016P065P034P014(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S8S48P016P065P034P014(0) <='1';
          else
          cVar1S8S48P016P065P034P014(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S9S48P016P065P034N014(0) <='1';
          else
          cVar1S9S48P016P065P034N014(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='1' AND E(10)='0' )then
          cVar1S10S48P016P065P067P063nsss(0) <='1';
          else
          cVar1S10S48P016P065P067P063nsss(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='1' AND E(10)='1' )then
          cVar1S11S48P016P065P067P063(0) <='1';
          else
          cVar1S11S48P016P065P067P063(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='1' AND E(10)='1' )then
          cVar1S12S48P016P065P067P063(0) <='1';
          else
          cVar1S12S48P016P065P067P063(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='0' AND E( 1)='0' )then
          cVar1S13S48P016P065N067P066(0) <='1';
          else
          cVar1S13S48P016P065N067P066(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='0' AND E( 1)='0' )then
          cVar1S14S48P016P065N067P066(0) <='1';
          else
          cVar1S14S48P016P065N067P066(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='0' AND E( 1)='0' )then
          cVar1S15S48P016P065N067P066(0) <='1';
          else
          cVar1S15S48P016P065N067P066(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='0' AND E( 1)='1' )then
          cVar1S16S48P016P065N067P066(0) <='1';
          else
          cVar1S16S48P016P065N067P066(0) <='0';
          end if;
        if(A(11)='0' AND D( 9)='1' AND E( 9)='0' AND E( 1)='1' )then
          cVar1S17S48P016P065N067P066(0) <='1';
          else
          cVar1S17S48P016P065N067P066(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='0' AND D(11)='0' )then
          cVar1S18S48P016P063P015P057(0) <='1';
          else
          cVar1S18S48P016P063P015P057(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='0' AND D(11)='0' )then
          cVar1S19S48P016P063P015P057(0) <='1';
          else
          cVar1S19S48P016P063P015P057(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='0' AND D(11)='0' )then
          cVar1S20S48P016P063P015P057(0) <='1';
          else
          cVar1S20S48P016P063P015P057(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='1' AND D( 3)='0' )then
          cVar1S21S48P016P063P015P056(0) <='1';
          else
          cVar1S21S48P016P063P015P056(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='1' AND D( 3)='0' )then
          cVar1S22S48P016P063P015P056(0) <='1';
          else
          cVar1S22S48P016P063P015P056(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='1' AND A( 2)='1' AND D( 3)='0' )then
          cVar1S23S48P016P063P015P056(0) <='1';
          else
          cVar1S23S48P016P063P015P056(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='0' )then
          cVar1S24S48P016N063P052P061(0) <='1';
          else
          cVar1S24S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='0' )then
          cVar1S25S48P016N063P052P061(0) <='1';
          else
          cVar1S25S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='0' )then
          cVar1S26S48P016N063P052P061(0) <='1';
          else
          cVar1S26S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='1' )then
          cVar1S27S48P016N063P052P061(0) <='1';
          else
          cVar1S27S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='1' )then
          cVar1S28S48P016N063P052P061(0) <='1';
          else
          cVar1S28S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='0' AND D(10)='1' )then
          cVar1S29S48P016N063P052P061(0) <='1';
          else
          cVar1S29S48P016N063P052P061(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='1' AND D( 2)='0' )then
          cVar1S30S48P016N063P052P060(0) <='1';
          else
          cVar1S30S48P016N063P052P060(0) <='0';
          end if;
        if(A(11)='1' AND E(10)='0' AND D( 4)='1' AND D( 2)='0' )then
          cVar1S31S48P016N063P052P060(0) <='1';
          else
          cVar1S31S48P016N063P052P060(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='1' AND E( 7)='1' )then
          cVar1S0S49P023P005P042nsss(0) <='1';
          else
          cVar1S0S49P023P005P042nsss(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='1' AND E( 7)='0' AND E(15)='1' )then
          cVar1S1S49P023P005N042P043nsss(0) <='1';
          else
          cVar1S1S49P023P005N042P043nsss(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S2S49P023N005P034P007(0) <='1';
          else
          cVar1S2S49P023N005P034P007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S3S49P023N005P034P007(0) <='1';
          else
          cVar1S3S49P023N005P034P007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S4S49P023N005P034N007(0) <='1';
          else
          cVar1S4S49P023N005P034N007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S5S49P023N005P034N007(0) <='1';
          else
          cVar1S5S49P023N005P034N007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S6S49P023N005P034N007(0) <='1';
          else
          cVar1S6S49P023N005P034N007(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='1' AND A( 7)='1' )then
          cVar1S7S49N023P022P043P005nsss(0) <='1';
          else
          cVar1S7S49N023P022P043P005nsss(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='1' AND A( 7)='0' )then
          cVar1S8S49N023P022P043N005(0) <='1';
          else
          cVar1S8S49N023P022P043N005(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='1' AND A( 7)='0' )then
          cVar1S9S49N023P022P043N005(0) <='1';
          else
          cVar1S9S49N023P022P043N005(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='1' AND A( 7)='0' )then
          cVar1S10S49N023P022P043N005(0) <='1';
          else
          cVar1S10S49N023P022P043N005(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar1S11S49N023P022N043P004nsss(0) <='1';
          else
          cVar1S11S49N023P022N043P004nsss(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='0' AND A(17)='0' )then
          cVar1S12S49N023P022N043N004(0) <='1';
          else
          cVar1S12S49N023P022N043N004(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='0' AND A(17)='0' )then
          cVar1S13S49N023P022N043N004(0) <='1';
          else
          cVar1S13S49N023P022N043N004(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='1' AND E(15)='0' AND A(17)='0' )then
          cVar1S14S49N023P022N043N004(0) <='1';
          else
          cVar1S14S49N023P022N043N004(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='1' AND B( 2)='0' )then
          cVar1S15S49N023N022P016P035(0) <='1';
          else
          cVar1S15S49N023N022P016P035(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='1' AND B( 2)='0' )then
          cVar1S16S49N023N022P016P035(0) <='1';
          else
          cVar1S16S49N023N022P016P035(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='1' AND B( 2)='0' )then
          cVar1S17S49N023N022P016P035(0) <='1';
          else
          cVar1S17S49N023N022P016P035(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='1' AND B( 2)='1' )then
          cVar1S18S49N023N022P016P035(0) <='1';
          else
          cVar1S18S49N023N022P016P035(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='1' )then
          cVar1S19S49N023N022N016P028(0) <='1';
          else
          cVar1S19S49N023N022N016P028(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='1' )then
          cVar1S20S49N023N022N016P028(0) <='1';
          else
          cVar1S20S49N023N022N016P028(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='1' )then
          cVar1S21S49N023N022N016P028(0) <='1';
          else
          cVar1S21S49N023N022N016P028(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='0' )then
          cVar1S22S49N023N022N016N028(0) <='1';
          else
          cVar1S22S49N023N022N016N028(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='0' )then
          cVar1S23S49N023N022N016N028(0) <='1';
          else
          cVar1S23S49N023N022N016N028(0) <='0';
          end if;
        if(B( 8)='0' AND B(18)='0' AND A(11)='0' AND B(15)='0' )then
          cVar1S24S49N023N022N016N028(0) <='1';
          else
          cVar1S24S49N023N022N016N028(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='1' AND E( 7)='1' )then
          cVar1S0S50P023P005P042nsss(0) <='1';
          else
          cVar1S0S50P023P005P042nsss(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='1' AND E( 7)='0' AND E(15)='1' )then
          cVar1S1S50P023P005N042P043nsss(0) <='1';
          else
          cVar1S1S50P023P005N042P043nsss(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S2S50P023N005P034P007(0) <='1';
          else
          cVar1S2S50P023N005P034P007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='1' )then
          cVar1S3S50P023N005P034P007(0) <='1';
          else
          cVar1S3S50P023N005P034P007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S4S50P023N005P034N007(0) <='1';
          else
          cVar1S4S50P023N005P034N007(0) <='0';
          end if;
        if(B( 8)='1' AND A( 7)='0' AND B(12)='0' AND A( 6)='0' )then
          cVar1S5S50P023N005P034N007(0) <='1';
          else
          cVar1S5S50P023N005P034N007(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='1' AND B( 5)='0' AND A(14)='1' )then
          cVar1S6S50N023P028P029P010(0) <='1';
          else
          cVar1S6S50N023P028P029P010(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='1' AND B( 5)='0' AND A(14)='0' )then
          cVar1S7S50N023P028P029N010(0) <='1';
          else
          cVar1S7S50N023P028P029N010(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='1' AND B( 5)='0' AND A(14)='0' )then
          cVar1S8S50N023P028P029N010(0) <='1';
          else
          cVar1S8S50N023P028P029N010(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='1' )then
          cVar1S9S50N023N028P053P025(0) <='1';
          else
          cVar1S9S50N023N028P053P025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='1' )then
          cVar1S10S50N023N028P053P025(0) <='1';
          else
          cVar1S10S50N023N028P053P025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='0' )then
          cVar1S11S50N023N028P053N025(0) <='1';
          else
          cVar1S11S50N023N028P053N025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='0' )then
          cVar1S12S50N023N028P053N025(0) <='1';
          else
          cVar1S12S50N023N028P053N025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='0' )then
          cVar1S13S50N023N028P053N025(0) <='1';
          else
          cVar1S13S50N023N028P053N025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='0' AND B( 7)='0' )then
          cVar1S14S50N023N028P053N025(0) <='1';
          else
          cVar1S14S50N023N028P053N025(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='1' AND B( 5)='1' )then
          cVar1S15S50N023N028P053P029(0) <='1';
          else
          cVar1S15S50N023N028P053P029(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='1' AND B( 5)='1' )then
          cVar1S16S50N023N028P053P029(0) <='1';
          else
          cVar1S16S50N023N028P053P029(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S17S50N023N028P053N029(0) <='1';
          else
          cVar1S17S50N023N028P053N029(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S18S50N023N028P053N029(0) <='1';
          else
          cVar1S18S50N023N028P053N029(0) <='0';
          end if;
        if(B( 8)='0' AND B(15)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S19S50N023N028P053N029(0) <='1';
          else
          cVar1S19S50N023N028P053N029(0) <='0';
          end if;
        if(B(15)='1' AND B( 5)='0' AND A(14)='1' AND B( 4)='0' )then
          cVar1S0S51P028P029P010P031(0) <='1';
          else
          cVar1S0S51P028P029P010P031(0) <='0';
          end if;
        if(B(15)='1' AND B( 5)='0' AND A(14)='1' AND B( 4)='0' )then
          cVar1S1S51P028P029P010P031(0) <='1';
          else
          cVar1S1S51P028P029P010P031(0) <='0';
          end if;
        if(B(15)='1' AND B( 5)='0' AND A(14)='1' AND B( 4)='0' )then
          cVar1S2S51P028P029P010P031(0) <='1';
          else
          cVar1S2S51P028P029P010P031(0) <='0';
          end if;
        if(B(15)='1' AND B( 5)='0' AND A(14)='0' AND A(15)='1' )then
          cVar1S3S51P028P029N010P008nsss(0) <='1';
          else
          cVar1S3S51P028P029N010P008nsss(0) <='0';
          end if;
        if(B(15)='1' AND B( 5)='0' AND A(14)='0' AND A(15)='0' )then
          cVar1S4S51P028P029N010N008(0) <='1';
          else
          cVar1S4S51P028P029N010N008(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='1' AND A( 7)='1' AND E( 7)='1' )then
          cVar1S5S51N028P023P005P042nsss(0) <='1';
          else
          cVar1S5S51N028P023P005P042nsss(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='1' AND A( 7)='1' AND E( 7)='0' )then
          cVar1S6S51N028P023P005N042(0) <='1';
          else
          cVar1S6S51N028P023P005N042(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='1' AND A( 7)='0' AND D(13)='0' )then
          cVar1S7S51N028P023N005P049(0) <='1';
          else
          cVar1S7S51N028P023N005P049(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='1' AND A( 7)='0' AND D(13)='0' )then
          cVar1S8S51N028P023N005P049(0) <='1';
          else
          cVar1S8S51N028P023N005P049(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S9S51N028N023P025P007nsss(0) <='1';
          else
          cVar1S9S51N028N023P025P007nsss(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S10S51N028N023P025N007(0) <='1';
          else
          cVar1S10S51N028N023P025N007(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S11S51N028N023P025N007(0) <='1';
          else
          cVar1S11S51N028N023P025N007(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S12S51N028N023N025P024(0) <='1';
          else
          cVar1S12S51N028N023N025P024(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S13S51N028N023N025P024(0) <='1';
          else
          cVar1S13S51N028N023N025P024(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S14S51N028N023N025P024(0) <='1';
          else
          cVar1S14S51N028N023N025P024(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S15S51N028N023N025N024(0) <='1';
          else
          cVar1S15S51N028N023N025N024(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S16S51N028N023N025N024(0) <='1';
          else
          cVar1S16S51N028N023N025N024(0) <='0';
          end if;
        if(B(15)='0' AND B( 8)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S17S51N028N023N025N024(0) <='1';
          else
          cVar1S17S51N028N023N025N024(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S0S52P045P043P005P068nsss(0) <='1';
          else
          cVar1S0S52P045P043P005P068nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S1S52P045P043N005P004nsss(0) <='1';
          else
          cVar1S1S52P045P043N005P004nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S2S52P045P043N005N004(0) <='1';
          else
          cVar1S2S52P045P043N005N004(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S3S52P045P043N005N004(0) <='1';
          else
          cVar1S3S52P045P043N005N004(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S4S52P045P043N005N004(0) <='1';
          else
          cVar1S4S52P045P043N005N004(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='1' AND A(16)='1' )then
          cVar1S5S52P045N043P047P006nsss(0) <='1';
          else
          cVar1S5S52P045N043P047P006nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='1' AND A(16)='0' )then
          cVar1S6S52P045N043P047N006(0) <='1';
          else
          cVar1S6S52P045N043P047N006(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='1' AND A(16)='0' )then
          cVar1S7S52P045N043P047N006(0) <='1';
          else
          cVar1S7S52P045N043P047N006(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='0' AND D( 5)='1' )then
          cVar1S8S52P045N043N047P048nsss(0) <='1';
          else
          cVar1S8S52P045N043N047P048nsss(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='0' AND D( 5)='0' )then
          cVar1S9S52P045N043N047N048(0) <='1';
          else
          cVar1S9S52P045N043N047N048(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='0' AND D( 5)='0' )then
          cVar1S10S52P045N043N047N048(0) <='1';
          else
          cVar1S10S52P045N043N047N048(0) <='0';
          end if;
        if(D(14)='1' AND E(15)='0' AND E(14)='0' AND D( 5)='0' )then
          cVar1S11S52P045N043N047N048(0) <='1';
          else
          cVar1S11S52P045N043N047N048(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='1' AND E(12)='1' )then
          cVar1S12S52N045P028P010P055(0) <='1';
          else
          cVar1S12S52N045P028P010P055(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='1' AND E(12)='0' )then
          cVar1S13S52N045P028P010N055(0) <='1';
          else
          cVar1S13S52N045P028P010N055(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='1' AND E(12)='0' )then
          cVar1S14S52N045P028P010N055(0) <='1';
          else
          cVar1S14S52N045P028P010N055(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar1S15S52N045P028N010P011(0) <='1';
          else
          cVar1S15S52N045P028N010P011(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar1S16S52N045P028N010P011(0) <='1';
          else
          cVar1S16S52N045P028N010P011(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar1S17S52N045P028N010P011(0) <='1';
          else
          cVar1S17S52N045P028N010P011(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='0' AND A( 4)='0' )then
          cVar1S18S52N045P028N010N011(0) <='1';
          else
          cVar1S18S52N045P028N010N011(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='1' AND A(14)='0' AND A( 4)='0' )then
          cVar1S19S52N045P028N010N011(0) <='1';
          else
          cVar1S19S52N045P028N010N011(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S20S52N045N028P040P021(0) <='1';
          else
          cVar1S20S52N045N028P040P021(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S21S52N045N028P040P021(0) <='1';
          else
          cVar1S21S52N045N028P040P021(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S22S52N045N028P040N021(0) <='1';
          else
          cVar1S22S52N045N028P040N021(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S23S52N045N028P040N021(0) <='1';
          else
          cVar1S23S52N045N028P040N021(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='1' )then
          cVar1S24S52N045N028N040P025(0) <='1';
          else
          cVar1S24S52N045N028N040P025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='1' )then
          cVar1S25S52N045N028N040P025(0) <='1';
          else
          cVar1S25S52N045N028N040P025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='1' )then
          cVar1S26S52N045N028N040P025(0) <='1';
          else
          cVar1S26S52N045N028N040P025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='0' )then
          cVar1S27S52N045N028N040N025(0) <='1';
          else
          cVar1S27S52N045N028N040N025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='0' )then
          cVar1S28S52N045N028N040N025(0) <='1';
          else
          cVar1S28S52N045N028N040N025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='0' )then
          cVar1S29S52N045N028N040N025(0) <='1';
          else
          cVar1S29S52N045N028N040N025(0) <='0';
          end if;
        if(D(14)='0' AND B(15)='0' AND D( 7)='0' AND B( 7)='0' )then
          cVar1S30S52N045N028N040N025(0) <='1';
          else
          cVar1S30S52N045N028N040N025(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='1' AND E( 1)='0' )then
          cVar1S0S53P025P007P066nsss(0) <='1';
          else
          cVar1S0S53P025P007P066nsss(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='1' AND E( 1)='1' AND B( 1)='1' )then
          cVar1S1S53P025P007P066P037nsss(0) <='1';
          else
          cVar1S1S53P025P007P066P037nsss(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='0' AND E( 6)='1' AND A(17)='1' )then
          cVar1S2S53P025N007P046P004nsss(0) <='1';
          else
          cVar1S2S53P025N007P046P004nsss(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='0' AND E( 6)='1' AND A(17)='0' )then
          cVar1S3S53P025N007P046N004(0) <='1';
          else
          cVar1S3S53P025N007P046N004(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='0' AND E( 6)='1' AND A(17)='0' )then
          cVar1S4S53P025N007P046N004(0) <='1';
          else
          cVar1S4S53P025N007P046N004(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='0' AND E( 6)='0' AND A( 8)='0' )then
          cVar1S5S53P025N007N046P003(0) <='1';
          else
          cVar1S5S53P025N007N046P003(0) <='0';
          end if;
        if(B( 7)='1' AND A( 6)='0' AND E( 6)='0' AND A( 8)='0' )then
          cVar1S6S53P025N007N046P003(0) <='1';
          else
          cVar1S6S53P025N007N046P003(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='1' AND E(12)='1' )then
          cVar1S7S53N025P028P010P055nsss(0) <='1';
          else
          cVar1S7S53N025P028P010P055nsss(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='1' AND E(12)='0' )then
          cVar1S8S53N025P028P010N055(0) <='1';
          else
          cVar1S8S53N025P028P010N055(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='1' AND E(12)='0' )then
          cVar1S9S53N025P028P010N055(0) <='1';
          else
          cVar1S9S53N025P028P010N055(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='0' AND B( 5)='0' )then
          cVar1S10S53N025P028N010P029(0) <='1';
          else
          cVar1S10S53N025P028N010P029(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='0' AND B( 5)='0' )then
          cVar1S11S53N025P028N010P029(0) <='1';
          else
          cVar1S11S53N025P028N010P029(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='1' AND A(14)='0' AND B( 5)='1' )then
          cVar1S12S53N025P028N010P029(0) <='1';
          else
          cVar1S12S53N025P028N010P029(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S13S53N025N028P040P021(0) <='1';
          else
          cVar1S13S53N025N028P040P021(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S14S53N025N028P040P021(0) <='1';
          else
          cVar1S14S53N025N028P040P021(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S15S53N025N028P040N021(0) <='1';
          else
          cVar1S15S53N025N028P040N021(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S16S53N025N028P040N021(0) <='1';
          else
          cVar1S16S53N025N028P040N021(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='1' )then
          cVar1S17S53N025N028N040P045(0) <='1';
          else
          cVar1S17S53N025N028N040P045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='1' )then
          cVar1S18S53N025N028N040P045(0) <='1';
          else
          cVar1S18S53N025N028N040P045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='1' )then
          cVar1S19S53N025N028N040P045(0) <='1';
          else
          cVar1S19S53N025N028N040P045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='0' )then
          cVar1S20S53N025N028N040N045(0) <='1';
          else
          cVar1S20S53N025N028N040N045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='0' )then
          cVar1S21S53N025N028N040N045(0) <='1';
          else
          cVar1S21S53N025N028N040N045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='0' )then
          cVar1S22S53N025N028N040N045(0) <='1';
          else
          cVar1S22S53N025N028N040N045(0) <='0';
          end if;
        if(B( 7)='0' AND B(15)='0' AND D( 7)='0' AND D(14)='0' )then
          cVar1S23S53N025N028N040N045(0) <='1';
          else
          cVar1S23S53N025N028N040N045(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S0S54P018P040P002nsss(0) <='1';
          else
          cVar1S0S54P018P040P002nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S1S54P018P040N002P004nsss(0) <='1';
          else
          cVar1S1S54P018P040N002P004nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S2S54P018P040N002N004(0) <='1';
          else
          cVar1S2S54P018P040N002N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S3S54P018P040N002N004(0) <='1';
          else
          cVar1S3S54P018P040N002N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S4S54P018P040N002N004(0) <='1';
          else
          cVar1S4S54P018P040N002N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='1' AND A(17)='1' )then
          cVar1S5S54P018N040P045P004nsss(0) <='1';
          else
          cVar1S5S54P018N040P045P004nsss(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S6S54P018N040P045N004(0) <='1';
          else
          cVar1S6S54P018N040P045N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S7S54P018N040P045N004(0) <='1';
          else
          cVar1S7S54P018N040P045N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S8S54P018N040P045N004(0) <='1';
          else
          cVar1S8S54P018N040P045N004(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='0' AND A( 2)='1' )then
          cVar1S9S54P018N040N045P015(0) <='1';
          else
          cVar1S9S54P018N040N045P015(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='0' AND A( 2)='1' )then
          cVar1S10S54P018N040N045P015(0) <='1';
          else
          cVar1S10S54P018N040N045P015(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='0' AND A( 2)='0' )then
          cVar1S11S54P018N040N045N015(0) <='1';
          else
          cVar1S11S54P018N040N045N015(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='0' AND A( 2)='0' )then
          cVar1S12S54P018N040N045N015(0) <='1';
          else
          cVar1S12S54P018N040N045N015(0) <='0';
          end if;
        if(A(10)='0' AND D( 7)='0' AND D(14)='0' AND A( 2)='0' )then
          cVar1S13S54P018N040N045N015(0) <='1';
          else
          cVar1S13S54P018N040N045N015(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S14S54P018P015P019P056(0) <='1';
          else
          cVar1S14S54P018P015P019P056(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S15S54P018P015P019P056(0) <='1';
          else
          cVar1S15S54P018P015P019P056(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S16S54P018P015P019P056(0) <='1';
          else
          cVar1S16S54P018P015P019P056(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S17S54P018P015P019P056(0) <='1';
          else
          cVar1S17S54P018P015P019P056(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='1' AND A( 0)='0' AND D(12)='1' )then
          cVar1S18S54P018P015N019P053nsss(0) <='1';
          else
          cVar1S18S54P018P015N019P053nsss(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='0' AND A( 6)='0' )then
          cVar1S19S54P018N015P019P007(0) <='1';
          else
          cVar1S19S54P018N015P019P007(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='0' AND A( 6)='0' )then
          cVar1S20S54P018N015P019P007(0) <='1';
          else
          cVar1S20S54P018N015P019P007(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='0' AND A( 6)='1' )then
          cVar1S21S54P018N015P019P007(0) <='1';
          else
          cVar1S21S54P018N015P019P007(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='0' AND A( 6)='1' )then
          cVar1S22S54P018N015P019P007(0) <='1';
          else
          cVar1S22S54P018N015P019P007(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='1' AND E(11)='1' )then
          cVar1S23S54P018N015P019P059(0) <='1';
          else
          cVar1S23S54P018N015P019P059(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='1' AND E(11)='1' )then
          cVar1S24S54P018N015P019P059(0) <='1';
          else
          cVar1S24S54P018N015P019P059(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='1' AND E(11)='0' )then
          cVar1S25S54P018N015P019N059(0) <='1';
          else
          cVar1S25S54P018N015P019N059(0) <='0';
          end if;
        if(A(10)='1' AND A( 2)='0' AND A( 0)='1' AND E(11)='0' )then
          cVar1S26S54P018N015P019N059(0) <='1';
          else
          cVar1S26S54P018N015P019N059(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' )then
          cVar1S0S55P040P002nsss(0) <='1';
          else
          cVar1S0S55P040P002nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='0' AND B( 9)='1' )then
          cVar1S1S55P040N002P015P021(0) <='1';
          else
          cVar1S1S55P040N002P015P021(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='0' AND B( 9)='1' )then
          cVar1S2S55P040N002P015P021(0) <='1';
          else
          cVar1S2S55P040N002P015P021(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='0' AND B( 9)='0' )then
          cVar1S3S55P040N002P015N021(0) <='1';
          else
          cVar1S3S55P040N002P015N021(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='0' AND B( 9)='0' )then
          cVar1S4S55P040N002P015N021(0) <='1';
          else
          cVar1S4S55P040N002P015N021(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='0' AND B( 9)='0' )then
          cVar1S5S55P040N002P015N021(0) <='1';
          else
          cVar1S5S55P040N002P015N021(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='1' AND A( 3)='1' )then
          cVar1S6S55P040N002P015P013nsss(0) <='1';
          else
          cVar1S6S55P040N002P015P013nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A( 2)='1' AND A( 3)='0' )then
          cVar1S7S55P040N002P015N013(0) <='1';
          else
          cVar1S7S55P040N002P015N013(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S8S55N040P045P005P068(0) <='1';
          else
          cVar1S8S55N040P045P005P068(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S9S55N040P045N005P004(0) <='1';
          else
          cVar1S9S55N040P045N005P004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S10S55N040P045N005P004(0) <='1';
          else
          cVar1S10S55N040P045N005P004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S11S55N040P045N005N004(0) <='1';
          else
          cVar1S11S55N040P045N005N004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S12S55N040P045N005N004(0) <='1';
          else
          cVar1S12S55N040P045N005N004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S13S55N040P045N005N004(0) <='1';
          else
          cVar1S13S55N040P045N005N004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S14S55N040P045N005N004(0) <='1';
          else
          cVar1S14S55N040P045N005N004(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='1' AND E(14)='0' )then
          cVar1S15S55N040N045P015P047(0) <='1';
          else
          cVar1S15S55N040N045P015P047(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='1' AND E(14)='0' )then
          cVar1S16S55N040N045P015P047(0) <='1';
          else
          cVar1S16S55N040N045P015P047(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='1' AND E(14)='0' )then
          cVar1S17S55N040N045P015P047(0) <='1';
          else
          cVar1S17S55N040N045P015P047(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='1' AND E(14)='0' )then
          cVar1S18S55N040N045P015P047(0) <='1';
          else
          cVar1S18S55N040N045P015P047(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='1' AND E(14)='1' )then
          cVar1S19S55N040N045P015P047(0) <='1';
          else
          cVar1S19S55N040N045P015P047(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='1' )then
          cVar1S20S55N040N045N015P028(0) <='1';
          else
          cVar1S20S55N040N045N015P028(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='1' )then
          cVar1S21S55N040N045N015P028(0) <='1';
          else
          cVar1S21S55N040N045N015P028(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='0' )then
          cVar1S22S55N040N045N015N028(0) <='1';
          else
          cVar1S22S55N040N045N015N028(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='0' )then
          cVar1S23S55N040N045N015N028(0) <='1';
          else
          cVar1S23S55N040N045N015N028(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='0' )then
          cVar1S24S55N040N045N015N028(0) <='1';
          else
          cVar1S24S55N040N045N015N028(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND A( 2)='0' AND B(15)='0' )then
          cVar1S25S55N040N045N015N028(0) <='1';
          else
          cVar1S25S55N040N045N015N028(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND D( 0)='0' AND A(13)='0' )then
          cVar1S0S56P045P005P068P012nsss(0) <='1';
          else
          cVar1S0S56P045P005P068P012nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='1' AND A( 3)='0' )then
          cVar1S1S56P045N005P004P013nsss(0) <='1';
          else
          cVar1S1S56P045N005P004P013nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S2S56P045N005N004P006(0) <='1';
          else
          cVar1S2S56P045N005N004P006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S3S56P045N005N004P006(0) <='1';
          else
          cVar1S3S56P045N005N004P006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S4S56P045N005N004N006(0) <='1';
          else
          cVar1S4S56P045N005N004N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S5S56P045N005N004N006(0) <='1';
          else
          cVar1S5S56P045N005N004N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S6S56P045N005N004N006(0) <='1';
          else
          cVar1S6S56P045N005N004N006(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='1' )then
          cVar1S7S56N045P040P021P002nsss(0) <='1';
          else
          cVar1S7S56N045P040P021P002nsss(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S8S56N045P040P021N002(0) <='1';
          else
          cVar1S8S56N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND E( 1)='0' )then
          cVar1S9S56N045P040N021P066(0) <='1';
          else
          cVar1S9S56N045P040N021P066(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND E( 1)='0' )then
          cVar1S10S56N045P040N021P066(0) <='1';
          else
          cVar1S10S56N045P040N021P066(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S11S56N045N040P018P043(0) <='1';
          else
          cVar1S11S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S12S56N045N040P018P043(0) <='1';
          else
          cVar1S12S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S13S56N045N040P018P043(0) <='1';
          else
          cVar1S13S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='1' )then
          cVar1S14S56N045N040P018P043(0) <='1';
          else
          cVar1S14S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='1' )then
          cVar1S15S56N045N040P018P043(0) <='1';
          else
          cVar1S15S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='1' )then
          cVar1S16S56N045N040P018P043(0) <='1';
          else
          cVar1S16S56N045N040P018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S17S56N045N040P018P060(0) <='1';
          else
          cVar1S17S56N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S18S56N045N040P018P060(0) <='1';
          else
          cVar1S18S56N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S19S56N045N040P018P060(0) <='1';
          else
          cVar1S19S56N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S20S56N045N040P018P060(0) <='1';
          else
          cVar1S20S56N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S21S56N045N040P018P060(0) <='1';
          else
          cVar1S21S56N045N040P018P060(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND B( 1)='0' )then
          cVar1S0S57P045P005P037nsss(0) <='1';
          else
          cVar1S0S57P045P005P037nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='1' AND A( 3)='0' )then
          cVar1S1S57P045N005P004P013nsss(0) <='1';
          else
          cVar1S1S57P045N005P004P013nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S2S57P045N005N004P006(0) <='1';
          else
          cVar1S2S57P045N005N004P006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar1S3S57P045N005N004P006(0) <='1';
          else
          cVar1S3S57P045N005N004P006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S4S57P045N005N004N006(0) <='1';
          else
          cVar1S4S57P045N005N004N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S5S57P045N005N004N006(0) <='1';
          else
          cVar1S5S57P045N005N004N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND A(17)='0' AND A(16)='0' )then
          cVar1S6S57P045N005N004N006(0) <='1';
          else
          cVar1S6S57P045N005N004N006(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='1' )then
          cVar1S7S57N045P040P021P002nsss(0) <='1';
          else
          cVar1S7S57N045P040P021P002nsss(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S8S57N045P040P021N002(0) <='1';
          else
          cVar1S8S57N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S9S57N045P040P021N002(0) <='1';
          else
          cVar1S9S57N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S10S57N045P040P021N002(0) <='1';
          else
          cVar1S10S57N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='1' )then
          cVar1S11S57N045P040N021P020(0) <='1';
          else
          cVar1S11S57N045P040N021P020(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S12S57N045P040N021N020(0) <='1';
          else
          cVar1S12S57N045P040N021N020(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND B(19)='0' )then
          cVar1S13S57N045P040N021N020(0) <='1';
          else
          cVar1S13S57N045P040N021N020(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S14S57N045N040P018P060(0) <='1';
          else
          cVar1S14S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S15S57N045N040P018P060(0) <='1';
          else
          cVar1S15S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S16S57N045N040P018P060(0) <='1';
          else
          cVar1S16S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S17S57N045N040P018P060(0) <='1';
          else
          cVar1S17S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S18S57N045N040P018P060(0) <='1';
          else
          cVar1S18S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S19S57N045N040P018P060(0) <='1';
          else
          cVar1S19S57N045N040P018P060(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S20S57N045N040N018P043(0) <='1';
          else
          cVar1S20S57N045N040N018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S21S57N045N040N018P043(0) <='1';
          else
          cVar1S21S57N045N040N018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='0' )then
          cVar1S22S57N045N040N018P043(0) <='1';
          else
          cVar1S22S57N045N040N018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='1' )then
          cVar1S23S57N045N040N018P043(0) <='1';
          else
          cVar1S23S57N045N040N018P043(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND A(10)='0' AND E(15)='1' )then
          cVar1S24S57N045N040N018P043(0) <='1';
          else
          cVar1S24S57N045N040N018P043(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S0S58P045P005P068nsss(0) <='1';
          else
          cVar1S0S58P045P005P068nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A(16)='1' )then
          cVar1S1S58P045N005P021P006(0) <='1';
          else
          cVar1S1S58P045N005P021P006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A(16)='0' )then
          cVar1S2S58P045N005P021N006(0) <='1';
          else
          cVar1S2S58P045N005P021N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A(16)='0' )then
          cVar1S3S58P045N005P021N006(0) <='1';
          else
          cVar1S3S58P045N005P021N006(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A(16)='0' )then
          cVar1S4S58P045N005P021N006(0) <='1';
          else
          cVar1S4S58P045N005P021N006(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S5S58N045P018P040P002nsss(0) <='1';
          else
          cVar1S5S58N045P018P040P002nsss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S6S58N045P018P040N002(0) <='1';
          else
          cVar1S6S58N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S7S58N045P018P040N002(0) <='1';
          else
          cVar1S7S58N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S8S58N045P018P040N002(0) <='1';
          else
          cVar1S8S58N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S9S58N045P018N040P043(0) <='1';
          else
          cVar1S9S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S10S58N045P018N040P043(0) <='1';
          else
          cVar1S10S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S11S58N045P018N040P043(0) <='1';
          else
          cVar1S11S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S12S58N045P018N040P043(0) <='1';
          else
          cVar1S12S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S13S58N045P018N040P043(0) <='1';
          else
          cVar1S13S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S14S58N045P018N040P043(0) <='1';
          else
          cVar1S14S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S15S58N045P018N040P043(0) <='1';
          else
          cVar1S15S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S16S58N045P018N040P043(0) <='1';
          else
          cVar1S16S58N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S17S58N045P018P019P056(0) <='1';
          else
          cVar1S17S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S18S58N045P018P019P056(0) <='1';
          else
          cVar1S18S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S19S58N045P018P019P056(0) <='1';
          else
          cVar1S19S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S20S58N045P018P019P056(0) <='1';
          else
          cVar1S20S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S21S58N045P018P019P056(0) <='1';
          else
          cVar1S21S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S22S58N045P018P019P056(0) <='1';
          else
          cVar1S22S58N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S23S58N045P018N019P024(0) <='1';
          else
          cVar1S23S58N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S24S58N045P018N019P024(0) <='1';
          else
          cVar1S24S58N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='1' )then
          cVar1S25S58N045P018N019P024(0) <='1';
          else
          cVar1S25S58N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='1' )then
          cVar1S26S58N045P018N019P024(0) <='1';
          else
          cVar1S26S58N045P018N019P024(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='1' AND A( 0)='1' )then
          cVar1S0S59P045P022P019nsss(0) <='1';
          else
          cVar1S0S59P045P022P019nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='1' AND A( 0)='0' AND A( 3)='0' )then
          cVar1S1S59P045P022N019P013nsss(0) <='1';
          else
          cVar1S1S59P045P022N019P013nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='0' AND B( 8)='1' )then
          cVar1S2S59P045N022P023nsss(0) <='1';
          else
          cVar1S2S59P045N022P023nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='0' AND B( 8)='0' AND A(16)='1' )then
          cVar1S3S59P045N022N023P006(0) <='1';
          else
          cVar1S3S59P045N022N023P006(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='0' AND B( 8)='0' AND A(16)='0' )then
          cVar1S4S59P045N022N023N006(0) <='1';
          else
          cVar1S4S59P045N022N023N006(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='0' AND B( 8)='0' AND A(16)='0' )then
          cVar1S5S59P045N022N023N006(0) <='1';
          else
          cVar1S5S59P045N022N023N006(0) <='0';
          end if;
        if(D(14)='1' AND B(18)='0' AND B( 8)='0' AND A(16)='0' )then
          cVar1S6S59P045N022N023N006(0) <='1';
          else
          cVar1S6S59P045N022N023N006(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='1' )then
          cVar1S7S59N045P040P021P002nsss(0) <='1';
          else
          cVar1S7S59N045P040P021P002nsss(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S8S59N045P040P021N002(0) <='1';
          else
          cVar1S8S59N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S9S59N045P040P021N002(0) <='1';
          else
          cVar1S9S59N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S10S59N045P040P021N002(0) <='1';
          else
          cVar1S10S59N045P040P021N002(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND E( 1)='0' )then
          cVar1S11S59N045P040N021P066nsss(0) <='1';
          else
          cVar1S11S59N045P040N021P066nsss(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='1' AND B( 9)='0' AND E( 1)='1' )then
          cVar1S12S59N045P040N021P066(0) <='1';
          else
          cVar1S12S59N045P040N021P066(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='1' AND A( 6)='1' )then
          cVar1S13S59N045N040P025P007(0) <='1';
          else
          cVar1S13S59N045N040P025P007(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S14S59N045N040P025N007(0) <='1';
          else
          cVar1S14S59N045N040P025N007(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S15S59N045N040P025N007(0) <='1';
          else
          cVar1S15S59N045N040P025N007(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='1' AND A( 6)='0' )then
          cVar1S16S59N045N040P025N007(0) <='1';
          else
          cVar1S16S59N045N040P025N007(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='0' AND A(10)='1' )then
          cVar1S17S59N045N040N025P018(0) <='1';
          else
          cVar1S17S59N045N040N025P018(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='0' AND A(10)='1' )then
          cVar1S18S59N045N040N025P018(0) <='1';
          else
          cVar1S18S59N045N040N025P018(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='0' AND A(10)='0' )then
          cVar1S19S59N045N040N025N018(0) <='1';
          else
          cVar1S19S59N045N040N025N018(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='0' AND A(10)='0' )then
          cVar1S20S59N045N040N025N018(0) <='1';
          else
          cVar1S20S59N045N040N025N018(0) <='0';
          end if;
        if(D(14)='0' AND D( 7)='0' AND B( 7)='0' AND A(10)='0' )then
          cVar1S21S59N045N040N025N018(0) <='1';
          else
          cVar1S21S59N045N040N025N018(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND B( 1)='0' )then
          cVar1S0S60P045P005P037nsss(0) <='1';
          else
          cVar1S0S60P045P005P037nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='1' )then
          cVar1S1S60P045N005P021P024(0) <='1';
          else
          cVar1S1S60P045N005P021P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='1' )then
          cVar1S2S60P045N005P021P024(0) <='1';
          else
          cVar1S2S60P045N005P021P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='1' )then
          cVar1S3S60P045N005P021P024(0) <='1';
          else
          cVar1S3S60P045N005P021P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='0' )then
          cVar1S4S60P045N005P021N024psss(0) <='1';
          else
          cVar1S4S60P045N005P021N024psss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S5S60N045P018P040P002(0) <='1';
          else
          cVar1S5S60N045P018P040P002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S6S60N045P018P040P002(0) <='1';
          else
          cVar1S6S60N045P018P040P002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S7S60N045P018P040P002(0) <='1';
          else
          cVar1S7S60N045P018P040P002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S8S60N045P018P040N002(0) <='1';
          else
          cVar1S8S60N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S9S60N045P018P040N002(0) <='1';
          else
          cVar1S9S60N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S10S60N045P018P040N002(0) <='1';
          else
          cVar1S10S60N045P018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S11S60N045P018N040P043(0) <='1';
          else
          cVar1S11S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S12S60N045P018N040P043(0) <='1';
          else
          cVar1S12S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S13S60N045P018N040P043(0) <='1';
          else
          cVar1S13S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='0' )then
          cVar1S14S60N045P018N040P043(0) <='1';
          else
          cVar1S14S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S15S60N045P018N040P043(0) <='1';
          else
          cVar1S15S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S16S60N045P018N040P043(0) <='1';
          else
          cVar1S16S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND E(15)='1' )then
          cVar1S17S60N045P018N040P043(0) <='1';
          else
          cVar1S17S60N045P018N040P043(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='1' AND B( 2)='1' )then
          cVar1S18S60N045P018P025P035nsss(0) <='1';
          else
          cVar1S18S60N045P018P025P035nsss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='1' AND B( 2)='0' )then
          cVar1S19S60N045P018P025N035(0) <='1';
          else
          cVar1S19S60N045P018P025N035(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='1' AND B( 2)='0' )then
          cVar1S20S60N045P018P025N035(0) <='1';
          else
          cVar1S20S60N045P018P025N035(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='0' AND B( 1)='0' )then
          cVar1S21S60N045P018N025P037(0) <='1';
          else
          cVar1S21S60N045P018N025P037(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='0' AND B( 1)='0' )then
          cVar1S22S60N045P018N025P037(0) <='1';
          else
          cVar1S22S60N045P018N025P037(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='0' AND B( 1)='1' )then
          cVar1S23S60N045P018N025P037(0) <='1';
          else
          cVar1S23S60N045P018N025P037(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='0' AND B( 1)='1' )then
          cVar1S24S60N045P018N025P037(0) <='1';
          else
          cVar1S24S60N045P018N025P037(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 7)='0' AND B( 1)='1' )then
          cVar1S25S60N045P018N025P037(0) <='1';
          else
          cVar1S25S60N045P018N025P037(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND D( 0)='0' AND A(13)='0' )then
          cVar1S0S61P045P005P068P012nsss(0) <='1';
          else
          cVar1S0S61P045P005P068P012nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='1' )then
          cVar1S1S61P045N005P021P024(0) <='1';
          else
          cVar1S1S61P045N005P021P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='1' )then
          cVar1S2S61P045N005P021P024(0) <='1';
          else
          cVar1S2S61P045N005P021P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='0' )then
          cVar1S3S61P045N005P021N024(0) <='1';
          else
          cVar1S3S61P045N005P021N024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='0' )then
          cVar1S4S61P045N005P021N024(0) <='1';
          else
          cVar1S4S61P045N005P021N024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND B(17)='0' )then
          cVar1S5S61P045N005P021N024(0) <='1';
          else
          cVar1S5S61P045N005P021N024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='1' )then
          cVar1S6S61N045P018P037P061(0) <='1';
          else
          cVar1S6S61N045P018P037P061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='1' )then
          cVar1S7S61N045P018P037P061(0) <='1';
          else
          cVar1S7S61N045P018P037P061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='1' )then
          cVar1S8S61N045P018P037P061(0) <='1';
          else
          cVar1S8S61N045P018P037P061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='0' )then
          cVar1S9S61N045P018P037N061(0) <='1';
          else
          cVar1S9S61N045P018P037N061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='0' )then
          cVar1S10S61N045P018P037N061(0) <='1';
          else
          cVar1S10S61N045P018P037N061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='0' AND D(10)='0' )then
          cVar1S11S61N045P018P037N061(0) <='1';
          else
          cVar1S11S61N045P018P037N061(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='1' AND E( 1)='0' )then
          cVar1S12S61N045P018P037P066(0) <='1';
          else
          cVar1S12S61N045P018P037P066(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='1' AND E( 1)='0' )then
          cVar1S13S61N045P018P037P066(0) <='1';
          else
          cVar1S13S61N045P018P037P066(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='1' AND E( 1)='1' )then
          cVar1S14S61N045P018P037P066(0) <='1';
          else
          cVar1S14S61N045P018P037P066(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND B( 1)='1' AND E( 1)='1' )then
          cVar1S15S61N045P018P037P066(0) <='1';
          else
          cVar1S15S61N045P018P037P066(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S16S61N045N018P040P002nsss(0) <='1';
          else
          cVar1S16S61N045N018P040P002nsss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S17S61N045N018P040N002(0) <='1';
          else
          cVar1S17S61N045N018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='1' AND A(18)='0' )then
          cVar1S18S61N045N018P040N002(0) <='1';
          else
          cVar1S18S61N045N018P040N002(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND A(19)='0' )then
          cVar1S19S61N045N018N040P000(0) <='1';
          else
          cVar1S19S61N045N018N040P000(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND A(19)='0' )then
          cVar1S20S61N045N018N040P000(0) <='1';
          else
          cVar1S20S61N045N018N040P000(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND A(19)='0' )then
          cVar1S21S61N045N018N040P000(0) <='1';
          else
          cVar1S21S61N045N018N040P000(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND D( 7)='0' AND A(19)='1' )then
          cVar1S22S61N045N018N040P000(0) <='1';
          else
          cVar1S22S61N045N018N040P000(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar1S0S62P045P005P068nsss(0) <='1';
          else
          cVar1S0S62P045P005P068nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='1' )then
          cVar1S1S62P045N005P027P024(0) <='1';
          else
          cVar1S1S62P045N005P027P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='1' )then
          cVar1S2S62P045N005P027P024(0) <='1';
          else
          cVar1S2S62P045N005P027P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='1' )then
          cVar1S3S62P045N005P027P024(0) <='1';
          else
          cVar1S3S62P045N005P027P024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='0' )then
          cVar1S4S62P045N005P027N024(0) <='1';
          else
          cVar1S4S62P045N005P027N024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='0' )then
          cVar1S5S62P045N005P027N024(0) <='1';
          else
          cVar1S5S62P045N005P027N024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='0' )then
          cVar1S6S62P045N005P027N024(0) <='1';
          else
          cVar1S6S62P045N005P027N024(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 6)='0' AND B(17)='0' )then
          cVar1S7S62P045N005P027N024(0) <='1';
          else
          cVar1S7S62P045N005P027N024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='1' )then
          cVar1S8S62N045P018P000P030(0) <='1';
          else
          cVar1S8S62N045P018P000P030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='1' )then
          cVar1S9S62N045P018P000P030(0) <='1';
          else
          cVar1S9S62N045P018P000P030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='0' )then
          cVar1S10S62N045P018P000N030(0) <='1';
          else
          cVar1S10S62N045P018P000N030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='0' )then
          cVar1S11S62N045P018P000N030(0) <='1';
          else
          cVar1S11S62N045P018P000N030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='0' )then
          cVar1S12S62N045P018P000N030(0) <='1';
          else
          cVar1S12S62N045P018P000N030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='0' AND B(14)='0' )then
          cVar1S13S62N045P018P000N030(0) <='1';
          else
          cVar1S13S62N045P018P000N030(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='1' AND D( 7)='1' )then
          cVar1S14S62N045P018P000P040nsss(0) <='1';
          else
          cVar1S14S62N045P018P000P040nsss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='1' AND D( 7)='0' )then
          cVar1S15S62N045P018P000N040(0) <='1';
          else
          cVar1S15S62N045P018P000N040(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND A(19)='1' AND D( 7)='0' )then
          cVar1S16S62N045P018P000N040(0) <='1';
          else
          cVar1S16S62N045P018P000N040(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='1' AND B( 2)='1' )then
          cVar1S17S62N045P018P061P035nsss(0) <='1';
          else
          cVar1S17S62N045P018P061P035nsss(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='1' AND B( 2)='0' )then
          cVar1S18S62N045P018P061N035(0) <='1';
          else
          cVar1S18S62N045P018P061N035(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='1' AND B( 2)='0' )then
          cVar1S19S62N045P018P061N035(0) <='1';
          else
          cVar1S19S62N045P018P061N035(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='1' AND B( 2)='0' )then
          cVar1S20S62N045P018P061N035(0) <='1';
          else
          cVar1S20S62N045P018P061N035(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='0' AND B( 7)='1' )then
          cVar1S21S62N045P018N061P025(0) <='1';
          else
          cVar1S21S62N045P018N061P025(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='0' AND B( 7)='1' )then
          cVar1S22S62N045P018N061P025(0) <='1';
          else
          cVar1S22S62N045P018N061P025(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='0' AND B( 7)='0' )then
          cVar1S23S62N045P018N061N025(0) <='1';
          else
          cVar1S23S62N045P018N061N025(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND D(10)='0' AND B( 7)='0' )then
          cVar1S24S62N045P018N061N025(0) <='1';
          else
          cVar1S24S62N045P018N061N025(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='1' AND B( 1)='0' )then
          cVar1S0S63P045P005P037nsss(0) <='1';
          else
          cVar1S0S63P045P005P037nsss(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A( 6)='1' )then
          cVar1S1S63P045N005P021P007(0) <='1';
          else
          cVar1S1S63P045N005P021P007(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A( 6)='0' )then
          cVar1S2S63P045N005P021N007(0) <='1';
          else
          cVar1S2S63P045N005P021N007(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A( 6)='0' )then
          cVar1S3S63P045N005P021N007(0) <='1';
          else
          cVar1S3S63P045N005P021N007(0) <='0';
          end if;
        if(D(14)='1' AND A( 7)='0' AND B( 9)='0' AND A( 6)='0' )then
          cVar1S4S63P045N005P021N007(0) <='1';
          else
          cVar1S4S63P045N005P021N007(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S5S63N045P018P019P056(0) <='1';
          else
          cVar1S5S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S6S63N045P018P019P056(0) <='1';
          else
          cVar1S6S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S7S63N045P018P019P056(0) <='1';
          else
          cVar1S7S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='0' )then
          cVar1S8S63N045P018P019P056(0) <='1';
          else
          cVar1S8S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S9S63N045P018P019P056(0) <='1';
          else
          cVar1S9S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S10S63N045P018P019P056(0) <='1';
          else
          cVar1S10S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='1' AND D( 3)='1' )then
          cVar1S11S63N045P018P019P056(0) <='1';
          else
          cVar1S11S63N045P018P019P056(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S12S63N045P018N019P024(0) <='1';
          else
          cVar1S12S63N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S13S63N045P018N019P024(0) <='1';
          else
          cVar1S13S63N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S14S63N045P018N019P024(0) <='1';
          else
          cVar1S14S63N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='0' )then
          cVar1S15S63N045P018N019P024(0) <='1';
          else
          cVar1S15S63N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='1' AND A( 0)='0' AND B(17)='1' )then
          cVar1S16S63N045P018N019P024(0) <='1';
          else
          cVar1S16S63N045P018N019P024(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='1' AND B( 4)='0' )then
          cVar1S17S63N045N018P030P031(0) <='1';
          else
          cVar1S17S63N045N018P030P031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='1' AND B( 4)='0' )then
          cVar1S18S63N045N018P030P031(0) <='1';
          else
          cVar1S18S63N045N018P030P031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='1' )then
          cVar1S19S63N045N018N030P031(0) <='1';
          else
          cVar1S19S63N045N018N030P031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='1' )then
          cVar1S20S63N045N018N030P031(0) <='1';
          else
          cVar1S20S63N045N018N030P031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='1' )then
          cVar1S21S63N045N018N030P031(0) <='1';
          else
          cVar1S21S63N045N018N030P031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='0' )then
          cVar1S22S63N045N018N030N031(0) <='1';
          else
          cVar1S22S63N045N018N030N031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='0' )then
          cVar1S23S63N045N018N030N031(0) <='1';
          else
          cVar1S23S63N045N018N030N031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='0' )then
          cVar1S24S63N045N018N030N031(0) <='1';
          else
          cVar1S24S63N045N018N030N031(0) <='0';
          end if;
        if(D(14)='0' AND A(10)='0' AND B(14)='0' AND B( 4)='0' )then
          cVar1S25S63N045N018N030N031(0) <='1';
          else
          cVar1S25S63N045N018N030N031(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='1' )then
          cVar1S0S64P018P069P011P029(0) <='1';
          else
          cVar1S0S64P018P069P011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='1' )then
          cVar1S1S64P018P069P011P029(0) <='1';
          else
          cVar1S1S64P018P069P011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='1' )then
          cVar1S2S64P018P069P011P029(0) <='1';
          else
          cVar1S2S64P018P069P011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='0' )then
          cVar1S3S64P018P069P011N029(0) <='1';
          else
          cVar1S3S64P018P069P011N029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='0' )then
          cVar1S4S64P018P069P011N029(0) <='1';
          else
          cVar1S4S64P018P069P011N029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='1' AND B( 5)='0' )then
          cVar1S5S64P018P069P011N029(0) <='1';
          else
          cVar1S5S64P018P069P011N029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='0' )then
          cVar1S6S64P018P069N011P029(0) <='1';
          else
          cVar1S6S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='0' )then
          cVar1S7S64P018P069N011P029(0) <='1';
          else
          cVar1S7S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='0' )then
          cVar1S8S64P018P069N011P029(0) <='1';
          else
          cVar1S8S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='0' )then
          cVar1S9S64P018P069N011P029(0) <='1';
          else
          cVar1S9S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='1' )then
          cVar1S10S64P018P069N011P029(0) <='1';
          else
          cVar1S10S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='0' AND A( 4)='0' AND B( 5)='1' )then
          cVar1S11S64P018P069N011P029(0) <='1';
          else
          cVar1S11S64P018P069N011P029(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='1' AND E( 9)='1' )then
          cVar1S12S64P018P069P019P067(0) <='1';
          else
          cVar1S12S64P018P069P019P067(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='1' AND E( 9)='1' )then
          cVar1S13S64P018P069P019P067(0) <='1';
          else
          cVar1S13S64P018P069P019P067(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='1' AND E( 9)='1' )then
          cVar1S14S64P018P069P019P067(0) <='1';
          else
          cVar1S14S64P018P069P019P067(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='1' AND E( 9)='0' )then
          cVar1S15S64P018P069P019N067(0) <='1';
          else
          cVar1S15S64P018P069P019N067(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S16S64P018P069N019P068(0) <='1';
          else
          cVar1S16S64P018P069N019P068(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='0' AND D( 0)='1' )then
          cVar1S17S64P018P069N019P068(0) <='1';
          else
          cVar1S17S64P018P069N019P068(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='0' AND D( 0)='0' )then
          cVar1S18S64P018P069N019N068(0) <='1';
          else
          cVar1S18S64P018P069N019N068(0) <='0';
          end if;
        if(A(10)='0' AND D( 8)='1' AND A( 0)='0' AND D( 0)='0' )then
          cVar1S19S64P018P069N019N068(0) <='1';
          else
          cVar1S19S64P018P069N019N068(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='1' AND A( 6)='0' AND A( 3)='1' )then
          cVar1S20S64P018P031P007P013(0) <='1';
          else
          cVar1S20S64P018P031P007P013(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='1' AND A( 6)='0' AND A( 3)='1' )then
          cVar1S21S64P018P031P007P013(0) <='1';
          else
          cVar1S21S64P018P031P007P013(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='1' AND A( 6)='0' AND A( 3)='1' )then
          cVar1S22S64P018P031P007P013(0) <='1';
          else
          cVar1S22S64P018P031P007P013(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='1' AND A( 6)='0' AND A( 3)='0' )then
          cVar1S23S64P018P031P007N013(0) <='1';
          else
          cVar1S23S64P018P031P007N013(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='1' AND A( 6)='0' AND A( 3)='0' )then
          cVar1S24S64P018P031P007N013(0) <='1';
          else
          cVar1S24S64P018P031P007N013(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='1' AND E(13)='1' )then
          cVar1S25S64P018N031P007P051nsss(0) <='1';
          else
          cVar1S25S64P018N031P007P051nsss(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='1' AND E(13)='0' )then
          cVar1S26S64P018N031P007N051(0) <='1';
          else
          cVar1S26S64P018N031P007N051(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='1' AND E(13)='0' )then
          cVar1S27S64P018N031P007N051(0) <='1';
          else
          cVar1S27S64P018N031P007N051(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='1' AND E(13)='0' )then
          cVar1S28S64P018N031P007N051(0) <='1';
          else
          cVar1S28S64P018N031P007N051(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S29S64P018N031N007P009(0) <='1';
          else
          cVar1S29S64P018N031N007P009(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S30S64P018N031N007P009(0) <='1';
          else
          cVar1S30S64P018N031N007P009(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S31S64P018N031N007N009(0) <='1';
          else
          cVar1S31S64P018N031N007N009(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S32S64P018N031N007N009(0) <='1';
          else
          cVar1S32S64P018N031N007N009(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S33S64P018N031N007N009(0) <='1';
          else
          cVar1S33S64P018N031N007N009(0) <='0';
          end if;
        if(A(10)='1' AND B( 4)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S34S64P018N031N007N009(0) <='1';
          else
          cVar1S34S64P018N031N007N009(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='0' AND D( 0)='1' )then
          cVar1S0S65P018P014P042P068(0) <='1';
          else
          cVar1S0S65P018P014P042P068(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='0' AND D( 0)='1' )then
          cVar1S1S65P018P014P042P068(0) <='1';
          else
          cVar1S1S65P018P014P042P068(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='0' AND D( 0)='0' )then
          cVar1S2S65P018P014P042N068(0) <='1';
          else
          cVar1S2S65P018P014P042N068(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='0' AND D( 0)='0' )then
          cVar1S3S65P018P014P042N068(0) <='1';
          else
          cVar1S3S65P018P014P042N068(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='1' AND A(17)='1' )then
          cVar1S4S65P018P014P042P004nsss(0) <='1';
          else
          cVar1S4S65P018P014P042P004nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='1' AND A(17)='0' )then
          cVar1S5S65P018P014P042N004(0) <='1';
          else
          cVar1S5S65P018P014P042N004(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='0' AND E( 7)='1' AND A(17)='0' )then
          cVar1S6S65P018P014P042N004(0) <='1';
          else
          cVar1S6S65P018P014P042N004(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='1' )then
          cVar1S7S65P018P014P045nsss(0) <='1';
          else
          cVar1S7S65P018P014P045nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='0' AND E( 6)='1' )then
          cVar1S8S65P018P014N045P046nsss(0) <='1';
          else
          cVar1S8S65P018P014N045P046nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='0' AND E( 6)='0' )then
          cVar1S9S65P018P014N045N046(0) <='1';
          else
          cVar1S9S65P018P014N045N046(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='0' AND E( 6)='0' )then
          cVar1S10S65P018P014N045N046(0) <='1';
          else
          cVar1S10S65P018P014N045N046(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='0' AND E( 6)='0' )then
          cVar1S11S65P018P014N045N046(0) <='1';
          else
          cVar1S11S65P018P014N045N046(0) <='0';
          end if;
        if(A(10)='1' AND A(12)='1' AND D(14)='0' AND E( 6)='0' )then
          cVar1S12S65P018P014N045N046(0) <='1';
          else
          cVar1S12S65P018P014N045N046(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='1' )then
          cVar1S13S65N018P041P020P002nsss(0) <='1';
          else
          cVar1S13S65N018P041P020P002nsss(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='0' )then
          cVar1S14S65N018P041P020N002(0) <='1';
          else
          cVar1S14S65N018P041P020N002(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='0' )then
          cVar1S15S65N018P041P020N002(0) <='1';
          else
          cVar1S15S65N018P041P020N002(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='1' )then
          cVar1S16S65N018P041N020P023(0) <='1';
          else
          cVar1S16S65N018P041N020P023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='0' )then
          cVar1S17S65N018P041N020N023(0) <='1';
          else
          cVar1S17S65N018P041N020N023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='0' )then
          cVar1S18S65N018P041N020N023(0) <='1';
          else
          cVar1S18S65N018P041N020N023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S19S65N018N041P039P045(0) <='1';
          else
          cVar1S19S65N018N041P039P045(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S20S65N018N041P039P045(0) <='1';
          else
          cVar1S20S65N018N041P039P045(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S21S65N018N041P039N045(0) <='1';
          else
          cVar1S21S65N018N041P039N045(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S22S65N018N041P039N045(0) <='1';
          else
          cVar1S22S65N018N041P039N045(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S23S65N018N041P039N045(0) <='1';
          else
          cVar1S23S65N018N041P039N045(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='1' )then
          cVar1S24S65N018N041P039P049nsss(0) <='1';
          else
          cVar1S24S65N018N041P039P049nsss(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='1' AND D(13)='0' )then
          cVar1S25S65N018N041P039N049(0) <='1';
          else
          cVar1S25S65N018N041P039N049(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='1' )then
          cVar1S0S66P018P041P020P002nsss(0) <='1';
          else
          cVar1S0S66P018P041P020P002nsss(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='0' )then
          cVar1S1S66P018P041P020N002(0) <='1';
          else
          cVar1S1S66P018P041P020N002(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='1' AND A(18)='0' )then
          cVar1S2S66P018P041P020N002(0) <='1';
          else
          cVar1S2S66P018P041P020N002(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='1' )then
          cVar1S3S66P018P041N020P023(0) <='1';
          else
          cVar1S3S66P018P041N020P023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='0' )then
          cVar1S4S66P018P041N020N023(0) <='1';
          else
          cVar1S4S66P018P041N020N023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='1' AND B(19)='0' AND B( 8)='0' )then
          cVar1S5S66P018P041N020N023(0) <='1';
          else
          cVar1S5S66P018P041N020N023(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='0' )then
          cVar1S6S66P018N041P039P020(0) <='1';
          else
          cVar1S6S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='0' )then
          cVar1S7S66P018N041P039P020(0) <='1';
          else
          cVar1S7S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='0' )then
          cVar1S8S66P018N041P039P020(0) <='1';
          else
          cVar1S8S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='0' )then
          cVar1S9S66P018N041P039P020(0) <='1';
          else
          cVar1S9S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='1' )then
          cVar1S10S66P018N041P039P020(0) <='1';
          else
          cVar1S10S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='1' )then
          cVar1S11S66P018N041P039P020(0) <='1';
          else
          cVar1S11S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='0' AND B(19)='1' )then
          cVar1S12S66P018N041P039P020(0) <='1';
          else
          cVar1S12S66P018N041P039P020(0) <='0';
          end if;
        if(A(10)='0' AND D(15)='0' AND B( 0)='1' AND A( 4)='0' )then
          cVar1S13S66P018N041P039P011(0) <='1';
          else
          cVar1S13S66P018N041P039P011(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='1' )then
          cVar1S14S66P018P068P057nsss(0) <='1';
          else
          cVar1S14S66P018P068P057nsss(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='0' AND E(10)='0' )then
          cVar1S15S66P018P068N057P063(0) <='1';
          else
          cVar1S15S66P018P068N057P063(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='0' AND E(10)='0' )then
          cVar1S16S66P018P068N057P063(0) <='1';
          else
          cVar1S16S66P018P068N057P063(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='0' AND E(10)='1' )then
          cVar1S17S66P018P068N057P063(0) <='1';
          else
          cVar1S17S66P018P068N057P063(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='0' AND E(10)='1' )then
          cVar1S18S66P018P068N057P063(0) <='1';
          else
          cVar1S18S66P018P068N057P063(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='1' AND D(11)='0' AND E(10)='1' )then
          cVar1S19S66P018P068N057P063(0) <='1';
          else
          cVar1S19S66P018P068N057P063(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S20S66P018N068P031P013(0) <='1';
          else
          cVar1S20S66P018N068P031P013(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S21S66P018N068P031N013(0) <='1';
          else
          cVar1S21S66P018N068P031N013(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S22S66P018N068P031N013(0) <='1';
          else
          cVar1S22S66P018N068P031N013(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='0' AND A( 7)='1' )then
          cVar1S23S66P018N068N031P005(0) <='1';
          else
          cVar1S23S66P018N068N031P005(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='0' AND A( 7)='0' )then
          cVar1S24S66P018N068N031N005(0) <='1';
          else
          cVar1S24S66P018N068N031N005(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='0' AND A( 7)='0' )then
          cVar1S25S66P018N068N031N005(0) <='1';
          else
          cVar1S25S66P018N068N031N005(0) <='0';
          end if;
        if(A(10)='1' AND D( 0)='0' AND B( 4)='0' AND A( 7)='0' )then
          cVar1S26S66P018N068N031N005(0) <='1';
          else
          cVar1S26S66P018N068N031N005(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='1' AND E(10)='0' AND A(10)='0' )then
          cVar1S0S67P009P027P063P018nsss(0) <='1';
          else
          cVar1S0S67P009P027P063P018nsss(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='1' AND E(10)='0' AND A(10)='1' )then
          cVar1S1S67P009P027P063P018(0) <='1';
          else
          cVar1S1S67P009P027P063P018(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='1' AND E(10)='0' AND A(10)='1' )then
          cVar1S2S67P009P027P063P018(0) <='1';
          else
          cVar1S2S67P009P027P063P018(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S3S67P009N027P049P026nsss(0) <='1';
          else
          cVar1S3S67P009N027P049P026nsss(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S4S67P009N027P049N026(0) <='1';
          else
          cVar1S4S67P009N027P049N026(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S5S67P009N027P049N026(0) <='1';
          else
          cVar1S5S67P009N027P049N026(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND A(12)='1' )then
          cVar1S6S67P009N027N049P014(0) <='1';
          else
          cVar1S6S67P009N027N049P014(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND A(12)='1' )then
          cVar1S7S67P009N027N049P014(0) <='1';
          else
          cVar1S7S67P009N027N049P014(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND A(12)='0' )then
          cVar1S8S67P009N027N049N014(0) <='1';
          else
          cVar1S8S67P009N027N049N014(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND A(12)='0' )then
          cVar1S9S67P009N027N049N014(0) <='1';
          else
          cVar1S9S67P009N027N049N014(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND A(12)='0' )then
          cVar1S10S67P009N027N049N014(0) <='1';
          else
          cVar1S10S67P009N027N049N014(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND B( 0)='1' )then
          cVar1S11S67N009P041P020P039nsss(0) <='1';
          else
          cVar1S11S67N009P041P020P039nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='1' )then
          cVar1S12S67N009P041N020P021nsss(0) <='1';
          else
          cVar1S12S67N009P041N020P021nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S13S67N009P041N020N021(0) <='1';
          else
          cVar1S13S67N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S14S67N009P041N020N021(0) <='1';
          else
          cVar1S14S67N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S15S67N009P041N020N021(0) <='1';
          else
          cVar1S15S67N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='1' )then
          cVar1S16S67N009N041P018P000(0) <='1';
          else
          cVar1S16S67N009N041P018P000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='1' )then
          cVar1S17S67N009N041P018P000(0) <='1';
          else
          cVar1S17S67N009N041P018P000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='0' )then
          cVar1S18S67N009N041P018N000(0) <='1';
          else
          cVar1S18S67N009N041P018N000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='0' )then
          cVar1S19S67N009N041P018N000(0) <='1';
          else
          cVar1S19S67N009N041P018N000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='0' )then
          cVar1S20S67N009N041P018N000(0) <='1';
          else
          cVar1S20S67N009N041P018N000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='1' AND A(19)='0' )then
          cVar1S21S67N009N041P018N000(0) <='1';
          else
          cVar1S21S67N009N041P018N000(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='0' AND B( 0)='0' )then
          cVar1S22S67N009N041N018P039(0) <='1';
          else
          cVar1S22S67N009N041N018P039(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='0' AND B( 0)='0' )then
          cVar1S23S67N009N041N018P039(0) <='1';
          else
          cVar1S23S67N009N041N018P039(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='0' AND B( 0)='0' )then
          cVar1S24S67N009N041N018P039(0) <='1';
          else
          cVar1S24S67N009N041N018P039(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='0' AND B( 0)='0' )then
          cVar1S25S67N009N041N018P039(0) <='1';
          else
          cVar1S25S67N009N041N018P039(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(10)='0' AND B( 0)='1' )then
          cVar1S26S67N009N041N018P039(0) <='1';
          else
          cVar1S26S67N009N041N018P039(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='1' AND E(10)='0' AND A(10)='0' )then
          cVar1S0S68P009P027P063P018nsss(0) <='1';
          else
          cVar1S0S68P009P027P063P018nsss(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='1' AND E(10)='0' AND A(10)='1' )then
          cVar1S1S68P009P027P063P018(0) <='1';
          else
          cVar1S1S68P009P027P063P018(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S2S68P009N027P049P026nsss(0) <='1';
          else
          cVar1S2S68P009N027P049P026nsss(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S3S68P009N027P049N026(0) <='1';
          else
          cVar1S3S68P009N027P049N026(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S4S68P009N027P049N026(0) <='1';
          else
          cVar1S4S68P009N027P049N026(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='1' )then
          cVar1S5S68P009N027N049P053(0) <='1';
          else
          cVar1S5S68P009N027N049P053(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='1' )then
          cVar1S6S68P009N027N049P053(0) <='1';
          else
          cVar1S6S68P009N027N049P053(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='0' )then
          cVar1S7S68P009N027N049N053(0) <='1';
          else
          cVar1S7S68P009N027N049N053(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='0' )then
          cVar1S8S68P009N027N049N053(0) <='1';
          else
          cVar1S8S68P009N027N049N053(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='0' )then
          cVar1S9S68P009N027N049N053(0) <='1';
          else
          cVar1S9S68P009N027N049N053(0) <='0';
          end if;
        if(A( 5)='1' AND B( 6)='0' AND D(13)='0' AND D(12)='0' )then
          cVar1S10S68P009N027N049N053(0) <='1';
          else
          cVar1S10S68P009N027N049N053(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S11S68N009P041P020P003nsss(0) <='1';
          else
          cVar1S11S68N009P041P020P003nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S12S68N009P041P020N003(0) <='1';
          else
          cVar1S12S68N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S13S68N009P041P020N003(0) <='1';
          else
          cVar1S13S68N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S14S68N009P041P020N003(0) <='1';
          else
          cVar1S14S68N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='1' )then
          cVar1S15S68N009P041N020P021(0) <='1';
          else
          cVar1S15S68N009P041N020P021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='1' )then
          cVar1S16S68N009P041N020P021(0) <='1';
          else
          cVar1S16S68N009P041N020P021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S17S68N009P041N020N021(0) <='1';
          else
          cVar1S17S68N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S18S68N009P041N020N021(0) <='1';
          else
          cVar1S18S68N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND B( 9)='0' )then
          cVar1S19S68N009P041N020N021(0) <='1';
          else
          cVar1S19S68N009P041N020N021(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='1' )then
          cVar1S20S68N009N041P016P031(0) <='1';
          else
          cVar1S20S68N009N041P016P031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='1' )then
          cVar1S21S68N009N041P016P031(0) <='1';
          else
          cVar1S21S68N009N041P016P031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='1' )then
          cVar1S22S68N009N041P016P031(0) <='1';
          else
          cVar1S22S68N009N041P016P031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='1' )then
          cVar1S23S68N009N041P016P031(0) <='1';
          else
          cVar1S23S68N009N041P016P031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='0' )then
          cVar1S24S68N009N041P016N031(0) <='1';
          else
          cVar1S24S68N009N041P016N031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='0' )then
          cVar1S25S68N009N041P016N031(0) <='1';
          else
          cVar1S25S68N009N041P016N031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='0' AND B( 4)='0' )then
          cVar1S26S68N009N041P016N031(0) <='1';
          else
          cVar1S26S68N009N041P016N031(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='1' AND E(11)='0' )then
          cVar1S27S68N009N041P016P059(0) <='1';
          else
          cVar1S27S68N009N041P016P059(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='1' AND E(11)='0' )then
          cVar1S28S68N009N041P016P059(0) <='1';
          else
          cVar1S28S68N009N041P016P059(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='1' AND E(11)='1' )then
          cVar1S29S68N009N041P016P059(0) <='1';
          else
          cVar1S29S68N009N041P016P059(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='1' AND E(11)='1' )then
          cVar1S30S68N009N041P016P059(0) <='1';
          else
          cVar1S30S68N009N041P016P059(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND A(11)='1' AND E(11)='1' )then
          cVar1S31S68N009N041P016P059(0) <='1';
          else
          cVar1S31S68N009N041P016P059(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND D( 2)='0' AND E( 9)='0' )then
          cVar1S0S69P009P049P060P067(0) <='1';
          else
          cVar1S0S69P009P049P060P067(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND D( 2)='0' AND E( 9)='0' )then
          cVar1S1S69P009P049P060P067(0) <='1';
          else
          cVar1S1S69P009P049P060P067(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND D( 2)='0' AND E( 9)='0' )then
          cVar1S2S69P009P049P060P067(0) <='1';
          else
          cVar1S2S69P009P049P060P067(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='1' AND B( 5)='1' )then
          cVar1S3S69P009N049P053P029nsss(0) <='1';
          else
          cVar1S3S69P009N049P053P029nsss(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S4S69P009N049P053N029(0) <='1';
          else
          cVar1S4S69P009N049P053N029(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S5S69P009N049P053N029(0) <='1';
          else
          cVar1S5S69P009N049P053N029(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S6S69P009N049N053P050(0) <='1';
          else
          cVar1S6S69P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S7S69P009N049N053P050(0) <='1';
          else
          cVar1S7S69P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S8S69P009N049N053P050(0) <='1';
          else
          cVar1S8S69P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S9S69P009N049N053N050(0) <='1';
          else
          cVar1S9S69P009N049N053N050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S10S69P009N049N053N050(0) <='1';
          else
          cVar1S10S69P009N049N053N050(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S11S69N009P041P020P003nsss(0) <='1';
          else
          cVar1S11S69N009P041P020P003nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S12S69N009P041P020N003(0) <='1';
          else
          cVar1S12S69N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S13S69N009P041P020N003(0) <='1';
          else
          cVar1S13S69N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S14S69N009P041P020N003(0) <='1';
          else
          cVar1S14S69N009P041P020N003(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='1' )then
          cVar1S15S69N009P041N020P001nsss(0) <='1';
          else
          cVar1S15S69N009P041N020P001nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S16S69N009P041N020N001(0) <='1';
          else
          cVar1S16S69N009P041N020N001(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S17S69N009P041N020N001(0) <='1';
          else
          cVar1S17S69N009P041N020N001(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S18S69N009P041N020N001(0) <='1';
          else
          cVar1S18S69N009P041N020N001(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S19S69N009N041P031P013(0) <='1';
          else
          cVar1S19S69N009N041P031P013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S20S69N009N041P031P013(0) <='1';
          else
          cVar1S20S69N009N041P031P013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S21S69N009N041P031P013(0) <='1';
          else
          cVar1S21S69N009N041P031P013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S22S69N009N041P031P013(0) <='1';
          else
          cVar1S22S69N009N041P031P013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S23S69N009N041P031N013(0) <='1';
          else
          cVar1S23S69N009N041P031N013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S24S69N009N041P031N013(0) <='1';
          else
          cVar1S24S69N009N041P031N013(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='0' )then
          cVar1S25S69N009N041N031P054(0) <='1';
          else
          cVar1S25S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='0' )then
          cVar1S26S69N009N041N031P054(0) <='1';
          else
          cVar1S26S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='0' )then
          cVar1S27S69N009N041N031P054(0) <='1';
          else
          cVar1S27S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='1' )then
          cVar1S28S69N009N041N031P054(0) <='1';
          else
          cVar1S28S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='1' )then
          cVar1S29S69N009N041N031P054(0) <='1';
          else
          cVar1S29S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='1' )then
          cVar1S30S69N009N041N031P054(0) <='1';
          else
          cVar1S30S69N009N041N031P054(0) <='0';
          end if;
        if(A( 5)='0' AND D(15)='0' AND B( 4)='0' AND E( 4)='1' )then
          cVar1S31S69N009N041N031P054(0) <='1';
          else
          cVar1S31S69N009N041N031P054(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S0S70P016P018P036P053(0) <='1';
          else
          cVar1S0S70P016P018P036P053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S1S70P016P018P036P053(0) <='1';
          else
          cVar1S1S70P016P018P036P053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='1' )then
          cVar1S2S70P016P018P036P053(0) <='1';
          else
          cVar1S2S70P016P018P036P053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S3S70P016P018P036N053(0) <='1';
          else
          cVar1S3S70P016P018P036N053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S4S70P016P018P036N053(0) <='1';
          else
          cVar1S4S70P016P018P036N053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S5S70P016P018P036N053(0) <='1';
          else
          cVar1S5S70P016P018P036N053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='0' AND D(12)='0' )then
          cVar1S6S70P016P018P036N053(0) <='1';
          else
          cVar1S6S70P016P018P036N053(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='1' AND A( 1)='1' )then
          cVar1S7S70P016P018P036P017(0) <='1';
          else
          cVar1S7S70P016P018P036P017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='1' AND A( 1)='1' )then
          cVar1S8S70P016P018P036P017(0) <='1';
          else
          cVar1S8S70P016P018P036P017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='1' AND A( 1)='0' )then
          cVar1S9S70P016P018P036N017(0) <='1';
          else
          cVar1S9S70P016P018P036N017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='1' AND A( 1)='0' )then
          cVar1S10S70P016P018P036N017(0) <='1';
          else
          cVar1S10S70P016P018P036N017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(11)='1' AND A( 1)='0' )then
          cVar1S11S70P016P018P036N017(0) <='1';
          else
          cVar1S11S70P016P018P036N017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='1' AND A( 1)='0' )then
          cVar1S12S70P016P018P045P017(0) <='1';
          else
          cVar1S12S70P016P018P045P017(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND B(16)='0' )then
          cVar1S13S70P016P018N045P026(0) <='1';
          else
          cVar1S13S70P016P018N045P026(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND B(16)='0' )then
          cVar1S14S70P016P018N045P026(0) <='1';
          else
          cVar1S14S70P016P018N045P026(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND B(16)='0' )then
          cVar1S15S70P016P018N045P026(0) <='1';
          else
          cVar1S15S70P016P018N045P026(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND B(16)='1' )then
          cVar1S16S70P016P018N045P026(0) <='1';
          else
          cVar1S16S70P016P018N045P026(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND B(16)='1' )then
          cVar1S17S70P016P018N045P026(0) <='1';
          else
          cVar1S17S70P016P018N045P026(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='0' AND D(15)='1' )then
          cVar1S18S70P016P035P053P041(0) <='1';
          else
          cVar1S18S70P016P035P053P041(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='0' AND D(15)='1' )then
          cVar1S19S70P016P035P053P041(0) <='1';
          else
          cVar1S19S70P016P035P053P041(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='0' AND D(15)='0' )then
          cVar1S20S70P016P035P053N041(0) <='1';
          else
          cVar1S20S70P016P035P053N041(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='0' AND D(15)='0' )then
          cVar1S21S70P016P035P053N041(0) <='1';
          else
          cVar1S21S70P016P035P053N041(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='0' AND D(15)='0' )then
          cVar1S22S70P016P035P053N041(0) <='1';
          else
          cVar1S22S70P016P035P053N041(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='1' AND B( 1)='1' )then
          cVar1S23S70P016P035P053P037(0) <='1';
          else
          cVar1S23S70P016P035P053P037(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='1' AND B( 1)='0' )then
          cVar1S24S70P016P035P053N037(0) <='1';
          else
          cVar1S24S70P016P035P053N037(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='0' AND D(12)='1' AND B( 1)='0' )then
          cVar1S25S70P016P035P053N037(0) <='1';
          else
          cVar1S25S70P016P035P053N037(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='1' AND B(13)='1' AND A(10)='1' )then
          cVar1S26S70P016P035P032P018nsss(0) <='1';
          else
          cVar1S26S70P016P035P032P018nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 2)='1' AND B(13)='0' AND B(12)='0' )then
          cVar1S27S70P016P035N032P034(0) <='1';
          else
          cVar1S27S70P016P035N032P034(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S0S71P041P020P003nsss(0) <='1';
          else
          cVar1S0S71P041P020P003nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='1' )then
          cVar1S1S71P041P020N003P002nsss(0) <='1';
          else
          cVar1S1S71P041P020N003P002nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='0' )then
          cVar1S2S71P041P020N003N002(0) <='1';
          else
          cVar1S2S71P041P020N003N002(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='1' AND A( 8)='0' AND A(18)='0' )then
          cVar1S3S71P041P020N003N002(0) <='1';
          else
          cVar1S3S71P041P020N003N002(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='1' )then
          cVar1S4S71P041N020P001nsss(0) <='1';
          else
          cVar1S4S71P041N020P001nsss(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='1' )then
          cVar1S5S71P041N020N001P005(0) <='1';
          else
          cVar1S5S71P041N020N001P005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='1' )then
          cVar1S6S71P041N020N001P005(0) <='1';
          else
          cVar1S6S71P041N020N001P005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='1' )then
          cVar1S7S71P041N020N001P005(0) <='1';
          else
          cVar1S7S71P041N020N001P005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='0' )then
          cVar1S8S71P041N020N001N005(0) <='1';
          else
          cVar1S8S71P041N020N001N005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='0' )then
          cVar1S9S71P041N020N001N005(0) <='1';
          else
          cVar1S9S71P041N020N001N005(0) <='0';
          end if;
        if(D(15)='1' AND B(19)='0' AND A( 9)='0' AND A( 7)='0' )then
          cVar1S10S71P041N020N001N005(0) <='1';
          else
          cVar1S10S71P041N020N001N005(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='1' AND B( 3)='0' )then
          cVar1S11S71N041P049P026P033(0) <='1';
          else
          cVar1S11S71N041P049P026P033(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S12S71N041P049N026P024(0) <='1';
          else
          cVar1S12S71N041P049N026P024(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S13S71N041P049N026P024(0) <='1';
          else
          cVar1S13S71N041P049N026P024(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='0' AND B(17)='0' )then
          cVar1S14S71N041P049N026N024(0) <='1';
          else
          cVar1S14S71N041P049N026N024(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='0' AND B(17)='0' )then
          cVar1S15S71N041P049N026N024(0) <='1';
          else
          cVar1S15S71N041P049N026N024(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='1' AND B(16)='0' AND B(17)='0' )then
          cVar1S16S71N041P049N026N024(0) <='1';
          else
          cVar1S16S71N041P049N026N024(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S17S71N041N049P039P045(0) <='1';
          else
          cVar1S17S71N041N049P039P045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S18S71N041N049P039P045(0) <='1';
          else
          cVar1S18S71N041N049P039P045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S19S71N041N049P039P045(0) <='1';
          else
          cVar1S19S71N041N049P039P045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S20S71N041N049P039N045(0) <='1';
          else
          cVar1S20S71N041N049P039N045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S21S71N041N049P039N045(0) <='1';
          else
          cVar1S21S71N041N049P039N045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S22S71N041N049P039N045(0) <='1';
          else
          cVar1S22S71N041N049P039N045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S23S71N041N049P039N045(0) <='1';
          else
          cVar1S23S71N041N049P039N045(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='1' AND B(11)='1' )then
          cVar1S24S71N041N049P039P036nsss(0) <='1';
          else
          cVar1S24S71N041N049P039P036nsss(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='1' AND B(11)='0' )then
          cVar1S25S71N041N049P039N036(0) <='1';
          else
          cVar1S25S71N041N049P039N036(0) <='0';
          end if;
        if(D(15)='0' AND D(13)='0' AND B( 0)='1' AND B(11)='0' )then
          cVar1S26S71N041N049P039N036(0) <='1';
          else
          cVar1S26S71N041N049P039N036(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='1' AND E( 7)='1' )then
          cVar1S0S72P016P018P023P042nsss(0) <='1';
          else
          cVar1S0S72P016P018P023P042nsss(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='1' AND E( 7)='0' )then
          cVar1S1S72P016P018P023N042(0) <='1';
          else
          cVar1S1S72P016P018P023N042(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='1' AND E( 7)='0' )then
          cVar1S2S72P016P018P023N042(0) <='1';
          else
          cVar1S2S72P016P018P023N042(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='1' )then
          cVar1S3S72P016P018N023P047(0) <='1';
          else
          cVar1S3S72P016P018N023P047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='1' )then
          cVar1S4S72P016P018N023P047(0) <='1';
          else
          cVar1S4S72P016P018N023P047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='1' )then
          cVar1S5S72P016P018N023P047(0) <='1';
          else
          cVar1S5S72P016P018N023P047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='0' )then
          cVar1S6S72P016P018N023N047(0) <='1';
          else
          cVar1S6S72P016P018N023N047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='0' )then
          cVar1S7S72P016P018N023N047(0) <='1';
          else
          cVar1S7S72P016P018N023N047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B( 8)='0' AND E(14)='0' )then
          cVar1S8S72P016P018N023N047(0) <='1';
          else
          cVar1S8S72P016P018N023N047(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='1' AND A( 2)='1' )then
          cVar1S9S72P016P018P045P015nsss(0) <='1';
          else
          cVar1S9S72P016P018P045P015nsss(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='1' AND A( 2)='0' )then
          cVar1S10S72P016P018P045N015(0) <='1';
          else
          cVar1S10S72P016P018P045N015(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='0' )then
          cVar1S11S72P016P018N045P013(0) <='1';
          else
          cVar1S11S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='0' )then
          cVar1S12S72P016P018N045P013(0) <='1';
          else
          cVar1S12S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='0' )then
          cVar1S13S72P016P018N045P013(0) <='1';
          else
          cVar1S13S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='0' )then
          cVar1S14S72P016P018N045P013(0) <='1';
          else
          cVar1S14S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='1' )then
          cVar1S15S72P016P018N045P013(0) <='1';
          else
          cVar1S15S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='1' )then
          cVar1S16S72P016P018N045P013(0) <='1';
          else
          cVar1S16S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(14)='0' AND A( 3)='1' )then
          cVar1S17S72P016P018N045P013(0) <='1';
          else
          cVar1S17S72P016P018N045P013(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='1' AND A( 4)='0' )then
          cVar1S18S72P016P033P041P011(0) <='1';
          else
          cVar1S18S72P016P033P041P011(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='1' AND A( 4)='0' )then
          cVar1S19S72P016P033P041P011(0) <='1';
          else
          cVar1S19S72P016P033P041P011(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='0' AND A( 5)='1' )then
          cVar1S20S72P016P033N041P009(0) <='1';
          else
          cVar1S20S72P016P033N041P009(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='0' AND A( 5)='1' )then
          cVar1S21S72P016P033N041P009(0) <='1';
          else
          cVar1S21S72P016P033N041P009(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='0' AND A( 5)='1' )then
          cVar1S22S72P016P033N041P009(0) <='1';
          else
          cVar1S22S72P016P033N041P009(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='0' AND A( 5)='0' )then
          cVar1S23S72P016P033N041N009(0) <='1';
          else
          cVar1S23S72P016P033N041N009(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='0' AND D(15)='0' AND A( 5)='0' )then
          cVar1S24S72P016P033N041N009(0) <='1';
          else
          cVar1S24S72P016P033N041N009(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='0' AND D( 0)='1' )then
          cVar1S25S72P016P033P069P068(0) <='1';
          else
          cVar1S25S72P016P033P069P068(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='0' AND D( 0)='1' )then
          cVar1S26S72P016P033P069P068(0) <='1';
          else
          cVar1S26S72P016P033P069P068(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='0' AND D( 0)='0' )then
          cVar1S27S72P016P033P069N068(0) <='1';
          else
          cVar1S27S72P016P033P069N068(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='0' AND D( 0)='0' )then
          cVar1S28S72P016P033P069N068(0) <='1';
          else
          cVar1S28S72P016P033P069N068(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='0' AND D( 0)='0' )then
          cVar1S29S72P016P033P069N068(0) <='1';
          else
          cVar1S29S72P016P033P069N068(0) <='0';
          end if;
        if(A(11)='1' AND B( 3)='1' AND D( 8)='1' AND E( 9)='1' )then
          cVar1S30S72P016P033P069P067(0) <='1';
          else
          cVar1S30S72P016P033P069P067(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='1' AND B(17)='1' )then
          cVar1S0S73P047P006P024nsss(0) <='1';
          else
          cVar1S0S73P047P006P024nsss(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S73P047P006N024P026nsss(0) <='1';
          else
          cVar1S1S73P047P006N024P026nsss(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='1' AND B(16)='1' )then
          cVar1S2S73P047N006P008P026nsss(0) <='1';
          else
          cVar1S2S73P047N006P008P026nsss(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='1' AND B(16)='0' )then
          cVar1S3S73P047N006P008N026(0) <='1';
          else
          cVar1S3S73P047N006P008N026(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='0' AND A( 6)='1' )then
          cVar1S4S73P047N006N008P007(0) <='1';
          else
          cVar1S4S73P047N006N008P007(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='0' AND A( 6)='0' )then
          cVar1S5S73P047N006N008N007(0) <='1';
          else
          cVar1S5S73P047N006N008N007(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='0' AND A( 6)='0' )then
          cVar1S6S73P047N006N008N007(0) <='1';
          else
          cVar1S6S73P047N006N008N007(0) <='0';
          end if;
        if(E(14)='1' AND A(16)='0' AND A(15)='0' AND A( 6)='0' )then
          cVar1S7S73P047N006N008N007(0) <='1';
          else
          cVar1S7S73P047N006N008N007(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='1' AND D( 3)='1' )then
          cVar1S8S73N047P031P013P056(0) <='1';
          else
          cVar1S8S73N047P031P013P056(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='1' AND D( 3)='1' )then
          cVar1S9S73N047P031P013P056(0) <='1';
          else
          cVar1S9S73N047P031P013P056(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='1' AND D( 3)='0' )then
          cVar1S10S73N047P031P013N056(0) <='1';
          else
          cVar1S10S73N047P031P013N056(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='1' AND D( 3)='0' )then
          cVar1S11S73N047P031P013N056(0) <='1';
          else
          cVar1S11S73N047P031P013N056(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='1' AND D( 3)='0' )then
          cVar1S12S73N047P031P013N056(0) <='1';
          else
          cVar1S12S73N047P031P013N056(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar1S13S73N047P031N013P011(0) <='1';
          else
          cVar1S13S73N047P031N013P011(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar1S14S73N047P031N013P011(0) <='1';
          else
          cVar1S14S73N047P031N013P011(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='0' AND A( 4)='0' )then
          cVar1S15S73N047P031N013N011(0) <='1';
          else
          cVar1S15S73N047P031N013N011(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='1' AND A( 3)='0' AND A( 4)='0' )then
          cVar1S16S73N047P031N013N011(0) <='1';
          else
          cVar1S16S73N047P031N013N011(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='1' )then
          cVar1S17S73N047N031P030P012(0) <='1';
          else
          cVar1S17S73N047N031P030P012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='1' )then
          cVar1S18S73N047N031P030P012(0) <='1';
          else
          cVar1S18S73N047N031P030P012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='1' )then
          cVar1S19S73N047N031P030P012(0) <='1';
          else
          cVar1S19S73N047N031P030P012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='0' )then
          cVar1S20S73N047N031P030N012(0) <='1';
          else
          cVar1S20S73N047N031P030N012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='0' )then
          cVar1S21S73N047N031P030N012(0) <='1';
          else
          cVar1S21S73N047N031P030N012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='1' AND A(13)='0' )then
          cVar1S22S73N047N031P030N012(0) <='1';
          else
          cVar1S22S73N047N031P030N012(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S23S73N047N031N030P057(0) <='1';
          else
          cVar1S23S73N047N031N030P057(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S24S73N047N031N030P057(0) <='1';
          else
          cVar1S24S73N047N031N030P057(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S25S73N047N031N030P057(0) <='1';
          else
          cVar1S25S73N047N031N030P057(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S26S73N047N031N030P057(0) <='1';
          else
          cVar1S26S73N047N031N030P057(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S27S73N047N031N030P057(0) <='1';
          else
          cVar1S27S73N047N031N030P057(0) <='0';
          end if;
        if(E(14)='0' AND B( 4)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S28S73N047N031N030P057(0) <='1';
          else
          cVar1S28S73N047N031N030P057(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='1' )then
          cVar1S0S74P064P066P027P009(0) <='1';
          else
          cVar1S0S74P064P066P027P009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='1' )then
          cVar1S1S74P064P066P027P009(0) <='1';
          else
          cVar1S1S74P064P066P027P009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='1' )then
          cVar1S2S74P064P066P027P009(0) <='1';
          else
          cVar1S2S74P064P066P027P009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='1' )then
          cVar1S3S74P064P066P027P009(0) <='1';
          else
          cVar1S3S74P064P066P027P009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S4S74P064P066P027N009(0) <='1';
          else
          cVar1S4S74P064P066P027N009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S5S74P064P066P027N009(0) <='1';
          else
          cVar1S5S74P064P066P027N009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='1' AND A( 5)='0' )then
          cVar1S6S74P064P066P027N009(0) <='1';
          else
          cVar1S6S74P064P066P027N009(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='1' )then
          cVar1S7S74P064P066N027P041(0) <='1';
          else
          cVar1S7S74P064P066N027P041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='1' )then
          cVar1S8S74P064P066N027P041(0) <='1';
          else
          cVar1S8S74P064P066N027P041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='1' )then
          cVar1S9S74P064P066N027P041(0) <='1';
          else
          cVar1S9S74P064P066N027P041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='1' )then
          cVar1S10S74P064P066N027P041(0) <='1';
          else
          cVar1S10S74P064P066N027P041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='0' )then
          cVar1S11S74P064P066N027N041(0) <='1';
          else
          cVar1S11S74P064P066N027N041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='0' )then
          cVar1S12S74P064P066N027N041(0) <='1';
          else
          cVar1S12S74P064P066N027N041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='0' )then
          cVar1S13S74P064P066N027N041(0) <='1';
          else
          cVar1S13S74P064P066N027N041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='0' AND B( 6)='0' AND D(15)='0' )then
          cVar1S14S74P064P066N027N041(0) <='1';
          else
          cVar1S14S74P064P066N027N041(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='1' AND A(16)='0' AND E(11)='0' )then
          cVar1S15S74P064P066P006P059(0) <='1';
          else
          cVar1S15S74P064P066P006P059(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='1' AND A(16)='0' AND E(11)='0' )then
          cVar1S16S74P064P066P006P059(0) <='1';
          else
          cVar1S16S74P064P066P006P059(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='1' AND A(16)='0' AND E(11)='1' )then
          cVar1S17S74P064P066P006P059(0) <='1';
          else
          cVar1S17S74P064P066P006P059(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='1' AND A(16)='1' AND B( 2)='0' )then
          cVar1S18S74P064P066P006P035(0) <='1';
          else
          cVar1S18S74P064P066P006P035(0) <='0';
          end if;
        if(D( 1)='0' AND E( 1)='1' AND A(16)='1' AND B( 2)='0' )then
          cVar1S19S74P064P066P006P035(0) <='1';
          else
          cVar1S19S74P064P066P006P035(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='0' AND E( 7)='1' AND A( 1)='0' )then
          cVar1S20S74P064P011P042P017nsss(0) <='1';
          else
          cVar1S20S74P064P011P042P017nsss(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='0' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S21S74P064P011N042P003(0) <='1';
          else
          cVar1S21S74P064P011N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='0' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S22S74P064P011N042P003(0) <='1';
          else
          cVar1S22S74P064P011N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='0' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S23S74P064P011N042P003(0) <='1';
          else
          cVar1S23S74P064P011N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='0' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S24S74P064P011N042P003(0) <='1';
          else
          cVar1S24S74P064P011N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='1' AND A( 1)='1' AND E( 4)='1' )then
          cVar1S25S74P064P011P017P054nsss(0) <='1';
          else
          cVar1S25S74P064P011P017P054nsss(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='1' AND A( 1)='1' AND E( 4)='0' )then
          cVar1S26S74P064P011P017N054(0) <='1';
          else
          cVar1S26S74P064P011P017N054(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='1' AND A( 1)='1' AND E( 4)='0' )then
          cVar1S27S74P064P011P017N054(0) <='1';
          else
          cVar1S27S74P064P011P017N054(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='1' AND A( 1)='0' AND A( 5)='1' )then
          cVar1S28S74P064P011N017P009(0) <='1';
          else
          cVar1S28S74P064P011N017P009(0) <='0';
          end if;
        if(D( 1)='1' AND A( 4)='1' AND A( 1)='0' AND A( 5)='0' )then
          cVar1S29S74P064P011N017N009(0) <='1';
          else
          cVar1S29S74P064P011N017N009(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='1' AND E(13)='1' )then
          cVar1S0S75P029P011P051nsss(0) <='1';
          else
          cVar1S0S75P029P011P051nsss(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='1' AND E(13)='0' AND E( 4)='1' )then
          cVar1S1S75P029P011N051P054(0) <='1';
          else
          cVar1S1S75P029P011N051P054(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='1' AND E(13)='0' AND E( 4)='1' )then
          cVar1S2S75P029P011N051P054(0) <='1';
          else
          cVar1S2S75P029P011N051P054(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='1' AND E(13)='0' AND E( 4)='0' )then
          cVar1S3S75P029P011N051N054(0) <='1';
          else
          cVar1S3S75P029P011N051N054(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='1' AND D( 4)='1' )then
          cVar1S4S75P029N011P010P052nsss(0) <='1';
          else
          cVar1S4S75P029N011P010P052nsss(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='1' AND D( 4)='0' )then
          cVar1S5S75P029N011P010N052(0) <='1';
          else
          cVar1S5S75P029N011P010N052(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='0' AND A( 5)='1' )then
          cVar1S6S75P029N011N010P009(0) <='1';
          else
          cVar1S6S75P029N011N010P009(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='0' AND A( 5)='1' )then
          cVar1S7S75P029N011N010P009(0) <='1';
          else
          cVar1S7S75P029N011N010P009(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='0' AND A( 5)='1' )then
          cVar1S8S75P029N011N010P009(0) <='1';
          else
          cVar1S8S75P029N011N010P009(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='0' AND A( 5)='0' )then
          cVar1S9S75P029N011N010N009(0) <='1';
          else
          cVar1S9S75P029N011N010N009(0) <='0';
          end if;
        if(B( 5)='1' AND A( 4)='0' AND A(14)='0' AND A( 5)='0' )then
          cVar1S10S75P029N011N010N009(0) <='1';
          else
          cVar1S10S75P029N011N010N009(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S11S75N029P041P020P003nsss(0) <='1';
          else
          cVar1S11S75N029P041P020P003nsss(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S12S75N029P041P020N003(0) <='1';
          else
          cVar1S12S75N029P041P020N003(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S13S75N029P041P020N003(0) <='1';
          else
          cVar1S13S75N029P041P020N003(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S14S75N029P041P020N003(0) <='1';
          else
          cVar1S14S75N029P041P020N003(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S15S75N029P041N020P005(0) <='1';
          else
          cVar1S15S75N029P041N020P005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S16S75N029P041N020P005(0) <='1';
          else
          cVar1S16S75N029P041N020P005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='1' )then
          cVar1S17S75N029P041N020P005(0) <='1';
          else
          cVar1S17S75N029P041N020P005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S18S75N029P041N020N005(0) <='1';
          else
          cVar1S18S75N029P041N020N005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='1' AND B(19)='0' AND A( 7)='0' )then
          cVar1S19S75N029P041N020N005(0) <='1';
          else
          cVar1S19S75N029P041N020N005(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='1' AND B( 8)='1' )then
          cVar1S20S75N029N041P045P023nsss(0) <='1';
          else
          cVar1S20S75N029N041P045P023nsss(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='1' AND B( 8)='0' )then
          cVar1S21S75N029N041P045N023(0) <='1';
          else
          cVar1S21S75N029N041P045N023(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='1' AND B( 8)='0' )then
          cVar1S22S75N029N041P045N023(0) <='1';
          else
          cVar1S22S75N029N041P045N023(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='1' AND B( 8)='0' )then
          cVar1S23S75N029N041P045N023(0) <='1';
          else
          cVar1S23S75N029N041P045N023(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='0' AND B( 6)='1' )then
          cVar1S24S75N029N041N045P027(0) <='1';
          else
          cVar1S24S75N029N041N045P027(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='0' AND B( 6)='1' )then
          cVar1S25S75N029N041N045P027(0) <='1';
          else
          cVar1S25S75N029N041N045P027(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='0' AND B( 6)='0' )then
          cVar1S26S75N029N041N045N027(0) <='1';
          else
          cVar1S26S75N029N041N045N027(0) <='0';
          end if;
        if(B( 5)='0' AND D(15)='0' AND D(14)='0' AND B( 6)='0' )then
          cVar1S27S75N029N041N045N027(0) <='1';
          else
          cVar1S27S75N029N041N045N027(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='0' AND A( 5)='1' )then
          cVar1S0S76P064P027P066P009(0) <='1';
          else
          cVar1S0S76P064P027P066P009(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='0' AND A( 5)='1' )then
          cVar1S1S76P064P027P066P009(0) <='1';
          else
          cVar1S1S76P064P027P066P009(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='0' AND A( 5)='0' )then
          cVar1S2S76P064P027P066N009(0) <='1';
          else
          cVar1S2S76P064P027P066N009(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='1' AND D( 0)='0' )then
          cVar1S3S76P064P027P066P068nsss(0) <='1';
          else
          cVar1S3S76P064P027P066P068nsss(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='1' AND D( 0)='1' )then
          cVar1S4S76P064P027P066P068(0) <='1';
          else
          cVar1S4S76P064P027P066P068(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='1' AND E( 1)='1' AND D( 0)='1' )then
          cVar1S5S76P064P027P066P068(0) <='1';
          else
          cVar1S5S76P064P027P066P068(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='1' )then
          cVar1S6S76P064N027P041P020(0) <='1';
          else
          cVar1S6S76P064N027P041P020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='1' )then
          cVar1S7S76P064N027P041P020(0) <='1';
          else
          cVar1S7S76P064N027P041P020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='1' )then
          cVar1S8S76P064N027P041P020(0) <='1';
          else
          cVar1S8S76P064N027P041P020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='0' )then
          cVar1S9S76P064N027P041N020(0) <='1';
          else
          cVar1S9S76P064N027P041N020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='0' )then
          cVar1S10S76P064N027P041N020(0) <='1';
          else
          cVar1S10S76P064N027P041N020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='1' AND B(19)='0' )then
          cVar1S11S76P064N027P041N020(0) <='1';
          else
          cVar1S11S76P064N027P041N020(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='0' )then
          cVar1S12S76P064N027N041P039(0) <='1';
          else
          cVar1S12S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='0' )then
          cVar1S13S76P064N027N041P039(0) <='1';
          else
          cVar1S13S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='0' )then
          cVar1S14S76P064N027N041P039(0) <='1';
          else
          cVar1S14S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='0' )then
          cVar1S15S76P064N027N041P039(0) <='1';
          else
          cVar1S15S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='1' )then
          cVar1S16S76P064N027N041P039(0) <='1';
          else
          cVar1S16S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='0' AND B( 6)='0' AND D(15)='0' AND B( 0)='1' )then
          cVar1S17S76P064N027N041P039(0) <='1';
          else
          cVar1S17S76P064N027N041P039(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='1' )then
          cVar1S18S76P064P042nsss(0) <='1';
          else
          cVar1S18S76P064P042nsss(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='0' AND B( 6)='0' )then
          cVar1S19S76P064N042P008P027(0) <='1';
          else
          cVar1S19S76P064N042P008P027(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='0' AND B( 6)='0' )then
          cVar1S20S76P064N042P008P027(0) <='1';
          else
          cVar1S20S76P064N042P008P027(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='0' AND B( 6)='0' )then
          cVar1S21S76P064N042P008P027(0) <='1';
          else
          cVar1S21S76P064N042P008P027(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='0' AND B( 6)='1' )then
          cVar1S22S76P064N042P008P027(0) <='1';
          else
          cVar1S22S76P064N042P008P027(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='1' AND A(14)='0' )then
          cVar1S23S76P064N042P008P010(0) <='1';
          else
          cVar1S23S76P064N042P008P010(0) <='0';
          end if;
        if(D( 1)='1' AND E( 7)='0' AND A(15)='1' AND A(14)='0' )then
          cVar1S24S76P064N042P008P010(0) <='1';
          else
          cVar1S24S76P064N042P008P010(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='1' AND B( 2)='0' )then
          cVar1S0S77P017P064P034P035(0) <='1';
          else
          cVar1S0S77P017P064P034P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='1' AND B( 2)='0' )then
          cVar1S1S77P017P064P034P035(0) <='1';
          else
          cVar1S1S77P017P064P034P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='1' AND B( 2)='1' )then
          cVar1S2S77P017P064P034P035(0) <='1';
          else
          cVar1S2S77P017P064P034P035(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='1' )then
          cVar1S3S77P017P064N034P020(0) <='1';
          else
          cVar1S3S77P017P064N034P020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='1' )then
          cVar1S4S77P017P064N034P020(0) <='1';
          else
          cVar1S4S77P017P064N034P020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='1' )then
          cVar1S5S77P017P064N034P020(0) <='1';
          else
          cVar1S5S77P017P064N034P020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='0' )then
          cVar1S6S77P017P064N034N020(0) <='1';
          else
          cVar1S6S77P017P064N034N020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='0' )then
          cVar1S7S77P017P064N034N020(0) <='1';
          else
          cVar1S7S77P017P064N034N020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='0' AND B(12)='0' AND B(19)='0' )then
          cVar1S8S77P017P064N034N020(0) <='1';
          else
          cVar1S8S77P017P064N034N020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND E( 5)='1' AND A(11)='0' )then
          cVar1S9S77P017P064P050P016nsss(0) <='1';
          else
          cVar1S9S77P017P064P050P016nsss(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND E( 5)='0' AND B(19)='0' )then
          cVar1S10S77P017P064N050P020(0) <='1';
          else
          cVar1S10S77P017P064N050P020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND E( 5)='0' AND B(19)='0' )then
          cVar1S11S77P017P064N050P020(0) <='1';
          else
          cVar1S11S77P017P064N050P020(0) <='0';
          end if;
        if(A( 1)='1' AND D( 1)='1' AND E( 5)='0' AND B(19)='0' )then
          cVar1S12S77P017P064N050P020(0) <='1';
          else
          cVar1S12S77P017P064N050P020(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S13S77N017P041P020P003nsss(0) <='1';
          else
          cVar1S13S77N017P041P020P003nsss(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S14S77N017P041P020N003(0) <='1';
          else
          cVar1S14S77N017P041P020N003(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S15S77N017P041P020N003(0) <='1';
          else
          cVar1S15S77N017P041P020N003(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='0' AND A( 2)='0' )then
          cVar1S16S77N017P041N020P015(0) <='1';
          else
          cVar1S16S77N017P041N020P015(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='0' AND A( 2)='0' )then
          cVar1S17S77N017P041N020P015(0) <='1';
          else
          cVar1S17S77N017P041N020P015(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='0' AND A( 2)='0' )then
          cVar1S18S77N017P041N020P015(0) <='1';
          else
          cVar1S18S77N017P041N020P015(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='1' AND B(19)='0' AND A( 2)='1' )then
          cVar1S19S77N017P041N020P015(0) <='1';
          else
          cVar1S19S77N017P041N020P015(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S20S77N017N041P062P027(0) <='1';
          else
          cVar1S20S77N017N041P062P027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S21S77N017N041P062P027(0) <='1';
          else
          cVar1S21S77N017N041P062P027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='1' )then
          cVar1S22S77N017N041P062P027(0) <='1';
          else
          cVar1S22S77N017N041P062P027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S23S77N017N041P062N027(0) <='1';
          else
          cVar1S23S77N017N041P062N027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S24S77N017N041P062N027(0) <='1';
          else
          cVar1S24S77N017N041P062N027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S25S77N017N041P062N027(0) <='1';
          else
          cVar1S25S77N017N041P062N027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='0' AND B( 6)='0' )then
          cVar1S26S77N017N041P062N027(0) <='1';
          else
          cVar1S26S77N017N041P062N027(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='1' AND A(14)='0' )then
          cVar1S27S77N017N041P062P010(0) <='1';
          else
          cVar1S27S77N017N041P062P010(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='1' AND A(14)='0' )then
          cVar1S28S77N017N041P062P010(0) <='1';
          else
          cVar1S28S77N017N041P062P010(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='1' AND A(14)='0' )then
          cVar1S29S77N017N041P062P010(0) <='1';
          else
          cVar1S29S77N017N041P062P010(0) <='0';
          end if;
        if(A( 1)='0' AND D(15)='0' AND E( 2)='1' AND A(14)='1' )then
          cVar1S30S77N017N041P062P010(0) <='1';
          else
          cVar1S30S77N017N041P062P010(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S0S78P062P063P007P025(0) <='1';
          else
          cVar1S0S78P062P063P007P025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S1S78P062P063P007P025(0) <='1';
          else
          cVar1S1S78P062P063P007P025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S2S78P062P063P007N025(0) <='1';
          else
          cVar1S2S78P062P063P007N025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S3S78P062P063P007N025(0) <='1';
          else
          cVar1S3S78P062P063P007N025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S4S78P062P063P007N025(0) <='1';
          else
          cVar1S4S78P062P063P007N025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S5S78P062P063P007N025(0) <='1';
          else
          cVar1S5S78P062P063P007N025(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='1' )then
          cVar1S6S78P062P063N007P029(0) <='1';
          else
          cVar1S6S78P062P063N007P029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='1' )then
          cVar1S7S78P062P063N007P029(0) <='1';
          else
          cVar1S7S78P062P063N007P029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='1' )then
          cVar1S8S78P062P063N007P029(0) <='1';
          else
          cVar1S8S78P062P063N007P029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='0' )then
          cVar1S9S78P062P063N007N029(0) <='1';
          else
          cVar1S9S78P062P063N007N029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='0' )then
          cVar1S10S78P062P063N007N029(0) <='1';
          else
          cVar1S10S78P062P063N007N029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='0' )then
          cVar1S11S78P062P063N007N029(0) <='1';
          else
          cVar1S11S78P062P063N007N029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='0' AND A( 6)='0' AND B( 5)='0' )then
          cVar1S12S78P062P063N007N029(0) <='1';
          else
          cVar1S12S78P062P063N007N029(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='1' AND E( 3)='0' )then
          cVar1S13S78P062P063P035P058(0) <='1';
          else
          cVar1S13S78P062P063P035P058(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='1' AND E( 3)='0' )then
          cVar1S14S78P062P063P035P058(0) <='1';
          else
          cVar1S14S78P062P063P035P058(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='1' AND E( 3)='0' )then
          cVar1S15S78P062P063P035P058(0) <='1';
          else
          cVar1S15S78P062P063P035P058(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='0' AND B(12)='1' )then
          cVar1S16S78P062P063N035P034(0) <='1';
          else
          cVar1S16S78P062P063N035P034(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='0' AND B(12)='1' )then
          cVar1S17S78P062P063N035P034(0) <='1';
          else
          cVar1S17S78P062P063N035P034(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='0' AND B(12)='0' )then
          cVar1S18S78P062P063N035N034(0) <='1';
          else
          cVar1S18S78P062P063N035N034(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='0' AND B(12)='0' )then
          cVar1S19S78P062P063N035N034(0) <='1';
          else
          cVar1S19S78P062P063N035N034(0) <='0';
          end if;
        if(E( 2)='0' AND E(10)='1' AND B( 2)='0' AND B(12)='0' )then
          cVar1S20S78P062P063N035N034(0) <='1';
          else
          cVar1S20S78P062P063N035N034(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='1' )then
          cVar1S21S78P062P026P027P060(0) <='1';
          else
          cVar1S21S78P062P026P027P060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='1' )then
          cVar1S22S78P062P026P027P060(0) <='1';
          else
          cVar1S22S78P062P026P027P060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='1' )then
          cVar1S23S78P062P026P027P060(0) <='1';
          else
          cVar1S23S78P062P026P027P060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='0' )then
          cVar1S24S78P062P026P027N060(0) <='1';
          else
          cVar1S24S78P062P026P027N060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='0' )then
          cVar1S25S78P062P026P027N060(0) <='1';
          else
          cVar1S25S78P062P026P027N060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='0' )then
          cVar1S26S78P062P026P027N060(0) <='1';
          else
          cVar1S26S78P062P026P027N060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 6)='0' AND D( 2)='0' )then
          cVar1S27S78P062P026P027N060(0) <='1';
          else
          cVar1S27S78P062P026P027N060(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='1' AND D( 0)='1' )then
          cVar1S28S78P062P026P068nsss(0) <='1';
          else
          cVar1S28S78P062P026P068nsss(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='1' AND D( 9)='0' AND B(15)='1' )then
          cVar1S0S79P051P008P065P028nsss(0) <='1';
          else
          cVar1S0S79P051P008P065P028nsss(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='1' AND D( 9)='0' AND B(15)='0' )then
          cVar1S1S79P051P008P065N028(0) <='1';
          else
          cVar1S1S79P051P008P065N028(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='1' AND D( 9)='0' AND B(15)='0' )then
          cVar1S2S79P051P008P065N028(0) <='1';
          else
          cVar1S2S79P051P008P065N028(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='1' )then
          cVar1S3S79P051N008P042nsss(0) <='1';
          else
          cVar1S3S79P051N008P042nsss(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='1' )then
          cVar1S4S79P051N008N042P009(0) <='1';
          else
          cVar1S4S79P051N008N042P009(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='1' )then
          cVar1S5S79P051N008N042P009(0) <='1';
          else
          cVar1S5S79P051N008N042P009(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='1' )then
          cVar1S6S79P051N008N042P009(0) <='1';
          else
          cVar1S6S79P051N008N042P009(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='0' )then
          cVar1S7S79P051N008N042N009(0) <='1';
          else
          cVar1S7S79P051N008N042N009(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='0' )then
          cVar1S8S79P051N008N042N009(0) <='1';
          else
          cVar1S8S79P051N008N042N009(0) <='0';
          end if;
        if(E(13)='1' AND A(15)='0' AND E( 7)='0' AND A( 5)='0' )then
          cVar1S9S79P051N008N042N009(0) <='1';
          else
          cVar1S9S79P051N008N042N009(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S10S79N051P041P020P003nsss(0) <='1';
          else
          cVar1S10S79N051P041P020P003nsss(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S11S79N051P041P020N003(0) <='1';
          else
          cVar1S11S79N051P041P020N003(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S12S79N051P041P020N003(0) <='1';
          else
          cVar1S12S79N051P041P020N003(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S13S79N051P041P020N003(0) <='1';
          else
          cVar1S13S79N051P041P020N003(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='1' )then
          cVar1S14S79N051P041N020P001nsss(0) <='1';
          else
          cVar1S14S79N051P041N020P001nsss(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S15S79N051P041N020N001(0) <='1';
          else
          cVar1S15S79N051P041N020N001(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S16S79N051P041N020N001(0) <='1';
          else
          cVar1S16S79N051P041N020N001(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='1' AND B(19)='0' AND A( 9)='0' )then
          cVar1S17S79N051P041N020N001(0) <='1';
          else
          cVar1S17S79N051P041N020N001(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='1' )then
          cVar1S18S79N051N041P047P026(0) <='1';
          else
          cVar1S18S79N051N041P047P026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='1' )then
          cVar1S19S79N051N041P047P026(0) <='1';
          else
          cVar1S19S79N051N041P047P026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='0' )then
          cVar1S20S79N051N041P047N026(0) <='1';
          else
          cVar1S20S79N051N041P047N026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='0' )then
          cVar1S21S79N051N041P047N026(0) <='1';
          else
          cVar1S21S79N051N041P047N026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='0' )then
          cVar1S22S79N051N041P047N026(0) <='1';
          else
          cVar1S22S79N051N041P047N026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='1' AND B(16)='0' )then
          cVar1S23S79N051N041P047N026(0) <='1';
          else
          cVar1S23S79N051N041P047N026(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='0' )then
          cVar1S24S79N051N041N047P049(0) <='1';
          else
          cVar1S24S79N051N041N047P049(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='0' )then
          cVar1S25S79N051N041N047P049(0) <='1';
          else
          cVar1S25S79N051N041N047P049(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='0' )then
          cVar1S26S79N051N041N047P049(0) <='1';
          else
          cVar1S26S79N051N041N047P049(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='1' )then
          cVar1S27S79N051N041N047P049(0) <='1';
          else
          cVar1S27S79N051N041N047P049(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='1' )then
          cVar1S28S79N051N041N047P049(0) <='1';
          else
          cVar1S28S79N051N041N047P049(0) <='0';
          end if;
        if(E(13)='0' AND D(15)='0' AND E(14)='0' AND D(13)='1' )then
          cVar1S29S79N051N041N047P049(0) <='1';
          else
          cVar1S29S79N051N041N047P049(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='1' )then
          cVar1S0S80P040P002P021nsss(0) <='1';
          else
          cVar1S0S80P040P002P021nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='1' )then
          cVar1S1S80P040P002N021P041nsss(0) <='1';
          else
          cVar1S1S80P040P002N021P041nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='0' )then
          cVar1S2S80P040P002N021N041(0) <='1';
          else
          cVar1S2S80P040P002N021N041(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='1' )then
          cVar1S3S80P040N002P057nsss(0) <='1';
          else
          cVar1S3S80P040N002P057nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S4S80P040N002N057P004(0) <='1';
          else
          cVar1S4S80P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S5S80P040N002N057P004(0) <='1';
          else
          cVar1S5S80P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S6S80P040N002N057P004(0) <='1';
          else
          cVar1S6S80P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='0' )then
          cVar1S7S80P040N002N057N004(0) <='1';
          else
          cVar1S7S80P040N002N057N004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='0' )then
          cVar1S8S80P040N002N057N004(0) <='1';
          else
          cVar1S8S80P040N002N057N004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='0' )then
          cVar1S9S80P040N002N057N004(0) <='1';
          else
          cVar1S9S80P040N002N057N004(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S10S80N040P021P007P025(0) <='1';
          else
          cVar1S10S80N040P021P007P025(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S11S80N040P021P007P025(0) <='1';
          else
          cVar1S11S80N040P021P007P025(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S12S80N040P021P007N025(0) <='1';
          else
          cVar1S12S80N040P021P007N025(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S13S80N040P021P007N025(0) <='1';
          else
          cVar1S13S80N040P021P007N025(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='1' )then
          cVar1S14S80N040P021N007P028(0) <='1';
          else
          cVar1S14S80N040P021N007P028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='1' )then
          cVar1S15S80N040P021N007P028(0) <='1';
          else
          cVar1S15S80N040P021N007P028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='0' )then
          cVar1S16S80N040P021N007N028(0) <='1';
          else
          cVar1S16S80N040P021N007N028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='0' )then
          cVar1S17S80N040P021N007N028(0) <='1';
          else
          cVar1S17S80N040P021N007N028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='0' )then
          cVar1S18S80N040P021N007N028(0) <='1';
          else
          cVar1S18S80N040P021N007N028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='0' AND A( 6)='0' AND B(15)='0' )then
          cVar1S19S80N040P021N007N028(0) <='1';
          else
          cVar1S19S80N040P021N007N028(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='1' AND E( 7)='1' )then
          cVar1S20S80N040P021P042nsss(0) <='1';
          else
          cVar1S20S80N040P021P042nsss(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='1' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S21S80N040P021N042P003(0) <='1';
          else
          cVar1S21S80N040P021N042P003(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='1' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S22S80N040P021N042P003(0) <='1';
          else
          cVar1S22S80N040P021N042P003(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='1' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S23S80N040P021N042N003(0) <='1';
          else
          cVar1S23S80N040P021N042N003(0) <='0';
          end if;
        if(D( 7)='0' AND B( 9)='1' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S24S80N040P021N042N003(0) <='1';
          else
          cVar1S24S80N040P021N042N003(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' )then
          cVar1S0S81P040P002nsss(0) <='1';
          else
          cVar1S0S81P040P002nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='1' )then
          cVar1S1S81P040N002P057nsss(0) <='1';
          else
          cVar1S1S81P040N002P057nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S2S81P040N002N057P004(0) <='1';
          else
          cVar1S2S81P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S3S81P040N002N057P004(0) <='1';
          else
          cVar1S3S81P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='1' )then
          cVar1S4S81P040N002N057P004(0) <='1';
          else
          cVar1S4S81P040N002N057P004(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND D(11)='0' AND A(17)='0' )then
          cVar1S5S81P040N002N057N004(0) <='1';
          else
          cVar1S5S81P040N002N057N004(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='1' AND B( 5)='0' AND D(12)='1' )then
          cVar1S6S81N040P028P029P053(0) <='1';
          else
          cVar1S6S81N040P028P029P053(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='1' AND B( 5)='0' AND D(12)='1' )then
          cVar1S7S81N040P028P029P053(0) <='1';
          else
          cVar1S7S81N040P028P029P053(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='1' AND B( 5)='0' AND D(12)='0' )then
          cVar1S8S81N040P028P029N053(0) <='1';
          else
          cVar1S8S81N040P028P029N053(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='1' AND B( 5)='0' AND D(12)='0' )then
          cVar1S9S81N040P028P029N053(0) <='1';
          else
          cVar1S9S81N040P028P029N053(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='1' )then
          cVar1S10S81N040N028P029P011(0) <='1';
          else
          cVar1S10S81N040N028P029P011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='1' )then
          cVar1S11S81N040N028P029P011(0) <='1';
          else
          cVar1S11S81N040N028P029P011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='1' )then
          cVar1S12S81N040N028P029P011(0) <='1';
          else
          cVar1S12S81N040N028P029P011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar1S13S81N040N028P029N011(0) <='1';
          else
          cVar1S13S81N040N028P029N011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar1S14S81N040N028P029N011(0) <='1';
          else
          cVar1S14S81N040N028P029N011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar1S15S81N040N028P029N011(0) <='1';
          else
          cVar1S15S81N040N028P029N011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar1S16S81N040N028P029N011(0) <='1';
          else
          cVar1S16S81N040N028P029N011(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='1' )then
          cVar1S17S81N040N028N029P007(0) <='1';
          else
          cVar1S17S81N040N028N029P007(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='1' )then
          cVar1S18S81N040N028N029P007(0) <='1';
          else
          cVar1S18S81N040N028N029P007(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='1' )then
          cVar1S19S81N040N028N029P007(0) <='1';
          else
          cVar1S19S81N040N028N029P007(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='0' )then
          cVar1S20S81N040N028N029N007(0) <='1';
          else
          cVar1S20S81N040N028N029N007(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='0' )then
          cVar1S21S81N040N028N029N007(0) <='1';
          else
          cVar1S21S81N040N028N029N007(0) <='0';
          end if;
        if(D( 7)='0' AND B(15)='0' AND B( 5)='0' AND A( 6)='0' )then
          cVar1S22S81N040N028N029N007(0) <='1';
          else
          cVar1S22S81N040N028N029N007(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='1' AND A( 5)='0' )then
          cVar1S0S82P062P007P025P009(0) <='1';
          else
          cVar1S0S82P062P007P025P009(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='1' AND A( 5)='1' )then
          cVar1S1S82P062P007P025P009(0) <='1';
          else
          cVar1S1S82P062P007P025P009(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='1' )then
          cVar1S2S82P062P007N025P003(0) <='1';
          else
          cVar1S2S82P062P007N025P003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='1' )then
          cVar1S3S82P062P007N025P003(0) <='1';
          else
          cVar1S3S82P062P007N025P003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='0' )then
          cVar1S4S82P062P007N025N003(0) <='1';
          else
          cVar1S4S82P062P007N025N003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='0' )then
          cVar1S5S82P062P007N025N003(0) <='1';
          else
          cVar1S5S82P062P007N025N003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='0' )then
          cVar1S6S82P062P007N025N003(0) <='1';
          else
          cVar1S6S82P062P007N025N003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='1' AND B( 7)='0' AND A( 8)='0' )then
          cVar1S7S82P062P007N025N003(0) <='1';
          else
          cVar1S7S82P062P007N025N003(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='0' )then
          cVar1S8S82P062N007P015P032(0) <='1';
          else
          cVar1S8S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='0' )then
          cVar1S9S82P062N007P015P032(0) <='1';
          else
          cVar1S9S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='0' )then
          cVar1S10S82P062N007P015P032(0) <='1';
          else
          cVar1S10S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='1' )then
          cVar1S11S82P062N007P015P032(0) <='1';
          else
          cVar1S11S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='1' )then
          cVar1S12S82P062N007P015P032(0) <='1';
          else
          cVar1S12S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='1' )then
          cVar1S13S82P062N007P015P032(0) <='1';
          else
          cVar1S13S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='0' AND B(13)='1' )then
          cVar1S14S82P062N007P015P032(0) <='1';
          else
          cVar1S14S82P062N007P015P032(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='1' AND B( 5)='1' )then
          cVar1S15S82P062N007P015P029(0) <='1';
          else
          cVar1S15S82P062N007P015P029(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='1' AND B( 5)='0' )then
          cVar1S16S82P062N007P015N029(0) <='1';
          else
          cVar1S16S82P062N007P015N029(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='1' AND B( 5)='0' )then
          cVar1S17S82P062N007P015N029(0) <='1';
          else
          cVar1S17S82P062N007P015N029(0) <='0';
          end if;
        if(E( 2)='0' AND A( 6)='0' AND A( 2)='1' AND B( 5)='0' )then
          cVar1S18S82P062N007P015N029(0) <='1';
          else
          cVar1S18S82P062N007P015N029(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 5)='0' AND E( 5)='1' )then
          cVar1S19S82P062P026P029P050(0) <='1';
          else
          cVar1S19S82P062P026P029P050(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 5)='0' AND E( 5)='1' )then
          cVar1S20S82P062P026P029P050(0) <='1';
          else
          cVar1S20S82P062P026P029P050(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S21S82P062P026P029N050(0) <='1';
          else
          cVar1S21S82P062P026P029N050(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 5)='0' AND E( 5)='0' )then
          cVar1S22S82P062P026P029N050(0) <='1';
          else
          cVar1S22S82P062P026P029N050(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='0' AND B( 5)='1' AND B(11)='0' )then
          cVar1S23S82P062P026P029P036(0) <='1';
          else
          cVar1S23S82P062P026P029P036(0) <='0';
          end if;
        if(E( 2)='1' AND B(16)='1' AND B( 1)='1' AND A( 0)='1' )then
          cVar1S24S82P062P026P037P019nsss(0) <='1';
          else
          cVar1S24S82P062P026P037P019nsss(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='1' AND E( 6)='1' AND A( 4)='0' )then
          cVar1S0S83P007P025P046P011nsss(0) <='1';
          else
          cVar1S0S83P007P025P046P011nsss(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='1' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S1S83P007P025N046P009(0) <='1';
          else
          cVar1S1S83P007P025N046P009(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='1' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S2S83P007P025N046P009(0) <='1';
          else
          cVar1S2S83P007P025N046P009(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='1' AND E( 6)='0' AND A( 5)='0' )then
          cVar1S3S83P007P025N046P009(0) <='1';
          else
          cVar1S3S83P007P025N046P009(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='0' AND E(10)='0' )then
          cVar1S4S83P007N025P034P063(0) <='1';
          else
          cVar1S4S83P007N025P034P063(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='0' AND E(10)='0' )then
          cVar1S5S83P007N025P034P063(0) <='1';
          else
          cVar1S5S83P007N025P034P063(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='0' AND E(10)='0' )then
          cVar1S6S83P007N025P034P063(0) <='1';
          else
          cVar1S6S83P007N025P034P063(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='0' AND E(10)='1' )then
          cVar1S7S83P007N025P034P063(0) <='1';
          else
          cVar1S7S83P007N025P034P063(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='0' AND E(10)='1' )then
          cVar1S8S83P007N025P034P063(0) <='1';
          else
          cVar1S8S83P007N025P034P063(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='1' AND A( 0)='1' )then
          cVar1S9S83P007N025P034P019(0) <='1';
          else
          cVar1S9S83P007N025P034P019(0) <='0';
          end if;
        if(A( 6)='1' AND B( 7)='0' AND B(12)='1' AND A( 0)='0' )then
          cVar1S10S83P007N025P034N019(0) <='1';
          else
          cVar1S10S83P007N025P034N019(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S11S83N007P040P002nsss(0) <='1';
          else
          cVar1S11S83N007P040P002nsss(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='1' AND A(18)='0' AND E(14)='1' )then
          cVar1S12S83N007P040N002P047nsss(0) <='1';
          else
          cVar1S12S83N007P040N002P047nsss(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='1' AND A(18)='0' AND E(14)='0' )then
          cVar1S13S83N007P040N002N047(0) <='1';
          else
          cVar1S13S83N007P040N002N047(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='1' AND A(18)='0' AND E(14)='0' )then
          cVar1S14S83N007P040N002N047(0) <='1';
          else
          cVar1S14S83N007P040N002N047(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='1' AND A(18)='0' AND E(14)='0' )then
          cVar1S15S83N007P040N002N047(0) <='1';
          else
          cVar1S15S83N007P040N002N047(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='1' AND B(10)='0' )then
          cVar1S16S83N007N040P015P038(0) <='1';
          else
          cVar1S16S83N007N040P015P038(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='1' AND B(10)='0' )then
          cVar1S17S83N007N040P015P038(0) <='1';
          else
          cVar1S17S83N007N040P015P038(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='1' )then
          cVar1S18S83N007N040N015P034(0) <='1';
          else
          cVar1S18S83N007N040N015P034(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='1' )then
          cVar1S19S83N007N040N015P034(0) <='1';
          else
          cVar1S19S83N007N040N015P034(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='0' )then
          cVar1S20S83N007N040N015N034(0) <='1';
          else
          cVar1S20S83N007N040N015N034(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='0' )then
          cVar1S21S83N007N040N015N034(0) <='1';
          else
          cVar1S21S83N007N040N015N034(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='0' )then
          cVar1S22S83N007N040N015N034(0) <='1';
          else
          cVar1S22S83N007N040N015N034(0) <='0';
          end if;
        if(A( 6)='0' AND D( 7)='0' AND A( 2)='0' AND B(12)='0' )then
          cVar1S23S83N007N040N015N034(0) <='1';
          else
          cVar1S23S83N007N040N015N034(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='1' AND A(18)='1' )then
          cVar1S0S84P040P021P002nsss(0) <='1';
          else
          cVar1S0S84P040P021P002nsss(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='1' AND A(18)='0' AND A(13)='0' )then
          cVar1S1S84P040P021N002P012(0) <='1';
          else
          cVar1S1S84P040P021N002P012(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='1' AND A(18)='0' AND A(13)='0' )then
          cVar1S2S84P040P021N002P012(0) <='1';
          else
          cVar1S2S84P040P021N002P012(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='1' AND A(18)='0' AND A(13)='0' )then
          cVar1S3S84P040P021N002P012(0) <='1';
          else
          cVar1S3S84P040P021N002P012(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='0' AND D(11)='1' )then
          cVar1S4S84P040N021P057nsss(0) <='1';
          else
          cVar1S4S84P040N021P057nsss(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='0' AND D(11)='0' AND A(15)='0' )then
          cVar1S5S84P040N021N057P008(0) <='1';
          else
          cVar1S5S84P040N021N057P008(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='0' AND D(11)='0' AND A(15)='0' )then
          cVar1S6S84P040N021N057P008(0) <='1';
          else
          cVar1S6S84P040N021N057P008(0) <='0';
          end if;
        if(D( 7)='1' AND B( 9)='0' AND D(11)='0' AND A(15)='0' )then
          cVar1S7S84P040N021N057P008(0) <='1';
          else
          cVar1S7S84P040N021N057P008(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='1' AND E( 6)='1' )then
          cVar1S8S84N040P007P025P046(0) <='1';
          else
          cVar1S8S84N040P007P025P046(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='1' AND E( 6)='0' )then
          cVar1S9S84N040P007P025N046(0) <='1';
          else
          cVar1S9S84N040P007P025N046(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='1' AND E( 6)='0' )then
          cVar1S10S84N040P007P025N046(0) <='1';
          else
          cVar1S10S84N040P007P025N046(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='1' AND E( 6)='0' )then
          cVar1S11S84N040P007P025N046(0) <='1';
          else
          cVar1S11S84N040P007P025N046(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='0' AND E(12)='0' )then
          cVar1S12S84N040P007N025P055(0) <='1';
          else
          cVar1S12S84N040P007N025P055(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='0' AND E(12)='0' )then
          cVar1S13S84N040P007N025P055(0) <='1';
          else
          cVar1S13S84N040P007N025P055(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='0' AND E(12)='0' )then
          cVar1S14S84N040P007N025P055(0) <='1';
          else
          cVar1S14S84N040P007N025P055(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='1' AND B( 7)='0' AND E(12)='1' )then
          cVar1S15S84N040P007N025P055(0) <='1';
          else
          cVar1S15S84N040P007N025P055(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='0' )then
          cVar1S16S84N040N007P015P001(0) <='1';
          else
          cVar1S16S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='0' )then
          cVar1S17S84N040N007P015P001(0) <='1';
          else
          cVar1S17S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='0' )then
          cVar1S18S84N040N007P015P001(0) <='1';
          else
          cVar1S18S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='1' )then
          cVar1S19S84N040N007P015P001(0) <='1';
          else
          cVar1S19S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='1' )then
          cVar1S20S84N040N007P015P001(0) <='1';
          else
          cVar1S20S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='0' AND A( 9)='1' )then
          cVar1S21S84N040N007P015P001(0) <='1';
          else
          cVar1S21S84N040N007P015P001(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='1' )then
          cVar1S22S84N040N007P015P035(0) <='1';
          else
          cVar1S22S84N040N007P015P035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='1' )then
          cVar1S23S84N040N007P015P035(0) <='1';
          else
          cVar1S23S84N040N007P015P035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='1' )then
          cVar1S24S84N040N007P015P035(0) <='1';
          else
          cVar1S24S84N040N007P015P035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='0' )then
          cVar1S25S84N040N007P015N035(0) <='1';
          else
          cVar1S25S84N040N007P015N035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='0' )then
          cVar1S26S84N040N007P015N035(0) <='1';
          else
          cVar1S26S84N040N007P015N035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='0' )then
          cVar1S27S84N040N007P015N035(0) <='1';
          else
          cVar1S27S84N040N007P015N035(0) <='0';
          end if;
        if(D( 7)='0' AND A( 6)='0' AND A( 2)='1' AND B( 2)='0' )then
          cVar1S28S84N040N007P015N035(0) <='1';
          else
          cVar1S28S84N040N007P015N035(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='1' AND A( 7)='1' )then
          cVar1S0S85P015P032P005nsss(0) <='1';
          else
          cVar1S0S85P015P032P005nsss(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='1' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S1S85P015P032N005P003(0) <='1';
          else
          cVar1S1S85P015P032N005P003(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='1' AND A( 7)='0' AND A( 8)='0' )then
          cVar1S2S85P015P032N005P003(0) <='1';
          else
          cVar1S2S85P015P032N005P003(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='1' AND A(15)='0' )then
          cVar1S3S85P015N032P011P008(0) <='1';
          else
          cVar1S3S85P015N032P011P008(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='1' AND A(15)='1' )then
          cVar1S4S85P015N032P011P008(0) <='1';
          else
          cVar1S4S85P015N032P011P008(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='0' AND A(19)='1' )then
          cVar1S5S85P015N032N011P000(0) <='1';
          else
          cVar1S5S85P015N032N011P000(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='0' AND A(19)='1' )then
          cVar1S6S85P015N032N011P000(0) <='1';
          else
          cVar1S6S85P015N032N011P000(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='0' AND A(19)='1' )then
          cVar1S7S85P015N032N011P000(0) <='1';
          else
          cVar1S7S85P015N032N011P000(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='0' AND A(19)='0' )then
          cVar1S8S85P015N032N011N000(0) <='1';
          else
          cVar1S8S85P015N032N011N000(0) <='0';
          end if;
        if(A( 2)='1' AND B(13)='0' AND A( 4)='0' AND A(19)='0' )then
          cVar1S9S85P015N032N011N000(0) <='1';
          else
          cVar1S9S85P015N032N011N000(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='1' )then
          cVar1S10S85N015P021P038nsss(0) <='1';
          else
          cVar1S10S85N015P021P038nsss(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S11S85N015P021N038P014(0) <='1';
          else
          cVar1S11S85N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S12S85N015P021N038P014(0) <='1';
          else
          cVar1S12S85N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S13S85N015P021N038P014(0) <='1';
          else
          cVar1S13S85N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='1' )then
          cVar1S14S85N015P021N038P014(0) <='1';
          else
          cVar1S14S85N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='1' AND A(17)='1' )then
          cVar1S15S85N015N021P044P004nsss(0) <='1';
          else
          cVar1S15S85N015N021P044P004nsss(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='1' AND A(17)='0' )then
          cVar1S16S85N015N021P044N004(0) <='1';
          else
          cVar1S16S85N015N021P044N004(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='1' AND A(17)='0' )then
          cVar1S17S85N015N021P044N004(0) <='1';
          else
          cVar1S17S85N015N021P044N004(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='1' AND A(17)='0' )then
          cVar1S18S85N015N021P044N004(0) <='1';
          else
          cVar1S18S85N015N021P044N004(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='0' AND A( 7)='0' )then
          cVar1S19S85N015N021N044P005(0) <='1';
          else
          cVar1S19S85N015N021N044P005(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='0' AND A( 7)='0' )then
          cVar1S20S85N015N021N044P005(0) <='1';
          else
          cVar1S20S85N015N021N044P005(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='0' AND A( 7)='0' )then
          cVar1S21S85N015N021N044P005(0) <='1';
          else
          cVar1S21S85N015N021N044P005(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='0' AND A( 7)='1' )then
          cVar1S22S85N015N021N044P005(0) <='1';
          else
          cVar1S22S85N015N021N044P005(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND D( 6)='0' AND A( 7)='1' )then
          cVar1S23S85N015N021N044P005(0) <='1';
          else
          cVar1S23S85N015N021N044P005(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='1' AND A(18)='1' )then
          cVar1S0S86P021P038P002nsss(0) <='1';
          else
          cVar1S0S86P021P038P002nsss(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S1S86P021P038N002P004nsss(0) <='1';
          else
          cVar1S1S86P021P038N002P004nsss(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S2S86P021P038N002N004(0) <='1';
          else
          cVar1S2S86P021P038N002N004(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S3S86P021P038N002N004(0) <='1';
          else
          cVar1S3S86P021P038N002N004(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='0' AND A(14)='0' AND E( 7)='1' )then
          cVar1S4S86P021N038P010P042nsss(0) <='1';
          else
          cVar1S4S86P021N038P010P042nsss(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='0' AND A(14)='0' AND E( 7)='0' )then
          cVar1S5S86P021N038P010N042(0) <='1';
          else
          cVar1S5S86P021N038P010N042(0) <='0';
          end if;
        if(B( 9)='1' AND B(10)='0' AND A(14)='1' AND A( 0)='1' )then
          cVar1S6S86P021N038P010P019nsss(0) <='1';
          else
          cVar1S6S86P021N038P010P019nsss(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='1' AND A( 8)='1' )then
          cVar1S7S86N021P020P039P003nsss(0) <='1';
          else
          cVar1S7S86N021P020P039P003nsss(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='1' AND A( 8)='0' )then
          cVar1S8S86N021P020P039N003(0) <='1';
          else
          cVar1S8S86N021P020P039N003(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='1' AND A( 8)='0' )then
          cVar1S9S86N021P020P039N003(0) <='1';
          else
          cVar1S9S86N021P020P039N003(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='1' AND A( 8)='0' )then
          cVar1S10S86N021P020P039N003(0) <='1';
          else
          cVar1S10S86N021P020P039N003(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='0' AND B( 4)='0' )then
          cVar1S11S86N021P020N039P031(0) <='1';
          else
          cVar1S11S86N021P020N039P031(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='0' AND B( 4)='0' )then
          cVar1S12S86N021P020N039P031(0) <='1';
          else
          cVar1S12S86N021P020N039P031(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='0' AND B( 4)='0' )then
          cVar1S13S86N021P020N039P031(0) <='1';
          else
          cVar1S13S86N021P020N039P031(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='1' AND B( 0)='0' AND B( 4)='0' )then
          cVar1S14S86N021P020N039P031(0) <='1';
          else
          cVar1S14S86N021P020N039P031(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='1' )then
          cVar1S15S86N021N020P002P015(0) <='1';
          else
          cVar1S15S86N021N020P002P015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='1' )then
          cVar1S16S86N021N020P002P015(0) <='1';
          else
          cVar1S16S86N021N020P002P015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='1' )then
          cVar1S17S86N021N020P002P015(0) <='1';
          else
          cVar1S17S86N021N020P002P015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='0' )then
          cVar1S18S86N021N020P002N015(0) <='1';
          else
          cVar1S18S86N021N020P002N015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='0' )then
          cVar1S19S86N021N020P002N015(0) <='1';
          else
          cVar1S19S86N021N020P002N015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='0' AND A( 2)='0' )then
          cVar1S20S86N021N020P002N015(0) <='1';
          else
          cVar1S20S86N021N020P002N015(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='1' AND A(17)='1' )then
          cVar1S21S86N021N020P002P004(0) <='1';
          else
          cVar1S21S86N021N020P002P004(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='1' AND A(17)='1' )then
          cVar1S22S86N021N020P002P004(0) <='1';
          else
          cVar1S22S86N021N020P002P004(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='1' AND A(17)='0' )then
          cVar1S23S86N021N020P002N004(0) <='1';
          else
          cVar1S23S86N021N020P002N004(0) <='0';
          end if;
        if(B( 9)='0' AND B(19)='0' AND A(18)='1' AND A(17)='0' )then
          cVar1S24S86N021N020P002N004(0) <='1';
          else
          cVar1S24S86N021N020P002N004(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='1' )then
          cVar1S0S87P015P055P061P032nsss(0) <='1';
          else
          cVar1S0S87P015P055P061P032nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='0' )then
          cVar1S1S87P015P055P061N032(0) <='1';
          else
          cVar1S1S87P015P055P061N032(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='0' )then
          cVar1S2S87P015P055P061N032(0) <='1';
          else
          cVar1S2S87P015P055P061N032(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='0' )then
          cVar1S3S87P015P055P061N032(0) <='1';
          else
          cVar1S3S87P015P055P061N032(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='0' AND B(19)='1' )then
          cVar1S4S87P015N055P021P020(0) <='1';
          else
          cVar1S4S87P015N055P021P020(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='0' AND B(19)='1' )then
          cVar1S5S87P015N055P021P020(0) <='1';
          else
          cVar1S5S87P015N055P021P020(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='0' AND B(19)='0' )then
          cVar1S6S87P015N055P021N020(0) <='1';
          else
          cVar1S6S87P015N055P021N020(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='0' AND B(19)='0' )then
          cVar1S7S87P015N055P021N020(0) <='1';
          else
          cVar1S7S87P015N055P021N020(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='0' AND B(19)='0' )then
          cVar1S8S87P015N055P021N020(0) <='1';
          else
          cVar1S8S87P015N055P021N020(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='1' AND E( 1)='1' )then
          cVar1S9S87P015N055P021P066nsss(0) <='1';
          else
          cVar1S9S87P015N055P021P066nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='1' AND E( 1)='0' )then
          cVar1S10S87P015N055P021N066(0) <='1';
          else
          cVar1S10S87P015N055P021N066(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B( 9)='1' AND E( 1)='0' )then
          cVar1S11S87P015N055P021N066(0) <='1';
          else
          cVar1S11S87P015N055P021N066(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='1' )then
          cVar1S12S87N015P021P038nsss(0) <='1';
          else
          cVar1S12S87N015P021P038nsss(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S13S87N015P021N038P014(0) <='1';
          else
          cVar1S13S87N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S14S87N015P021N038P014(0) <='1';
          else
          cVar1S14S87N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S15S87N015P021N038P014(0) <='1';
          else
          cVar1S15S87N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='0' )then
          cVar1S16S87N015P021N038P014(0) <='1';
          else
          cVar1S16S87N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='1' AND B(10)='0' AND A(12)='1' )then
          cVar1S17S87N015P021N038P014(0) <='1';
          else
          cVar1S17S87N015P021N038P014(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='1' AND B( 0)='1' )then
          cVar1S18S87N015N021P020P039nsss(0) <='1';
          else
          cVar1S18S87N015N021P020P039nsss(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='1' AND B( 0)='0' )then
          cVar1S19S87N015N021P020N039(0) <='1';
          else
          cVar1S19S87N015N021P020N039(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='1' AND B( 0)='0' )then
          cVar1S20S87N015N021P020N039(0) <='1';
          else
          cVar1S20S87N015N021P020N039(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='0' )then
          cVar1S21S87N015N021N020P057(0) <='1';
          else
          cVar1S21S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='0' )then
          cVar1S22S87N015N021N020P057(0) <='1';
          else
          cVar1S22S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='0' )then
          cVar1S23S87N015N021N020P057(0) <='1';
          else
          cVar1S23S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='1' )then
          cVar1S24S87N015N021N020P057(0) <='1';
          else
          cVar1S24S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='1' )then
          cVar1S25S87N015N021N020P057(0) <='1';
          else
          cVar1S25S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='1' )then
          cVar1S26S87N015N021N020P057(0) <='1';
          else
          cVar1S26S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND B( 9)='0' AND B(19)='0' AND D(11)='1' )then
          cVar1S27S87N015N021N020P057(0) <='1';
          else
          cVar1S27S87N015N021N020P057(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='1' )then
          cVar1S0S88P015P057P055P039(0) <='1';
          else
          cVar1S0S88P015P057P055P039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='1' )then
          cVar1S1S88P015P057P055P039(0) <='1';
          else
          cVar1S1S88P015P057P055P039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='0' )then
          cVar1S2S88P015P057P055N039(0) <='1';
          else
          cVar1S2S88P015P057P055N039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='0' )then
          cVar1S3S88P015P057P055N039(0) <='1';
          else
          cVar1S3S88P015P057P055N039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='0' )then
          cVar1S4S88P015P057P055N039(0) <='1';
          else
          cVar1S4S88P015P057P055N039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='0' AND B( 0)='0' )then
          cVar1S5S88P015P057P055N039(0) <='1';
          else
          cVar1S5S88P015P057P055N039(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='1' AND D( 8)='1' )then
          cVar1S6S88P015P057P055P069nsss(0) <='1';
          else
          cVar1S6S88P015P057P055P069nsss(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='1' AND D( 8)='0' )then
          cVar1S7S88P015P057P055N069(0) <='1';
          else
          cVar1S7S88P015P057P055N069(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='1' AND D( 8)='0' )then
          cVar1S8S88P015P057P055N069(0) <='1';
          else
          cVar1S8S88P015P057P055N069(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='0' AND E(12)='1' AND D( 8)='0' )then
          cVar1S9S88P015P057P055N069(0) <='1';
          else
          cVar1S9S88P015P057P055N069(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='1' AND E(12)='1' )then
          cVar1S10S88P015P057P010P055(0) <='1';
          else
          cVar1S10S88P015P057P010P055(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='1' AND E(12)='1' )then
          cVar1S11S88P015P057P010P055(0) <='1';
          else
          cVar1S11S88P015P057P010P055(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar1S12S88P015P057N010P013(0) <='1';
          else
          cVar1S12S88P015P057N010P013(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar1S13S88P015P057N010P013(0) <='1';
          else
          cVar1S13S88P015P057N010P013(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S14S88P015P057N010N013(0) <='1';
          else
          cVar1S14S88P015P057N010N013(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S15S88P015P057N010N013(0) <='1';
          else
          cVar1S15S88P015P057N010N013(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S16S88P015P057N010N013(0) <='1';
          else
          cVar1S16S88P015P057N010N013(0) <='0';
          end if;
        if(A( 2)='0' AND D(11)='1' AND A(14)='0' AND A( 3)='0' )then
          cVar1S17S88P015P057N010N013(0) <='1';
          else
          cVar1S17S88P015P057N010N013(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='1' )then
          cVar1S18S88P015P055P061P032nsss(0) <='1';
          else
          cVar1S18S88P015P055P061P032nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='0' )then
          cVar1S19S88P015P055P061N032(0) <='1';
          else
          cVar1S19S88P015P055P061N032(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='1' AND D(10)='0' AND B(13)='0' )then
          cVar1S20S88P015P055P061N032(0) <='1';
          else
          cVar1S20S88P015P055P061N032(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='1' AND A(18)='1' )then
          cVar1S21S88P015N055P020P002nsss(0) <='1';
          else
          cVar1S21S88P015N055P020P002nsss(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='1' AND A(18)='0' )then
          cVar1S22S88P015N055P020N002(0) <='1';
          else
          cVar1S22S88P015N055P020N002(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='0' AND A( 5)='1' )then
          cVar1S23S88P015N055N020P009(0) <='1';
          else
          cVar1S23S88P015N055N020P009(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='0' AND A( 5)='1' )then
          cVar1S24S88P015N055N020P009(0) <='1';
          else
          cVar1S24S88P015N055N020P009(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='0' AND A( 5)='0' )then
          cVar1S25S88P015N055N020N009(0) <='1';
          else
          cVar1S25S88P015N055N020N009(0) <='0';
          end if;
        if(A( 2)='1' AND E(12)='0' AND B(19)='0' AND A( 5)='0' )then
          cVar1S26S88P015N055N020N009(0) <='1';
          else
          cVar1S26S88P015N055N020N009(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='1' )then
          cVar1S0S89P015P013P008P059(0) <='1';
          else
          cVar1S0S89P015P013P008P059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='1' )then
          cVar1S1S89P015P013P008P059(0) <='1';
          else
          cVar1S1S89P015P013P008P059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='1' )then
          cVar1S2S89P015P013P008P059(0) <='1';
          else
          cVar1S2S89P015P013P008P059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='0' )then
          cVar1S3S89P015P013P008N059(0) <='1';
          else
          cVar1S3S89P015P013P008N059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='0' )then
          cVar1S4S89P015P013P008N059(0) <='1';
          else
          cVar1S4S89P015P013P008N059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='0' AND E(11)='0' )then
          cVar1S5S89P015P013P008N059(0) <='1';
          else
          cVar1S5S89P015P013P008N059(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='1' AND A( 0)='1' )then
          cVar1S6S89P015P013P008P019(0) <='1';
          else
          cVar1S6S89P015P013P008P019(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='1' AND A( 0)='1' )then
          cVar1S7S89P015P013P008P019(0) <='1';
          else
          cVar1S7S89P015P013P008P019(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND A(15)='1' AND A( 0)='0' )then
          cVar1S8S89P015P013P008N019(0) <='1';
          else
          cVar1S8S89P015P013P008N019(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='0' AND E(12)='1' )then
          cVar1S9S89P015P013P059P055(0) <='1';
          else
          cVar1S9S89P015P013P059P055(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='0' AND E(12)='0' )then
          cVar1S10S89P015P013P059N055(0) <='1';
          else
          cVar1S10S89P015P013P059N055(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='0' AND E(12)='0' )then
          cVar1S11S89P015P013P059N055(0) <='1';
          else
          cVar1S11S89P015P013P059N055(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='0' AND E(12)='0' )then
          cVar1S12S89P015P013P059N055(0) <='1';
          else
          cVar1S12S89P015P013P059N055(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='0' AND E(12)='0' )then
          cVar1S13S89P015P013P059N055(0) <='1';
          else
          cVar1S13S89P015P013P059N055(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='1' AND D(10)='1' )then
          cVar1S14S89P015P013P059P061(0) <='1';
          else
          cVar1S14S89P015P013P059P061(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND E(11)='1' AND D(10)='1' )then
          cVar1S15S89P015P013P059P061(0) <='1';
          else
          cVar1S15S89P015P013P059P061(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='1' AND B(19)='1' AND A( 8)='1' )then
          cVar1S16S89N015P039P020P003nsss(0) <='1';
          else
          cVar1S16S89N015P039P020P003nsss(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S17S89N015P039P020N003(0) <='1';
          else
          cVar1S17S89N015P039P020N003(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='1' AND B(19)='1' AND A( 8)='0' )then
          cVar1S18S89N015P039P020N003(0) <='1';
          else
          cVar1S18S89N015P039P020N003(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='1' AND B(19)='0' AND A( 1)='0' )then
          cVar1S19S89N015P039N020P017(0) <='1';
          else
          cVar1S19S89N015P039N020P017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='1' AND B(19)='0' AND A( 1)='0' )then
          cVar1S20S89N015P039N020P017(0) <='1';
          else
          cVar1S20S89N015P039N020P017(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='1' AND B( 7)='1' )then
          cVar1S21S89N015N039P044P025(0) <='1';
          else
          cVar1S21S89N015N039P044P025(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='1' AND B( 7)='0' )then
          cVar1S22S89N015N039P044N025(0) <='1';
          else
          cVar1S22S89N015N039P044N025(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='1' AND B( 7)='0' )then
          cVar1S23S89N015N039P044N025(0) <='1';
          else
          cVar1S23S89N015N039P044N025(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='1' AND B( 7)='0' )then
          cVar1S24S89N015N039P044N025(0) <='1';
          else
          cVar1S24S89N015N039P044N025(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='0' AND B(10)='1' )then
          cVar1S25S89N015N039N044P038(0) <='1';
          else
          cVar1S25S89N015N039N044P038(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='0' AND B(10)='1' )then
          cVar1S26S89N015N039N044P038(0) <='1';
          else
          cVar1S26S89N015N039N044P038(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='0' AND B(10)='0' )then
          cVar1S27S89N015N039N044N038(0) <='1';
          else
          cVar1S27S89N015N039N044N038(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='0' AND B(10)='0' )then
          cVar1S28S89N015N039N044N038(0) <='1';
          else
          cVar1S28S89N015N039N044N038(0) <='0';
          end if;
        if(A( 2)='0' AND B( 0)='0' AND D( 6)='0' AND B(10)='0' )then
          cVar1S29S89N015N039N044N038(0) <='1';
          else
          cVar1S29S89N015N039N044N038(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='1' )then
          cVar1S0S90P020P039P010P003nsss(0) <='1';
          else
          cVar1S0S90P020P039P010P003nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='0' )then
          cVar1S1S90P020P039P010N003(0) <='1';
          else
          cVar1S1S90P020P039P010N003(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='1' )then
          cVar1S2S90P020N039P025nsss(0) <='1';
          else
          cVar1S2S90P020N039P025nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S3S90P020N039N025P031(0) <='1';
          else
          cVar1S3S90P020N039N025P031(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S4S90P020N039N025P031(0) <='1';
          else
          cVar1S4S90P020N039N025P031(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='1' )then
          cVar1S5S90N020P040P021P002nsss(0) <='1';
          else
          cVar1S5S90N020P040P021P002nsss(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S6S90N020P040P021N002(0) <='1';
          else
          cVar1S6S90N020P040P021N002(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S7S90N020P040P021N002(0) <='1';
          else
          cVar1S7S90N020P040P021N002(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='1' AND A(18)='0' )then
          cVar1S8S90N020P040P021N002(0) <='1';
          else
          cVar1S8S90N020P040P021N002(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='0' AND D(11)='1' )then
          cVar1S9S90N020P040N021P057nsss(0) <='1';
          else
          cVar1S9S90N020P040N021P057nsss(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='1' AND B( 9)='0' AND D(11)='0' )then
          cVar1S10S90N020P040N021N057(0) <='1';
          else
          cVar1S10S90N020P040N021N057(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S11S90N020N040P039P045(0) <='1';
          else
          cVar1S11S90N020N040P039P045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S12S90N020N040P039P045(0) <='1';
          else
          cVar1S12S90N020N040P039P045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='1' )then
          cVar1S13S90N020N040P039P045(0) <='1';
          else
          cVar1S13S90N020N040P039P045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S14S90N020N040P039N045(0) <='1';
          else
          cVar1S14S90N020N040P039N045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S15S90N020N040P039N045(0) <='1';
          else
          cVar1S15S90N020N040P039N045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S16S90N020N040P039N045(0) <='1';
          else
          cVar1S16S90N020N040P039N045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='0' AND D(14)='0' )then
          cVar1S17S90N020N040P039N045(0) <='1';
          else
          cVar1S17S90N020N040P039N045(0) <='0';
          end if;
        if(B(19)='0' AND D( 7)='0' AND B( 0)='1' AND A( 7)='1' )then
          cVar1S18S90N020N040P039P005nsss(0) <='1';
          else
          cVar1S18S90N020N040P039P005nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='1' )then
          cVar1S0S91P020P039P010P003nsss(0) <='1';
          else
          cVar1S0S91P020P039P010P003nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='0' )then
          cVar1S1S91P020P039P010N003(0) <='1';
          else
          cVar1S1S91P020P039P010N003(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='1' )then
          cVar1S2S91P020N039P025nsss(0) <='1';
          else
          cVar1S2S91P020N039P025nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B(17)='1' )then
          cVar1S3S91P020N039N025P024nsss(0) <='1';
          else
          cVar1S3S91P020N039N025P024nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S4S91P020N039N025N024(0) <='1';
          else
          cVar1S4S91P020N039N025N024(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B(17)='0' )then
          cVar1S5S91P020N039N025N024(0) <='1';
          else
          cVar1S5S91P020N039N025N024(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='1' AND A(10)='0' )then
          cVar1S6S91N020P045P004P018nsss(0) <='1';
          else
          cVar1S6S91N020P045P004P018nsss(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='1' AND A(10)='1' )then
          cVar1S7S91N020P045P004P018(0) <='1';
          else
          cVar1S7S91N020P045P004P018(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='1' )then
          cVar1S8S91N020P045N004P006(0) <='1';
          else
          cVar1S8S91N020P045N004P006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='1' )then
          cVar1S9S91N020P045N004P006(0) <='1';
          else
          cVar1S9S91N020P045N004P006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S10S91N020P045N004N006(0) <='1';
          else
          cVar1S10S91N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S11S91N020P045N004N006(0) <='1';
          else
          cVar1S11S91N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S12S91N020P045N004N006(0) <='1';
          else
          cVar1S12S91N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S13S91N020N045P040P021nsss(0) <='1';
          else
          cVar1S13S91N020N045P040P021nsss(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S14S91N020N045P040N021(0) <='1';
          else
          cVar1S14S91N020N045P040N021(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S15S91N020N045P040N021(0) <='1';
          else
          cVar1S15S91N020N045P040N021(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='1' )then
          cVar1S16S91N020N045N040P055(0) <='1';
          else
          cVar1S16S91N020N045N040P055(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='1' )then
          cVar1S17S91N020N045N040P055(0) <='1';
          else
          cVar1S17S91N020N045N040P055(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='1' )then
          cVar1S18S91N020N045N040P055(0) <='1';
          else
          cVar1S18S91N020N045N040P055(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='0' )then
          cVar1S19S91N020N045N040N055(0) <='1';
          else
          cVar1S19S91N020N045N040N055(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='0' )then
          cVar1S20S91N020N045N040N055(0) <='1';
          else
          cVar1S20S91N020N045N040N055(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND E(12)='0' )then
          cVar1S21S91N020N045N040N055(0) <='1';
          else
          cVar1S21S91N020N045N040N055(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='1' )then
          cVar1S0S92P020P039P010P003nsss(0) <='1';
          else
          cVar1S0S92P020P039P010P003nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='0' )then
          cVar1S1S92P020P039P010N003(0) <='1';
          else
          cVar1S1S92P020P039P010N003(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='1' AND A(14)='0' AND A( 8)='0' )then
          cVar1S2S92P020P039P010N003(0) <='1';
          else
          cVar1S2S92P020P039P010N003(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='1' )then
          cVar1S3S92P020N039P025nsss(0) <='1';
          else
          cVar1S3S92P020N039P025nsss(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S4S92P020N039N025P031(0) <='1';
          else
          cVar1S4S92P020N039N025P031(0) <='0';
          end if;
        if(B(19)='1' AND B( 0)='0' AND B( 7)='0' AND B( 4)='0' )then
          cVar1S5S92P020N039N025P031(0) <='1';
          else
          cVar1S5S92P020N039N025P031(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='1' AND A(10)='0' )then
          cVar1S6S92N020P045P004P018nsss(0) <='1';
          else
          cVar1S6S92N020P045P004P018nsss(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='1' AND A(10)='1' )then
          cVar1S7S92N020P045P004P018(0) <='1';
          else
          cVar1S7S92N020P045P004P018(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='1' )then
          cVar1S8S92N020P045N004P006(0) <='1';
          else
          cVar1S8S92N020P045N004P006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='1' )then
          cVar1S9S92N020P045N004P006(0) <='1';
          else
          cVar1S9S92N020P045N004P006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S10S92N020P045N004N006(0) <='1';
          else
          cVar1S10S92N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S11S92N020P045N004N006(0) <='1';
          else
          cVar1S11S92N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='1' AND A(17)='0' AND A(16)='0' )then
          cVar1S12S92N020P045N004N006(0) <='1';
          else
          cVar1S12S92N020P045N004N006(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar1S13S92N020N045P040P021nsss(0) <='1';
          else
          cVar1S13S92N020N045P040P021nsss(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S14S92N020N045P040N021(0) <='1';
          else
          cVar1S14S92N020N045P040N021(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='1' AND B( 9)='0' )then
          cVar1S15S92N020N045P040N021(0) <='1';
          else
          cVar1S15S92N020N045P040N021(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S16S92N020N045N040P044(0) <='1';
          else
          cVar1S16S92N020N045N040P044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S17S92N020N045N040P044(0) <='1';
          else
          cVar1S17S92N020N045N040P044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='1' )then
          cVar1S18S92N020N045N040P044(0) <='1';
          else
          cVar1S18S92N020N045N040P044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S19S92N020N045N040N044(0) <='1';
          else
          cVar1S19S92N020N045N040N044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S20S92N020N045N040N044(0) <='1';
          else
          cVar1S20S92N020N045N040N044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S21S92N020N045N040N044(0) <='1';
          else
          cVar1S21S92N020N045N040N044(0) <='0';
          end if;
        if(B(19)='0' AND D(14)='0' AND D( 7)='0' AND D( 6)='0' )then
          cVar1S22S92N020N045N040N044(0) <='1';
          else
          cVar1S22S92N020N045N040N044(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='1' )then
          cVar1S0S93P040P002P021nsss(0) <='1';
          else
          cVar1S0S93P040P002P021nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='1' )then
          cVar1S1S93P040P002N021P041nsss(0) <='1';
          else
          cVar1S1S93P040P002N021P041nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='0' )then
          cVar1S2S93P040P002N021N041(0) <='1';
          else
          cVar1S2S93P040P002N021N041(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='1' )then
          cVar1S3S93P040N002P004P022nsss(0) <='1';
          else
          cVar1S3S93P040N002P004P022nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='0' )then
          cVar1S4S93P040N002P004N022(0) <='1';
          else
          cVar1S4S93P040N002P004N022(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='0' )then
          cVar1S5S93P040N002P004N022(0) <='1';
          else
          cVar1S5S93P040N002P004N022(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='0' AND A(19)='1' )then
          cVar1S6S93P040N002N004P000nsss(0) <='1';
          else
          cVar1S6S93P040N002N004P000nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='0' AND A(19)='0' )then
          cVar1S7S93P040N002N004N000(0) <='1';
          else
          cVar1S7S93P040N002N004N000(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='0' AND A(19)='0' )then
          cVar1S8S93P040N002N004N000(0) <='1';
          else
          cVar1S8S93P040N002N004N000(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='0' AND A(19)='0' )then
          cVar1S9S93P040N002N004N000(0) <='1';
          else
          cVar1S9S93P040N002N004N000(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='1' AND A( 0)='1' )then
          cVar1S10S93N040P045P022P019nsss(0) <='1';
          else
          cVar1S10S93N040P045P022P019nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='1' AND A( 0)='0' )then
          cVar1S11S93N040P045P022N019(0) <='1';
          else
          cVar1S11S93N040P045P022N019(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='1' AND A( 0)='0' )then
          cVar1S12S93N040P045P022N019(0) <='1';
          else
          cVar1S12S93N040P045P022N019(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='1' AND A( 0)='0' )then
          cVar1S13S93N040P045P022N019(0) <='1';
          else
          cVar1S13S93N040P045P022N019(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='0' AND B( 8)='1' )then
          cVar1S14S93N040P045N022P023(0) <='1';
          else
          cVar1S14S93N040P045N022P023(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='0' AND B( 8)='0' )then
          cVar1S15S93N040P045N022N023(0) <='1';
          else
          cVar1S15S93N040P045N022N023(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='1' AND B(18)='0' AND B( 8)='0' )then
          cVar1S16S93N040P045N022N023(0) <='1';
          else
          cVar1S16S93N040P045N022N023(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='1' AND B( 0)='1' )then
          cVar1S17S93N040N045P020P039(0) <='1';
          else
          cVar1S17S93N040N045P020P039(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='1' AND B( 0)='1' )then
          cVar1S18S93N040N045P020P039(0) <='1';
          else
          cVar1S18S93N040N045P020P039(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='1' AND B( 0)='1' )then
          cVar1S19S93N040N045P020P039(0) <='1';
          else
          cVar1S19S93N040N045P020P039(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='1' AND B( 0)='0' )then
          cVar1S20S93N040N045P020N039(0) <='1';
          else
          cVar1S20S93N040N045P020N039(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='1' AND B( 0)='0' )then
          cVar1S21S93N040N045P020N039(0) <='1';
          else
          cVar1S21S93N040N045P020N039(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S22S93N040N045N020P044(0) <='1';
          else
          cVar1S22S93N040N045N020P044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S23S93N040N045N020P044(0) <='1';
          else
          cVar1S23S93N040N045N020P044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='1' )then
          cVar1S24S93N040N045N020P044(0) <='1';
          else
          cVar1S24S93N040N045N020P044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S25S93N040N045N020N044(0) <='1';
          else
          cVar1S25S93N040N045N020N044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S26S93N040N045N020N044(0) <='1';
          else
          cVar1S26S93N040N045N020N044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S27S93N040N045N020N044(0) <='1';
          else
          cVar1S27S93N040N045N020N044(0) <='0';
          end if;
        if(D( 7)='0' AND D(14)='0' AND B(19)='0' AND D( 6)='0' )then
          cVar1S28S93N040N045N020N044(0) <='1';
          else
          cVar1S28S93N040N045N020N044(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='1' )then
          cVar1S0S94P040P002P021nsss(0) <='1';
          else
          cVar1S0S94P040P002P021nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='1' )then
          cVar1S1S94P040P002N021P041nsss(0) <='1';
          else
          cVar1S1S94P040P002N021P041nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='1' AND B( 9)='0' AND D(15)='0' )then
          cVar1S2S94P040P002N021N041(0) <='1';
          else
          cVar1S2S94P040P002N021N041(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='1' )then
          cVar1S3S94P040N002P004P022nsss(0) <='1';
          else
          cVar1S3S94P040N002P004P022nsss(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='0' )then
          cVar1S4S94P040N002P004N022(0) <='1';
          else
          cVar1S4S94P040N002P004N022(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='1' AND B(18)='0' )then
          cVar1S5S94P040N002P004N022(0) <='1';
          else
          cVar1S5S94P040N002P004N022(0) <='0';
          end if;
        if(D( 7)='1' AND A(18)='0' AND A(17)='0' AND B(19)='0' )then
          cVar1S6S94P040N002N004P020nsss(0) <='1';
          else
          cVar1S6S94P040N002N004P020nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='1' AND D( 5)='0' )then
          cVar1S7S94N040P044P006P048(0) <='1';
          else
          cVar1S7S94N040P044P006P048(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='1' AND D( 5)='0' )then
          cVar1S8S94N040P044P006P048(0) <='1';
          else
          cVar1S8S94N040P044P006P048(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='1' )then
          cVar1S9S94N040P044N006P023(0) <='1';
          else
          cVar1S9S94N040P044N006P023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='1' )then
          cVar1S10S94N040P044N006P023(0) <='1';
          else
          cVar1S10S94N040P044N006P023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='1' )then
          cVar1S11S94N040P044N006P023(0) <='1';
          else
          cVar1S11S94N040P044N006P023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='0' )then
          cVar1S12S94N040P044N006N023(0) <='1';
          else
          cVar1S12S94N040P044N006N023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='0' )then
          cVar1S13S94N040P044N006N023(0) <='1';
          else
          cVar1S13S94N040P044N006N023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='1' AND A(16)='0' AND B( 8)='0' )then
          cVar1S14S94N040P044N006N023(0) <='1';
          else
          cVar1S14S94N040P044N006N023(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='1' )then
          cVar1S15S94N040N044P042P020(0) <='1';
          else
          cVar1S15S94N040N044P042P020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='1' )then
          cVar1S16S94N040N044P042P020(0) <='1';
          else
          cVar1S16S94N040N044P042P020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='0' )then
          cVar1S17S94N040N044P042N020(0) <='1';
          else
          cVar1S17S94N040N044P042N020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='0' )then
          cVar1S18S94N040N044P042N020(0) <='1';
          else
          cVar1S18S94N040N044P042N020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='0' )then
          cVar1S19S94N040N044P042N020(0) <='1';
          else
          cVar1S19S94N040N044P042N020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='0' AND B(19)='0' )then
          cVar1S20S94N040N044P042N020(0) <='1';
          else
          cVar1S20S94N040N044P042N020(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='1' )then
          cVar1S21S94N040N044P042P058nsss(0) <='1';
          else
          cVar1S21S94N040N044P042P058nsss(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='0' )then
          cVar1S22S94N040N044P042N058(0) <='1';
          else
          cVar1S22S94N040N044P042N058(0) <='0';
          end if;
        if(D( 7)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='0' )then
          cVar1S23S94N040N044P042N058(0) <='1';
          else
          cVar1S23S94N040N044P042N058(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S0S95P044P023P005nsss(0) <='1';
          else
          cVar1S0S95P044P023P005nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar1S1S95P044P023N005P004nsss(0) <='1';
          else
          cVar1S1S95P044P023N005P004nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S2S95P044P023N005N004(0) <='1';
          else
          cVar1S2S95P044P023N005N004(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='1' AND A( 7)='0' AND A(17)='0' )then
          cVar1S3S95P044P023N005N004(0) <='1';
          else
          cVar1S3S95P044P023N005N004(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='1' )then
          cVar1S4S95P044N023P051nsss(0) <='1';
          else
          cVar1S4S95P044N023P051nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='0' AND D(11)='1' )then
          cVar1S5S95P044N023N051P057nsss(0) <='1';
          else
          cVar1S5S95P044N023N051P057nsss(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='0' AND D(11)='0' )then
          cVar1S6S95P044N023N051N057(0) <='1';
          else
          cVar1S6S95P044N023N051N057(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='0' AND D(11)='0' )then
          cVar1S7S95P044N023N051N057(0) <='1';
          else
          cVar1S7S95P044N023N051N057(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='0' AND D(11)='0' )then
          cVar1S8S95P044N023N051N057(0) <='1';
          else
          cVar1S8S95P044N023N051N057(0) <='0';
          end if;
        if(D( 6)='1' AND B( 8)='0' AND E(13)='0' AND D(11)='0' )then
          cVar1S9S95P044N023N051N057(0) <='1';
          else
          cVar1S9S95P044N023N051N057(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='1' )then
          cVar1S10S95N044P040P002nsss(0) <='1';
          else
          cVar1S10S95N044P040P002nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S11S95N044P040N002P004(0) <='1';
          else
          cVar1S11S95N044P040N002P004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S12S95N044P040N002P004(0) <='1';
          else
          cVar1S12S95N044P040N002P004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='1' )then
          cVar1S13S95N044P040N002P004(0) <='1';
          else
          cVar1S13S95N044P040N002P004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S14S95N044P040N002N004(0) <='1';
          else
          cVar1S14S95N044P040N002N004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S15S95N044P040N002N004(0) <='1';
          else
          cVar1S15S95N044P040N002N004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='1' AND A(18)='0' AND A(17)='0' )then
          cVar1S16S95N044P040N002N004(0) <='1';
          else
          cVar1S16S95N044P040N002N004(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='1' AND B(18)='1' )then
          cVar1S17S95N044N040P045P022nsss(0) <='1';
          else
          cVar1S17S95N044N040P045P022nsss(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S18S95N044N040P045N022(0) <='1';
          else
          cVar1S18S95N044N040P045N022(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S19S95N044N040P045N022(0) <='1';
          else
          cVar1S19S95N044N040P045N022(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S20S95N044N040P045N022(0) <='1';
          else
          cVar1S20S95N044N040P045N022(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S21S95N044N040N045P020(0) <='1';
          else
          cVar1S21S95N044N040N045P020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S22S95N044N040N045P020(0) <='1';
          else
          cVar1S22S95N044N040N045P020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S23S95N044N040N045P020(0) <='1';
          else
          cVar1S23S95N044N040N045P020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S24S95N044N040N045P020(0) <='1';
          else
          cVar1S24S95N044N040N045P020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S25S95N044N040N045N020(0) <='1';
          else
          cVar1S25S95N044N040N045N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S26S95N044N040N045N020(0) <='1';
          else
          cVar1S26S95N044N040N045N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S27S95N044N040N045N020(0) <='1';
          else
          cVar1S27S95N044N040N045N020(0) <='0';
          end if;
        if(D( 6)='0' AND D( 7)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S28S95N044N040N045N020(0) <='1';
          else
          cVar1S28S95N044N040N045N020(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='1' AND B( 8)='1' )then
          cVar1S0S96P044P004P023nsss(0) <='1';
          else
          cVar1S0S96P044P004P023nsss(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='1' AND B( 8)='0' AND B(18)='1' )then
          cVar1S1S96P044P004N023P022(0) <='1';
          else
          cVar1S1S96P044P004N023P022(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='1' )then
          cVar1S2S96P044N004P021nsss(0) <='1';
          else
          cVar1S2S96P044N004P021nsss(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='1' )then
          cVar1S3S96P044N004N021P005(0) <='1';
          else
          cVar1S3S96P044N004N021P005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S4S96P044N004N021N005(0) <='1';
          else
          cVar1S4S96P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S5S96P044N004N021N005(0) <='1';
          else
          cVar1S5S96P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S6S96P044N004N021N005(0) <='1';
          else
          cVar1S6S96P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S7S96P044N004N021N005(0) <='1';
          else
          cVar1S7S96P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S8S96N044P016P012P056(0) <='1';
          else
          cVar1S8S96N044P016P012P056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S9S96N044P016P012P056(0) <='1';
          else
          cVar1S9S96N044P016P012P056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S10S96N044P016P012N056(0) <='1';
          else
          cVar1S10S96N044P016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S11S96N044P016P012N056(0) <='1';
          else
          cVar1S11S96N044P016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S12S96N044P016P012N056(0) <='1';
          else
          cVar1S12S96N044P016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S13S96N044P016P012N056(0) <='1';
          else
          cVar1S13S96N044P016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='1' )then
          cVar1S14S96N044P016N012P053(0) <='1';
          else
          cVar1S14S96N044P016N012P053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='1' )then
          cVar1S15S96N044P016N012P053(0) <='1';
          else
          cVar1S15S96N044P016N012P053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='0' )then
          cVar1S16S96N044P016N012N053(0) <='1';
          else
          cVar1S16S96N044P016N012N053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='0' )then
          cVar1S17S96N044P016N012N053(0) <='1';
          else
          cVar1S17S96N044P016N012N053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S18S96N044P016P052P059(0) <='1';
          else
          cVar1S18S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S19S96N044P016P052P059(0) <='1';
          else
          cVar1S19S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S20S96N044P016P052P059(0) <='1';
          else
          cVar1S20S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S21S96N044P016P052P059(0) <='1';
          else
          cVar1S21S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S22S96N044P016P052P059(0) <='1';
          else
          cVar1S22S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S23S96N044P016P052P059(0) <='1';
          else
          cVar1S23S96N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='1' AND D( 9)='1' )then
          cVar1S24S96N044P016P052P065nsss(0) <='1';
          else
          cVar1S24S96N044P016P052P065nsss(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='1' AND D( 9)='0' )then
          cVar1S25S96N044P016P052N065(0) <='1';
          else
          cVar1S25S96N044P016P052N065(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='1' AND D( 9)='0' )then
          cVar1S26S96N044P016P052N065(0) <='1';
          else
          cVar1S26S96N044P016P052N065(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='1' AND B( 8)='1' )then
          cVar1S0S97P044P004P023nsss(0) <='1';
          else
          cVar1S0S97P044P004P023nsss(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='1' AND B( 8)='0' AND A(11)='0' )then
          cVar1S1S97P044P004N023P016(0) <='1';
          else
          cVar1S1S97P044P004N023P016(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='1' )then
          cVar1S2S97P044N004P021nsss(0) <='1';
          else
          cVar1S2S97P044N004P021nsss(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='1' )then
          cVar1S3S97P044N004N021P005(0) <='1';
          else
          cVar1S3S97P044N004N021P005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='1' )then
          cVar1S4S97P044N004N021P005(0) <='1';
          else
          cVar1S4S97P044N004N021P005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S5S97P044N004N021N005(0) <='1';
          else
          cVar1S5S97P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S6S97P044N004N021N005(0) <='1';
          else
          cVar1S6S97P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='1' AND A(17)='0' AND B( 9)='0' AND A( 7)='0' )then
          cVar1S7S97P044N004N021N005(0) <='1';
          else
          cVar1S7S97P044N004N021N005(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S8S97N044P016P052P059(0) <='1';
          else
          cVar1S8S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S9S97N044P016P052P059(0) <='1';
          else
          cVar1S9S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='0' )then
          cVar1S10S97N044P016P052P059(0) <='1';
          else
          cVar1S10S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S11S97N044P016P052P059(0) <='1';
          else
          cVar1S11S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S12S97N044P016P052P059(0) <='1';
          else
          cVar1S12S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='0' AND E(11)='1' )then
          cVar1S13S97N044P016P052P059(0) <='1';
          else
          cVar1S13S97N044P016P052P059(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='1' AND D( 9)='1' )then
          cVar1S14S97N044P016P052P065nsss(0) <='1';
          else
          cVar1S14S97N044P016P052P065nsss(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='1' AND D( 4)='1' AND D( 9)='0' )then
          cVar1S15S97N044P016P052N065(0) <='1';
          else
          cVar1S15S97N044P016P052N065(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S16S97N044N016P012P056(0) <='1';
          else
          cVar1S16S97N044N016P012P056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S17S97N044N016P012P056(0) <='1';
          else
          cVar1S17S97N044N016P012P056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S18S97N044N016P012N056(0) <='1';
          else
          cVar1S18S97N044N016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S19S97N044N016P012N056(0) <='1';
          else
          cVar1S19S97N044N016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S20S97N044N016P012N056(0) <='1';
          else
          cVar1S20S97N044N016P012N056(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='1' )then
          cVar1S21S97N044N016N012P053(0) <='1';
          else
          cVar1S21S97N044N016N012P053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='1' )then
          cVar1S22S97N044N016N012P053(0) <='1';
          else
          cVar1S22S97N044N016N012P053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='1' )then
          cVar1S23S97N044N016N012P053(0) <='1';
          else
          cVar1S23S97N044N016N012P053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='0' )then
          cVar1S24S97N044N016N012N053(0) <='1';
          else
          cVar1S24S97N044N016N012N053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='0' )then
          cVar1S25S97N044N016N012N053(0) <='1';
          else
          cVar1S25S97N044N016N012N053(0) <='0';
          end if;
        if(D( 6)='0' AND A(11)='0' AND A(13)='0' AND D(12)='0' )then
          cVar1S26S97N044N016N012N053(0) <='1';
          else
          cVar1S26S97N044N016N012N053(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='1' AND B( 8)='1' )then
          cVar1S0S98P016P044P004P023nsss(0) <='1';
          else
          cVar1S0S98P016P044P004P023nsss(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='1' AND B( 8)='0' )then
          cVar1S1S98P016P044P004N023(0) <='1';
          else
          cVar1S1S98P016P044P004N023(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='0' AND E(14)='1' )then
          cVar1S2S98P016P044N004P047nsss(0) <='1';
          else
          cVar1S2S98P016P044N004P047nsss(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='0' AND E(14)='0' )then
          cVar1S3S98P016P044N004N047(0) <='1';
          else
          cVar1S3S98P016P044N004N047(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='0' AND E(14)='0' )then
          cVar1S4S98P016P044N004N047(0) <='1';
          else
          cVar1S4S98P016P044N004N047(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='1' AND A(17)='0' AND E(14)='0' )then
          cVar1S5S98P016P044N004N047(0) <='1';
          else
          cVar1S5S98P016P044N004N047(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S6S98P016N044P012P056(0) <='1';
          else
          cVar1S6S98P016N044P012P056(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='1' AND D( 3)='1' )then
          cVar1S7S98P016N044P012P056(0) <='1';
          else
          cVar1S7S98P016N044P012P056(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S8S98P016N044P012N056(0) <='1';
          else
          cVar1S8S98P016N044P012N056(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S9S98P016N044P012N056(0) <='1';
          else
          cVar1S9S98P016N044P012N056(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='1' AND D( 3)='0' )then
          cVar1S10S98P016N044P012N056(0) <='1';
          else
          cVar1S10S98P016N044P012N056(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='0' )then
          cVar1S11S98P016N044N012P032(0) <='1';
          else
          cVar1S11S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='0' )then
          cVar1S12S98P016N044N012P032(0) <='1';
          else
          cVar1S12S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='0' )then
          cVar1S13S98P016N044N012P032(0) <='1';
          else
          cVar1S13S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='1' )then
          cVar1S14S98P016N044N012P032(0) <='1';
          else
          cVar1S14S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='1' )then
          cVar1S15S98P016N044N012P032(0) <='1';
          else
          cVar1S15S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='0' AND D( 6)='0' AND A(13)='0' AND B(13)='1' )then
          cVar1S16S98P016N044N012P032(0) <='1';
          else
          cVar1S16S98P016N044N012P032(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='1' AND D(12)='1' )then
          cVar1S17S98P016P021P037P053nsss(0) <='1';
          else
          cVar1S17S98P016P021P037P053nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='1' AND D(12)='0' )then
          cVar1S18S98P016P021P037N053(0) <='1';
          else
          cVar1S18S98P016P021P037N053(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='0' )then
          cVar1S19S98P016P021N037P047(0) <='1';
          else
          cVar1S19S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='0' )then
          cVar1S20S98P016P021N037P047(0) <='1';
          else
          cVar1S20S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='0' )then
          cVar1S21S98P016P021N037P047(0) <='1';
          else
          cVar1S21S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='1' )then
          cVar1S22S98P016P021N037P047(0) <='1';
          else
          cVar1S22S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='1' )then
          cVar1S23S98P016P021N037P047(0) <='1';
          else
          cVar1S23S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND B( 1)='0' AND E(14)='1' )then
          cVar1S24S98P016P021N037P047(0) <='1';
          else
          cVar1S24S98P016P021N037P047(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='1' )then
          cVar1S25S98P016P021P069P038nsss(0) <='1';
          else
          cVar1S25S98P016P021P069P038nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='0' )then
          cVar1S26S98P016P021P069N038(0) <='1';
          else
          cVar1S26S98P016P021P069N038(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='0' )then
          cVar1S27S98P016P021P069N038(0) <='1';
          else
          cVar1S27S98P016P021P069N038(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='1' )then
          cVar1S0S99P044P051nsss(0) <='1';
          else
          cVar1S0S99P044P051nsss(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='1' )then
          cVar1S1S99P044N051P057nsss(0) <='1';
          else
          cVar1S1S99P044N051P057nsss(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='0' AND B(13)='1' )then
          cVar1S2S99P044N051N057P032nsss(0) <='1';
          else
          cVar1S2S99P044N051N057P032nsss(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='0' AND B(13)='0' )then
          cVar1S3S99P044N051N057N032(0) <='1';
          else
          cVar1S3S99P044N051N057N032(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='0' AND B(13)='0' )then
          cVar1S4S99P044N051N057N032(0) <='1';
          else
          cVar1S4S99P044N051N057N032(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='0' AND B(13)='0' )then
          cVar1S5S99P044N051N057N032(0) <='1';
          else
          cVar1S5S99P044N051N057N032(0) <='0';
          end if;
        if(D( 6)='1' AND E(13)='0' AND D(11)='0' AND B(13)='0' )then
          cVar1S6S99P044N051N057N032(0) <='1';
          else
          cVar1S6S99P044N051N057N032(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='1' AND B( 0)='1' )then
          cVar1S7S99N044P062P003P039(0) <='1';
          else
          cVar1S7S99N044P062P003P039(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='1' AND B( 0)='1' )then
          cVar1S8S99N044P062P003P039(0) <='1';
          else
          cVar1S8S99N044P062P003P039(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='1' AND B( 0)='0' )then
          cVar1S9S99N044P062P003N039(0) <='1';
          else
          cVar1S9S99N044P062P003N039(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='1' AND B( 0)='0' )then
          cVar1S10S99N044P062P003N039(0) <='1';
          else
          cVar1S10S99N044P062P003N039(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='1' AND B( 0)='0' )then
          cVar1S11S99N044P062P003N039(0) <='1';
          else
          cVar1S11S99N044P062P003N039(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='0' )then
          cVar1S12S99N044P062N003P042(0) <='1';
          else
          cVar1S12S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='0' )then
          cVar1S13S99N044P062N003P042(0) <='1';
          else
          cVar1S13S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='0' )then
          cVar1S14S99N044P062N003P042(0) <='1';
          else
          cVar1S14S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='0' )then
          cVar1S15S99N044P062N003P042(0) <='1';
          else
          cVar1S15S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='1' )then
          cVar1S16S99N044P062N003P042(0) <='1';
          else
          cVar1S16S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='1' )then
          cVar1S17S99N044P062N003P042(0) <='1';
          else
          cVar1S17S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='0' AND A( 8)='0' AND E( 7)='1' )then
          cVar1S18S99N044P062N003P042(0) <='1';
          else
          cVar1S18S99N044P062N003P042(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='1' AND D(12)='1' )then
          cVar1S19S99N044P062P063P053nsss(0) <='1';
          else
          cVar1S19S99N044P062P063P053nsss(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='1' AND D(12)='0' )then
          cVar1S20S99N044P062P063N053(0) <='1';
          else
          cVar1S20S99N044P062P063N053(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='1' AND D(12)='0' )then
          cVar1S21S99N044P062P063N053(0) <='1';
          else
          cVar1S21S99N044P062P063N053(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='0' )then
          cVar1S22S99N044P062N063P009(0) <='1';
          else
          cVar1S22S99N044P062N063P009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='0' )then
          cVar1S23S99N044P062N063P009(0) <='1';
          else
          cVar1S23S99N044P062N063P009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='0' )then
          cVar1S24S99N044P062N063P009(0) <='1';
          else
          cVar1S24S99N044P062N063P009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='0' )then
          cVar1S25S99N044P062N063P009(0) <='1';
          else
          cVar1S25S99N044P062N063P009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='1' )then
          cVar1S26S99N044P062N063P009(0) <='1';
          else
          cVar1S26S99N044P062N063P009(0) <='0';
          end if;
        if(D( 6)='0' AND E( 2)='1' AND E(10)='0' AND A( 5)='1' )then
          cVar1S27S99N044P062N063P009(0) <='1';
          else
          cVar1S27S99N044P062N063P009(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='1' )then
          cVar1S0S100P015P044P004nsss(0) <='1';
          else
          cVar1S0S100P015P044P004nsss(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND B( 9)='1' )then
          cVar1S1S100P015P044N004P021nsss(0) <='1';
          else
          cVar1S1S100P015P044N004P021nsss(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND B( 9)='0' )then
          cVar1S2S100P015P044N004N021(0) <='1';
          else
          cVar1S2S100P015P044N004N021(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND B( 9)='0' )then
          cVar1S3S100P015P044N004N021(0) <='1';
          else
          cVar1S3S100P015P044N004N021(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND B( 9)='0' )then
          cVar1S4S100P015P044N004N021(0) <='1';
          else
          cVar1S4S100P015P044N004N021(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='0' AND D(14)='1' )then
          cVar1S5S100P015N044P062P045nsss(0) <='1';
          else
          cVar1S5S100P015N044P062P045nsss(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='0' AND D(14)='0' )then
          cVar1S6S100P015N044P062N045(0) <='1';
          else
          cVar1S6S100P015N044P062N045(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='0' AND D(14)='0' )then
          cVar1S7S100P015N044P062N045(0) <='1';
          else
          cVar1S7S100P015N044P062N045(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='0' AND D(14)='0' )then
          cVar1S8S100P015N044P062N045(0) <='1';
          else
          cVar1S8S100P015N044P062N045(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='1' )then
          cVar1S9S100P015N044P062P017(0) <='1';
          else
          cVar1S9S100P015N044P062P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='1' )then
          cVar1S10S100P015N044P062P017(0) <='1';
          else
          cVar1S10S100P015N044P062P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='1' )then
          cVar1S11S100P015N044P062P017(0) <='1';
          else
          cVar1S11S100P015N044P062P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='1' )then
          cVar1S12S100P015N044P062P017(0) <='1';
          else
          cVar1S12S100P015N044P062P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar1S13S100P015N044P062N017(0) <='1';
          else
          cVar1S13S100P015N044P062N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar1S14S100P015N044P062N017(0) <='1';
          else
          cVar1S14S100P015N044P062N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar1S15S100P015N044P062N017(0) <='1';
          else
          cVar1S15S100P015N044P062N017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND E( 2)='1' AND A( 1)='0' )then
          cVar1S16S100P015N044P062N017(0) <='1';
          else
          cVar1S16S100P015N044P062N017(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND B(13)='1' )then
          cVar1S17S100P015P013P056P032(0) <='1';
          else
          cVar1S17S100P015P013P056P032(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND B(13)='1' )then
          cVar1S18S100P015P013P056P032(0) <='1';
          else
          cVar1S18S100P015P013P056P032(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND B(13)='0' )then
          cVar1S19S100P015P013P056N032(0) <='1';
          else
          cVar1S19S100P015P013P056N032(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND B(13)='0' )then
          cVar1S20S100P015P013P056N032(0) <='1';
          else
          cVar1S20S100P015P013P056N032(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND B(13)='0' )then
          cVar1S21S100P015P013P056N032(0) <='1';
          else
          cVar1S21S100P015P013P056N032(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='1' AND D( 0)='1' )then
          cVar1S22S100P015P013P056P068(0) <='1';
          else
          cVar1S22S100P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='1' AND D( 0)='0' )then
          cVar1S23S100P015P013P056N068(0) <='1';
          else
          cVar1S23S100P015P013P056N068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='1' )then
          cVar1S24S100P015P013P025nsss(0) <='1';
          else
          cVar1S24S100P015P013P025nsss(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='1' )then
          cVar1S25S100P015P013N025P066(0) <='1';
          else
          cVar1S25S100P015P013N025P066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='1' )then
          cVar1S26S100P015P013N025P066(0) <='1';
          else
          cVar1S26S100P015P013N025P066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='1' )then
          cVar1S27S100P015P013N025P066(0) <='1';
          else
          cVar1S27S100P015P013N025P066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='0' )then
          cVar1S28S100P015P013N025N066(0) <='1';
          else
          cVar1S28S100P015P013N025N066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='0' )then
          cVar1S29S100P015P013N025N066(0) <='1';
          else
          cVar1S29S100P015P013N025N066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 1)='0' )then
          cVar1S30S100P015P013N025N066(0) <='1';
          else
          cVar1S30S100P015P013N025N066(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='0' )then
          cVar1S0S101P015P013P056P068(0) <='1';
          else
          cVar1S0S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='0' )then
          cVar1S1S101P015P013P056P068(0) <='1';
          else
          cVar1S1S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='1' )then
          cVar1S2S101P015P013P056P068(0) <='1';
          else
          cVar1S2S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='1' )then
          cVar1S3S101P015P013P056P068(0) <='1';
          else
          cVar1S3S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='1' )then
          cVar1S4S101P015P013P056P068(0) <='1';
          else
          cVar1S4S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='0' AND D( 0)='1' )then
          cVar1S5S101P015P013P056P068(0) <='1';
          else
          cVar1S5S101P015P013P056P068(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='1' AND E( 5)='1' )then
          cVar1S6S101P015P013P056P050nsss(0) <='1';
          else
          cVar1S6S101P015P013P056P050nsss(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='1' AND E( 5)='0' )then
          cVar1S7S101P015P013P056N050(0) <='1';
          else
          cVar1S7S101P015P013P056N050(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='0' AND D( 3)='1' AND E( 5)='0' )then
          cVar1S8S101P015P013P056N050(0) <='1';
          else
          cVar1S8S101P015P013P056N050(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='1' )then
          cVar1S9S101P015P013P025nsss(0) <='1';
          else
          cVar1S9S101P015P013P025nsss(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 5)='0' )then
          cVar1S10S101P015P013N025P050(0) <='1';
          else
          cVar1S10S101P015P013N025P050(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 5)='0' )then
          cVar1S11S101P015P013N025P050(0) <='1';
          else
          cVar1S11S101P015P013N025P050(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 5)='0' )then
          cVar1S12S101P015P013N025P050(0) <='1';
          else
          cVar1S12S101P015P013N025P050(0) <='0';
          end if;
        if(A( 2)='1' AND A( 3)='1' AND B( 7)='0' AND E( 5)='1' )then
          cVar1S13S101P015P013N025P050(0) <='1';
          else
          cVar1S13S101P015P013N025P050(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='1' AND A( 1)='0' )then
          cVar1S14S101N015P044P025P017(0) <='1';
          else
          cVar1S14S101N015P044P025P017(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='1' AND A( 1)='1' )then
          cVar1S15S101N015P044P025P017psss(0) <='1';
          else
          cVar1S15S101N015P044P025P017psss(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='0' AND A( 7)='1' )then
          cVar1S16S101N015P044N025P005(0) <='1';
          else
          cVar1S16S101N015P044N025P005(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='0' AND A( 7)='0' )then
          cVar1S17S101N015P044N025N005(0) <='1';
          else
          cVar1S17S101N015P044N025N005(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='0' AND A( 7)='0' )then
          cVar1S18S101N015P044N025N005(0) <='1';
          else
          cVar1S18S101N015P044N025N005(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND B( 7)='0' AND A( 7)='0' )then
          cVar1S19S101N015P044N025N005(0) <='1';
          else
          cVar1S19S101N015P044N025N005(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='1' AND D( 4)='0' )then
          cVar1S20S101N015N044P016P052(0) <='1';
          else
          cVar1S20S101N015N044P016P052(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='1' AND D( 4)='0' )then
          cVar1S21S101N015N044P016P052(0) <='1';
          else
          cVar1S21S101N015N044P016P052(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='1' AND D( 4)='0' )then
          cVar1S22S101N015N044P016P052(0) <='1';
          else
          cVar1S22S101N015N044P016P052(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='1' AND D( 4)='0' )then
          cVar1S23S101N015N044P016P052(0) <='1';
          else
          cVar1S23S101N015N044P016P052(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='1' AND D( 4)='1' )then
          cVar1S24S101N015N044P016P052(0) <='1';
          else
          cVar1S24S101N015N044P016P052(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='1' )then
          cVar1S25S101N015N044N016P012(0) <='1';
          else
          cVar1S25S101N015N044N016P012(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='1' )then
          cVar1S26S101N015N044N016P012(0) <='1';
          else
          cVar1S26S101N015N044N016P012(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='1' )then
          cVar1S27S101N015N044N016P012(0) <='1';
          else
          cVar1S27S101N015N044N016P012(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='1' )then
          cVar1S28S101N015N044N016P012(0) <='1';
          else
          cVar1S28S101N015N044N016P012(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='0' )then
          cVar1S29S101N015N044N016N012(0) <='1';
          else
          cVar1S29S101N015N044N016N012(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND A(11)='0' AND A(13)='0' )then
          cVar1S30S101N015N044N016N012(0) <='1';
          else
          cVar1S30S101N015N044N016N012(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='1' )then
          cVar1S0S102P016P015P044nsss(0) <='1';
          else
          cVar1S0S102P016P015P044nsss(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='0' )then
          cVar1S1S102P016P015N044P032(0) <='1';
          else
          cVar1S1S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='0' )then
          cVar1S2S102P016P015N044P032(0) <='1';
          else
          cVar1S2S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='0' )then
          cVar1S3S102P016P015N044P032(0) <='1';
          else
          cVar1S3S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='0' )then
          cVar1S4S102P016P015N044P032(0) <='1';
          else
          cVar1S4S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='1' )then
          cVar1S5S102P016P015N044P032(0) <='1';
          else
          cVar1S5S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='1' )then
          cVar1S6S102P016P015N044P032(0) <='1';
          else
          cVar1S6S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='0' AND D( 6)='0' AND B(13)='1' )then
          cVar1S7S102P016P015N044P032(0) <='1';
          else
          cVar1S7S102P016P015N044P032(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='0' )then
          cVar1S8S102P016P015P043P017(0) <='1';
          else
          cVar1S8S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='0' )then
          cVar1S9S102P016P015P043P017(0) <='1';
          else
          cVar1S9S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='0' )then
          cVar1S10S102P016P015P043P017(0) <='1';
          else
          cVar1S10S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='1' )then
          cVar1S11S102P016P015P043P017(0) <='1';
          else
          cVar1S11S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='1' )then
          cVar1S12S102P016P015P043P017(0) <='1';
          else
          cVar1S12S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='1' )then
          cVar1S13S102P016P015P043P017(0) <='1';
          else
          cVar1S13S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='0' AND A( 1)='1' )then
          cVar1S14S102P016P015P043P017(0) <='1';
          else
          cVar1S14S102P016P015P043P017(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='1' AND A( 7)='1' )then
          cVar1S15S102P016P015P043P005nsss(0) <='1';
          else
          cVar1S15S102P016P015P043P005nsss(0) <='0';
          end if;
        if(A(11)='0' AND A( 2)='1' AND E(15)='1' AND A( 7)='0' )then
          cVar1S16S102P016P015P043N005(0) <='1';
          else
          cVar1S16S102P016P015P043N005(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='0' AND D( 3)='0' )then
          cVar1S17S102P016P021P012P056(0) <='1';
          else
          cVar1S17S102P016P021P012P056(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='0' AND D( 3)='0' )then
          cVar1S18S102P016P021P012P056(0) <='1';
          else
          cVar1S18S102P016P021P012P056(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='0' AND D( 3)='1' )then
          cVar1S19S102P016P021P012P056(0) <='1';
          else
          cVar1S19S102P016P021P012P056(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='0' AND D( 3)='1' )then
          cVar1S20S102P016P021P012P056(0) <='1';
          else
          cVar1S20S102P016P021P012P056(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='1' AND D( 7)='1' )then
          cVar1S21S102P016P021P012P040nsss(0) <='1';
          else
          cVar1S21S102P016P021P012P040nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='1' AND D( 7)='0' )then
          cVar1S22S102P016P021P012N040(0) <='1';
          else
          cVar1S22S102P016P021P012N040(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='1' AND D( 7)='0' )then
          cVar1S23S102P016P021P012N040(0) <='1';
          else
          cVar1S23S102P016P021P012N040(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='0' AND A(13)='1' AND D( 7)='0' )then
          cVar1S24S102P016P021P012N040(0) <='1';
          else
          cVar1S24S102P016P021P012N040(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='1' )then
          cVar1S25S102P016P021P069P038nsss(0) <='1';
          else
          cVar1S25S102P016P021P069P038nsss(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='0' )then
          cVar1S26S102P016P021P069N038(0) <='1';
          else
          cVar1S26S102P016P021P069N038(0) <='0';
          end if;
        if(A(11)='1' AND B( 9)='1' AND D( 8)='0' AND B(10)='0' )then
          cVar1S27S102P016P021P069N038(0) <='1';
          else
          cVar1S27S102P016P021P069N038(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='0' AND B(12)='0' )then
          cVar1S0S103P015P017P063P034(0) <='1';
          else
          cVar1S0S103P015P017P063P034(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='0' AND B(12)='0' )then
          cVar1S1S103P015P017P063P034(0) <='1';
          else
          cVar1S1S103P015P017P063P034(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='0' AND B(12)='0' )then
          cVar1S2S103P015P017P063P034(0) <='1';
          else
          cVar1S2S103P015P017P063P034(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='0' AND B(12)='1' )then
          cVar1S3S103P015P017P063P034(0) <='1';
          else
          cVar1S3S103P015P017P063P034(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='0' AND B(12)='1' )then
          cVar1S4S103P015P017P063P034(0) <='1';
          else
          cVar1S4S103P015P017P063P034(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='1' AND B( 2)='1' )then
          cVar1S5S103P015P017P063P035(0) <='1';
          else
          cVar1S5S103P015P017P063P035(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='1' AND B( 2)='0' )then
          cVar1S6S103P015P017P063N035(0) <='1';
          else
          cVar1S6S103P015P017P063N035(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='1' AND B( 2)='0' )then
          cVar1S7S103P015P017P063N035(0) <='1';
          else
          cVar1S7S103P015P017P063N035(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='0' AND E(10)='1' AND B( 2)='0' )then
          cVar1S8S103P015P017P063N035(0) <='1';
          else
          cVar1S8S103P015P017P063N035(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND B( 2)='0' AND A(12)='1' )then
          cVar1S9S103P015P017P035P014(0) <='1';
          else
          cVar1S9S103P015P017P035P014(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S10S103P015P017P035N014(0) <='1';
          else
          cVar1S10S103P015P017P035N014(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S11S103P015P017P035N014(0) <='1';
          else
          cVar1S11S103P015P017P035N014(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND B( 2)='0' AND A(12)='0' )then
          cVar1S12S103P015P017P035N014(0) <='1';
          else
          cVar1S12S103P015P017P035N014(0) <='0';
          end if;
        if(A( 2)='1' AND A( 1)='1' AND B( 2)='1' AND D( 9)='1' )then
          cVar1S13S103P015P017P035P065(0) <='1';
          else
          cVar1S13S103P015P017P035P065(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='1' AND B( 8)='1' )then
          cVar1S14S103N015P044P004P023nsss(0) <='1';
          else
          cVar1S14S103N015P044P004P023nsss(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='1' AND B( 8)='0' )then
          cVar1S15S103N015P044P004N023(0) <='1';
          else
          cVar1S15S103N015P044P004N023(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND A( 6)='1' )then
          cVar1S16S103N015P044N004P007(0) <='1';
          else
          cVar1S16S103N015P044N004P007(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND A( 6)='1' )then
          cVar1S17S103N015P044N004P007(0) <='1';
          else
          cVar1S17S103N015P044N004P007(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND A( 6)='0' )then
          cVar1S18S103N015P044N004N007(0) <='1';
          else
          cVar1S18S103N015P044N004N007(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND A( 6)='0' )then
          cVar1S19S103N015P044N004N007(0) <='1';
          else
          cVar1S19S103N015P044N004N007(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='1' AND A(17)='0' AND A( 6)='0' )then
          cVar1S20S103N015P044N004N007(0) <='1';
          else
          cVar1S20S103N015P044N004N007(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S21S103N015N044P031P013(0) <='1';
          else
          cVar1S21S103N015N044P031P013(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar1S22S103N015N044P031P013(0) <='1';
          else
          cVar1S22S103N015N044P031P013(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S23S103N015N044P031N013(0) <='1';
          else
          cVar1S23S103N015N044P031N013(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S24S103N015N044P031N013(0) <='1';
          else
          cVar1S24S103N015N044P031N013(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='1' AND A( 3)='0' )then
          cVar1S25S103N015N044P031N013(0) <='1';
          else
          cVar1S25S103N015N044P031N013(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='1' )then
          cVar1S26S103N015N044N031P030(0) <='1';
          else
          cVar1S26S103N015N044N031P030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='1' )then
          cVar1S27S103N015N044N031P030(0) <='1';
          else
          cVar1S27S103N015N044N031P030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='1' )then
          cVar1S28S103N015N044N031P030(0) <='1';
          else
          cVar1S28S103N015N044N031P030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='1' )then
          cVar1S29S103N015N044N031P030(0) <='1';
          else
          cVar1S29S103N015N044N031P030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='0' )then
          cVar1S30S103N015N044N031N030(0) <='1';
          else
          cVar1S30S103N015N044N031N030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='0' )then
          cVar1S31S103N015N044N031N030(0) <='1';
          else
          cVar1S31S103N015N044N031N030(0) <='0';
          end if;
        if(A( 2)='0' AND D( 6)='0' AND B( 4)='0' AND B(14)='0' )then
          cVar1S32S103N015N044N031N030(0) <='1';
          else
          cVar1S32S103N015N044N031N030(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='1' AND D( 2)='0' AND B(15)='0' )then
          cVar1S0S104P015P005P060P028(0) <='1';
          else
          cVar1S0S104P015P005P060P028(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='1' AND D( 2)='0' AND B(15)='0' )then
          cVar1S1S104P015P005P060P028(0) <='1';
          else
          cVar1S1S104P015P005P060P028(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='1' AND D( 2)='0' AND B(15)='1' )then
          cVar1S2S104P015P005P060P028(0) <='1';
          else
          cVar1S2S104P015P005P060P028(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='1' AND D( 2)='1' AND A( 1)='1' )then
          cVar1S3S104P015P005P060P017nsss(0) <='1';
          else
          cVar1S3S104P015P005P060P017nsss(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='1' AND D( 4)='1' )then
          cVar1S4S104P015N005P063P052(0) <='1';
          else
          cVar1S4S104P015N005P063P052(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='1' AND D( 4)='0' )then
          cVar1S5S104P015N005P063N052(0) <='1';
          else
          cVar1S5S104P015N005P063N052(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='1' AND D( 4)='0' )then
          cVar1S6S104P015N005P063N052(0) <='1';
          else
          cVar1S6S104P015N005P063N052(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='1' AND D( 4)='0' )then
          cVar1S7S104P015N005P063N052(0) <='1';
          else
          cVar1S7S104P015N005P063N052(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='0' )then
          cVar1S8S104P015N005N063P017(0) <='1';
          else
          cVar1S8S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='0' )then
          cVar1S9S104P015N005N063P017(0) <='1';
          else
          cVar1S9S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='0' )then
          cVar1S10S104P015N005N063P017(0) <='1';
          else
          cVar1S10S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='1' )then
          cVar1S11S104P015N005N063P017(0) <='1';
          else
          cVar1S11S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='1' )then
          cVar1S12S104P015N005N063P017(0) <='1';
          else
          cVar1S12S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='1' )then
          cVar1S13S104P015N005N063P017(0) <='1';
          else
          cVar1S13S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='0' AND A( 7)='0' AND E(10)='0' AND A( 1)='1' )then
          cVar1S14S104P015N005N063P017(0) <='1';
          else
          cVar1S14S104P015N005N063P017(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='1' AND D( 2)='0' AND D( 9)='0' )then
          cVar1S15S104P015P029P060P065(0) <='1';
          else
          cVar1S15S104P015P029P060P065(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='1' AND D( 2)='0' AND D( 9)='0' )then
          cVar1S16S104P015P029P060P065(0) <='1';
          else
          cVar1S16S104P015P029P060P065(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='1' AND D( 2)='0' AND D( 9)='0' )then
          cVar1S17S104P015P029P060P065(0) <='1';
          else
          cVar1S17S104P015P029P060P065(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='0' AND A( 5)='0' )then
          cVar1S18S104P015N029P056P009(0) <='1';
          else
          cVar1S18S104P015N029P056P009(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='0' AND A( 5)='0' )then
          cVar1S19S104P015N029P056P009(0) <='1';
          else
          cVar1S19S104P015N029P056P009(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='0' AND A( 5)='0' )then
          cVar1S20S104P015N029P056P009(0) <='1';
          else
          cVar1S20S104P015N029P056P009(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='0' AND A( 5)='1' )then
          cVar1S21S104P015N029P056P009(0) <='1';
          else
          cVar1S21S104P015N029P056P009(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='0' AND A( 5)='1' )then
          cVar1S22S104P015N029P056P009(0) <='1';
          else
          cVar1S22S104P015N029P056P009(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='1' AND B( 4)='1' )then
          cVar1S23S104P015N029P056P031(0) <='1';
          else
          cVar1S23S104P015N029P056P031(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='1' AND B( 4)='0' )then
          cVar1S24S104P015N029P056N031(0) <='1';
          else
          cVar1S24S104P015N029P056N031(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='1' AND B( 4)='0' )then
          cVar1S25S104P015N029P056N031(0) <='1';
          else
          cVar1S25S104P015N029P056N031(0) <='0';
          end if;
        if(A( 2)='1' AND B( 5)='0' AND D( 3)='1' AND B( 4)='0' )then
          cVar1S26S104P015N029P056N031(0) <='1';
          else
          cVar1S26S104P015N029P056N031(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar1S0S105P017P015P018P013(0) <='1';
          else
          cVar1S0S105P017P015P018P013(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='0' AND A( 3)='0' )then
          cVar1S1S105P017P015P018P013(0) <='1';
          else
          cVar1S1S105P017P015P018P013(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S2S105P017P015P018P013(0) <='1';
          else
          cVar1S2S105P017P015P018P013(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S3S105P017P015P018P013(0) <='1';
          else
          cVar1S3S105P017P015P018P013(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar1S4S105P017P015P018P013(0) <='1';
          else
          cVar1S4S105P017P015P018P013(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='1' AND D( 2)='1' )then
          cVar1S5S105P017P015P018P060nsss(0) <='1';
          else
          cVar1S5S105P017P015P018P060nsss(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S6S105P017P015P018N060(0) <='1';
          else
          cVar1S6S105P017P015P018N060(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='0' AND A(10)='1' AND D( 2)='0' )then
          cVar1S7S105P017P015P018N060(0) <='1';
          else
          cVar1S7S105P017P015P018N060(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S8S105P017P015P058P048(0) <='1';
          else
          cVar1S8S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S9S105P017P015P058P048(0) <='1';
          else
          cVar1S9S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S10S105P017P015P058P048(0) <='1';
          else
          cVar1S10S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='0' )then
          cVar1S11S105P017P015P058P048(0) <='1';
          else
          cVar1S11S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='1' )then
          cVar1S12S105P017P015P058P048(0) <='1';
          else
          cVar1S12S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='0' AND D( 5)='1' )then
          cVar1S13S105P017P015P058P048(0) <='1';
          else
          cVar1S13S105P017P015P058P048(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='1' AND B( 2)='0' )then
          cVar1S14S105P017P015P058P035(0) <='1';
          else
          cVar1S14S105P017P015P058P035(0) <='0';
          end if;
        if(A( 1)='1' AND A( 2)='1' AND E( 3)='1' AND B( 2)='0' )then
          cVar1S15S105P017P015P058P035(0) <='1';
          else
          cVar1S15S105P017P015P058P035(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S16S105N017P015P034P014(0) <='1';
          else
          cVar1S16S105N017P015P034P014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S17S105N017P015P034P014(0) <='1';
          else
          cVar1S17S105N017P015P034P014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S18S105N017P015P034P014(0) <='1';
          else
          cVar1S18S105N017P015P034P014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S19S105N017P015P034N014(0) <='1';
          else
          cVar1S19S105N017P015P034N014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S20S105N017P015P034N014(0) <='1';
          else
          cVar1S20S105N017P015P034N014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S21S105N017P015P034N014(0) <='1';
          else
          cVar1S21S105N017P015P034N014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S22S105N017P015P034N014(0) <='1';
          else
          cVar1S22S105N017P015P034N014(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='0' )then
          cVar1S23S105N017P015N034P065(0) <='1';
          else
          cVar1S23S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='0' )then
          cVar1S24S105N017P015N034P065(0) <='1';
          else
          cVar1S24S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='0' )then
          cVar1S25S105N017P015N034P065(0) <='1';
          else
          cVar1S25S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='1' )then
          cVar1S26S105N017P015N034P065(0) <='1';
          else
          cVar1S26S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='1' )then
          cVar1S27S105N017P015N034P065(0) <='1';
          else
          cVar1S27S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='0' AND B(12)='0' AND D( 9)='1' )then
          cVar1S28S105N017P015N034P065(0) <='1';
          else
          cVar1S28S105N017P015N034P065(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='1' AND A(17)='1' )then
          cVar1S29S105N017P015P005P004nsss(0) <='1';
          else
          cVar1S29S105N017P015P005P004nsss(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='1' AND A(17)='0' )then
          cVar1S30S105N017P015P005N004(0) <='1';
          else
          cVar1S30S105N017P015P005N004(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='1' AND A(17)='0' )then
          cVar1S31S105N017P015P005N004(0) <='1';
          else
          cVar1S31S105N017P015P005N004(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='0' )then
          cVar1S32S105N017P015N005P043(0) <='1';
          else
          cVar1S32S105N017P015N005P043(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='0' )then
          cVar1S33S105N017P015N005P043(0) <='1';
          else
          cVar1S33S105N017P015N005P043(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='0' )then
          cVar1S34S105N017P015N005P043(0) <='1';
          else
          cVar1S34S105N017P015N005P043(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='1' )then
          cVar1S35S105N017P015N005P043(0) <='1';
          else
          cVar1S35S105N017P015N005P043(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='1' )then
          cVar1S36S105N017P015N005P043(0) <='1';
          else
          cVar1S36S105N017P015N005P043(0) <='0';
          end if;
        if(A( 1)='0' AND A( 2)='1' AND A( 7)='0' AND E(15)='1' )then
          cVar1S37S105N017P015N005P043(0) <='1';
          else
          cVar1S37S105N017P015N005P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='1' AND B(18)='1' )then
          cVar1S0S106P065P015P045P022(0) <='1';
          else
          cVar1S0S106P065P015P045P022(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S1S106P065P015P045N022(0) <='1';
          else
          cVar1S1S106P065P015P045N022(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='0' )then
          cVar1S2S106P065P015N045P043(0) <='1';
          else
          cVar1S2S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='0' )then
          cVar1S3S106P065P015N045P043(0) <='1';
          else
          cVar1S3S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='0' )then
          cVar1S4S106P065P015N045P043(0) <='1';
          else
          cVar1S4S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='1' )then
          cVar1S5S106P065P015N045P043(0) <='1';
          else
          cVar1S5S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='1' )then
          cVar1S6S106P065P015N045P043(0) <='1';
          else
          cVar1S6S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='0' AND D(14)='0' AND E(15)='1' )then
          cVar1S7S106P065P015N045P043(0) <='1';
          else
          cVar1S7S106P065P015N045P043(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='1' AND D( 2)='0' )then
          cVar1S8S106P065P015P029P060(0) <='1';
          else
          cVar1S8S106P065P015P029P060(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='0' )then
          cVar1S9S106P065P015N029P014(0) <='1';
          else
          cVar1S9S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='0' )then
          cVar1S10S106P065P015N029P014(0) <='1';
          else
          cVar1S10S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='0' )then
          cVar1S11S106P065P015N029P014(0) <='1';
          else
          cVar1S11S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='1' )then
          cVar1S12S106P065P015N029P014(0) <='1';
          else
          cVar1S12S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='1' )then
          cVar1S13S106P065P015N029P014(0) <='1';
          else
          cVar1S13S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='0' AND A( 2)='1' AND B( 5)='0' AND A(12)='1' )then
          cVar1S14S106P065P015N029P014(0) <='1';
          else
          cVar1S14S106P065P015N029P014(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='1' )then
          cVar1S15S106P065P052nsss(0) <='1';
          else
          cVar1S15S106P065P052nsss(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='1' )then
          cVar1S16S106P065N052P035P017(0) <='1';
          else
          cVar1S16S106P065N052P035P017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='1' )then
          cVar1S17S106P065N052P035P017(0) <='1';
          else
          cVar1S17S106P065N052P035P017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='1' )then
          cVar1S18S106P065N052P035P017(0) <='1';
          else
          cVar1S18S106P065N052P035P017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='0' )then
          cVar1S19S106P065N052P035N017(0) <='1';
          else
          cVar1S19S106P065N052P035N017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='0' )then
          cVar1S20S106P065N052P035N017(0) <='1';
          else
          cVar1S20S106P065N052P035N017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='1' AND A( 1)='0' )then
          cVar1S21S106P065N052P035N017(0) <='1';
          else
          cVar1S21S106P065N052P035N017(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='0' AND B(12)='1' )then
          cVar1S22S106P065N052N035P034(0) <='1';
          else
          cVar1S22S106P065N052N035P034(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='0' AND B(12)='1' )then
          cVar1S23S106P065N052N035P034(0) <='1';
          else
          cVar1S23S106P065N052N035P034(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='0' AND B(12)='0' )then
          cVar1S24S106P065N052N035N034(0) <='1';
          else
          cVar1S24S106P065N052N035N034(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='0' AND B(12)='0' )then
          cVar1S25S106P065N052N035N034(0) <='1';
          else
          cVar1S25S106P065N052N035N034(0) <='0';
          end if;
        if(D( 9)='1' AND D( 4)='0' AND B( 2)='0' AND B(12)='0' )then
          cVar1S26S106P065N052N035N034(0) <='1';
          else
          cVar1S26S106P065N052N035N034(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='1' )then
          cVar1S0S107P052P065nsss(0) <='1';
          else
          cVar1S0S107P052P065nsss(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='1' AND A( 5)='0' )then
          cVar1S1S107P052N065P010P009(0) <='1';
          else
          cVar1S1S107P052N065P010P009(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='1' AND A( 5)='0' )then
          cVar1S2S107P052N065P010P009(0) <='1';
          else
          cVar1S2S107P052N065P010P009(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='1' )then
          cVar1S3S107P052N065N010P067(0) <='1';
          else
          cVar1S3S107P052N065N010P067(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='1' )then
          cVar1S4S107P052N065N010P067(0) <='1';
          else
          cVar1S4S107P052N065N010P067(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='0' )then
          cVar1S5S107P052N065N010N067(0) <='1';
          else
          cVar1S5S107P052N065N010N067(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='0' )then
          cVar1S6S107P052N065N010N067(0) <='1';
          else
          cVar1S6S107P052N065N010N067(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='0' )then
          cVar1S7S107P052N065N010N067(0) <='1';
          else
          cVar1S7S107P052N065N010N067(0) <='0';
          end if;
        if(D( 4)='1' AND D( 9)='0' AND A(14)='0' AND E( 9)='0' )then
          cVar1S8S107P052N065N010N067(0) <='1';
          else
          cVar1S8S107P052N065N010N067(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='1' AND A( 7)='1' )then
          cVar1S9S107N052P044P025P005nsss(0) <='1';
          else
          cVar1S9S107N052P044P025P005nsss(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='1' AND A( 7)='0' )then
          cVar1S10S107N052P044P025N005(0) <='1';
          else
          cVar1S10S107N052P044P025N005(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='1' AND A( 7)='0' )then
          cVar1S11S107N052P044P025N005(0) <='1';
          else
          cVar1S11S107N052P044P025N005(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='0' AND E( 9)='1' )then
          cVar1S12S107N052P044N025P067nsss(0) <='1';
          else
          cVar1S12S107N052P044N025P067nsss(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='0' AND E( 9)='0' )then
          cVar1S13S107N052P044N025N067(0) <='1';
          else
          cVar1S13S107N052P044N025N067(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='0' AND E( 9)='0' )then
          cVar1S14S107N052P044N025N067(0) <='1';
          else
          cVar1S14S107N052P044N025N067(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='1' AND B( 7)='0' AND E( 9)='0' )then
          cVar1S15S107N052P044N025N067(0) <='1';
          else
          cVar1S15S107N052P044N025N067(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S16S107N052N044P058P033(0) <='1';
          else
          cVar1S16S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S17S107N052N044P058P033(0) <='1';
          else
          cVar1S17S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='0' AND B( 3)='0' )then
          cVar1S18S107N052N044P058P033(0) <='1';
          else
          cVar1S18S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='0' AND B( 3)='1' )then
          cVar1S19S107N052N044P058P033(0) <='1';
          else
          cVar1S19S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='1' )then
          cVar1S20S107N052N044P058P033(0) <='1';
          else
          cVar1S20S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='1' )then
          cVar1S21S107N052N044P058P033(0) <='1';
          else
          cVar1S21S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='1' )then
          cVar1S22S107N052N044P058P033(0) <='1';
          else
          cVar1S22S107N052N044P058P033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S23S107N052N044P058N033(0) <='1';
          else
          cVar1S23S107N052N044P058N033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S24S107N052N044P058N033(0) <='1';
          else
          cVar1S24S107N052N044P058N033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S25S107N052N044P058N033(0) <='1';
          else
          cVar1S25S107N052N044P058N033(0) <='0';
          end if;
        if(D( 4)='0' AND D( 6)='0' AND E( 3)='1' AND B( 3)='0' )then
          cVar1S26S107N052N044P058N033(0) <='1';
          else
          cVar1S26S107N052N044P058N033(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='1' )then
          cVar1S0S108P058P033P060P006(0) <='1';
          else
          cVar1S0S108P058P033P060P006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='1' )then
          cVar1S1S108P058P033P060P006(0) <='1';
          else
          cVar1S1S108P058P033P060P006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='1' )then
          cVar1S2S108P058P033P060P006(0) <='1';
          else
          cVar1S2S108P058P033P060P006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='0' )then
          cVar1S3S108P058P033P060N006(0) <='1';
          else
          cVar1S3S108P058P033P060N006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='0' )then
          cVar1S4S108P058P033P060N006(0) <='1';
          else
          cVar1S4S108P058P033P060N006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='0' AND A(16)='0' )then
          cVar1S5S108P058P033P060N006(0) <='1';
          else
          cVar1S5S108P058P033P060N006(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='1' AND E( 1)='1' )then
          cVar1S6S108P058P033P060P066(0) <='1';
          else
          cVar1S6S108P058P033P060P066(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='1' AND E( 1)='1' )then
          cVar1S7S108P058P033P060P066(0) <='1';
          else
          cVar1S7S108P058P033P060P066(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='1' AND E( 1)='0' )then
          cVar1S8S108P058P033P060N066(0) <='1';
          else
          cVar1S8S108P058P033P060N066(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='1' AND E( 1)='0' )then
          cVar1S9S108P058P033P060N066(0) <='1';
          else
          cVar1S9S108P058P033P060N066(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='0' AND D( 2)='1' AND E( 1)='0' )then
          cVar1S10S108P058P033P060N066(0) <='1';
          else
          cVar1S10S108P058P033P060N066(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='1' AND A(16)='0' AND E(13)='0' )then
          cVar1S11S108P058P033P006P051(0) <='1';
          else
          cVar1S11S108P058P033P006P051(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='1' AND A(16)='0' AND E(13)='0' )then
          cVar1S12S108P058P033P006P051(0) <='1';
          else
          cVar1S12S108P058P033P006P051(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='1' AND A(16)='0' AND E(13)='0' )then
          cVar1S13S108P058P033P006P051(0) <='1';
          else
          cVar1S13S108P058P033P006P051(0) <='0';
          end if;
        if(E( 3)='0' AND B( 3)='1' AND A(16)='1' AND A( 1)='0' )then
          cVar1S14S108P058P033P006P017(0) <='1';
          else
          cVar1S14S108P058P033P006P017(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='1' AND B( 3)='1' )then
          cVar1S15S108P058P006P013P033(0) <='1';
          else
          cVar1S15S108P058P006P013P033(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='1' AND B( 3)='1' )then
          cVar1S16S108P058P006P013P033(0) <='1';
          else
          cVar1S16S108P058P006P013P033(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='1' AND B( 3)='0' )then
          cVar1S17S108P058P006P013N033(0) <='1';
          else
          cVar1S17S108P058P006P013N033(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='1' AND B( 3)='0' )then
          cVar1S18S108P058P006P013N033(0) <='1';
          else
          cVar1S18S108P058P006P013N033(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='1' AND B( 3)='0' )then
          cVar1S19S108P058P006P013N033(0) <='1';
          else
          cVar1S19S108P058P006P013N033(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='0' AND A(12)='1' )then
          cVar1S20S108P058P006N013P014(0) <='1';
          else
          cVar1S20S108P058P006N013P014(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='0' AND A(12)='1' )then
          cVar1S21S108P058P006N013P014(0) <='1';
          else
          cVar1S21S108P058P006N013P014(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='0' AND A(12)='0' )then
          cVar1S22S108P058P006N013N014(0) <='1';
          else
          cVar1S22S108P058P006N013N014(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='0' AND A(12)='0' )then
          cVar1S23S108P058P006N013N014(0) <='1';
          else
          cVar1S23S108P058P006N013N014(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='0' AND A( 3)='0' AND A(12)='0' )then
          cVar1S24S108P058P006N013N014(0) <='1';
          else
          cVar1S24S108P058P006N013N014(0) <='0';
          end if;
        if(E( 3)='1' AND A(16)='1' AND A( 1)='1' )then
          cVar1S25S108P058P006P017nsss(0) <='1';
          else
          cVar1S25S108P058P006P017nsss(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='1' AND A(11)='0' AND A(10)='0' )then
          cVar1S0S109P045P004P016P018nsss(0) <='1';
          else
          cVar1S0S109P045P004P016P018nsss(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='1' AND B(17)='1' )then
          cVar1S1S109P045N004P006P024nsss(0) <='1';
          else
          cVar1S1S109P045N004P006P024nsss(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='1' AND B(17)='0' )then
          cVar1S2S109P045N004P006N024(0) <='1';
          else
          cVar1S2S109P045N004P006N024(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='0' AND B( 8)='1' )then
          cVar1S3S109P045N004N006P023nsss(0) <='1';
          else
          cVar1S3S109P045N004N006P023nsss(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='0' AND B( 8)='0' )then
          cVar1S4S109P045N004N006N023(0) <='1';
          else
          cVar1S4S109P045N004N006N023(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='0' AND B( 8)='0' )then
          cVar1S5S109P045N004N006N023(0) <='1';
          else
          cVar1S5S109P045N004N006N023(0) <='0';
          end if;
        if(D(14)='1' AND A(17)='0' AND A(16)='0' AND B( 8)='0' )then
          cVar1S6S109P045N004N006N023(0) <='1';
          else
          cVar1S6S109P045N004N006N023(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='1' AND E( 4)='1' )then
          cVar1S7S109N045P029P011P054(0) <='1';
          else
          cVar1S7S109N045P029P011P054(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='1' AND E( 4)='1' )then
          cVar1S8S109N045P029P011P054(0) <='1';
          else
          cVar1S8S109N045P029P011P054(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='1' AND E( 4)='0' )then
          cVar1S9S109N045P029P011N054(0) <='1';
          else
          cVar1S9S109N045P029P011N054(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='1' AND E( 4)='0' )then
          cVar1S10S109N045P029P011N054(0) <='1';
          else
          cVar1S10S109N045P029P011N054(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='1' AND E( 4)='0' )then
          cVar1S11S109N045P029P011N054(0) <='1';
          else
          cVar1S11S109N045P029P011N054(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='0' AND A(14)='1' )then
          cVar1S12S109N045P029N011P010(0) <='1';
          else
          cVar1S12S109N045P029N011P010(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='0' AND A(14)='1' )then
          cVar1S13S109N045P029N011P010(0) <='1';
          else
          cVar1S13S109N045P029N011P010(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='0' AND A(14)='0' )then
          cVar1S14S109N045P029N011N010(0) <='1';
          else
          cVar1S14S109N045P029N011N010(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='0' AND A(14)='0' )then
          cVar1S15S109N045P029N011N010(0) <='1';
          else
          cVar1S15S109N045P029N011N010(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='1' AND A( 4)='0' AND A(14)='0' )then
          cVar1S16S109N045P029N011N010(0) <='1';
          else
          cVar1S16S109N045P029N011N010(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='1' )then
          cVar1S17S109N045N029P011P007(0) <='1';
          else
          cVar1S17S109N045N029P011P007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='1' )then
          cVar1S18S109N045N029P011P007(0) <='1';
          else
          cVar1S18S109N045N029P011P007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='1' )then
          cVar1S19S109N045N029P011P007(0) <='1';
          else
          cVar1S19S109N045N029P011P007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='0' )then
          cVar1S20S109N045N029P011N007(0) <='1';
          else
          cVar1S20S109N045N029P011N007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='0' )then
          cVar1S21S109N045N029P011N007(0) <='1';
          else
          cVar1S21S109N045N029P011N007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='0' AND A( 6)='0' )then
          cVar1S22S109N045N029P011N007(0) <='1';
          else
          cVar1S22S109N045N029P011N007(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='0' )then
          cVar1S23S109N045N029P011P069(0) <='1';
          else
          cVar1S23S109N045N029P011P069(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='0' )then
          cVar1S24S109N045N029P011P069(0) <='1';
          else
          cVar1S24S109N045N029P011P069(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='0' )then
          cVar1S25S109N045N029P011P069(0) <='1';
          else
          cVar1S25S109N045N029P011P069(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='0' )then
          cVar1S26S109N045N029P011P069(0) <='1';
          else
          cVar1S26S109N045N029P011P069(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='1' )then
          cVar1S27S109N045N029P011P069(0) <='1';
          else
          cVar1S27S109N045N029P011P069(0) <='0';
          end if;
        if(D(14)='0' AND B( 5)='0' AND A( 4)='1' AND D( 8)='1' )then
          cVar1S28S109N045N029P011P069(0) <='1';
          else
          cVar1S28S109N045N029P011P069(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S0S110P011P029P007P025(0) <='1';
          else
          cVar1S0S110P011P029P007P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S1S110P011P029P007P025(0) <='1';
          else
          cVar1S1S110P011P029P007P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S2S110P011P029P007P025(0) <='1';
          else
          cVar1S2S110P011P029P007P025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S3S110P011P029P007N025(0) <='1';
          else
          cVar1S3S110P011P029P007N025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S4S110P011P029P007N025(0) <='1';
          else
          cVar1S4S110P011P029P007N025(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='0' )then
          cVar1S5S110P011P029N007P049(0) <='1';
          else
          cVar1S5S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='0' )then
          cVar1S6S110P011P029N007P049(0) <='1';
          else
          cVar1S6S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='0' )then
          cVar1S7S110P011P029N007P049(0) <='1';
          else
          cVar1S7S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='0' )then
          cVar1S8S110P011P029N007P049(0) <='1';
          else
          cVar1S8S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='1' )then
          cVar1S9S110P011P029N007P049(0) <='1';
          else
          cVar1S9S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='1' )then
          cVar1S10S110P011P029N007P049(0) <='1';
          else
          cVar1S10S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='1' )then
          cVar1S11S110P011P029N007P049(0) <='1';
          else
          cVar1S11S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='0' AND A( 6)='0' AND D(13)='1' )then
          cVar1S12S110P011P029N007P049(0) <='1';
          else
          cVar1S12S110P011P029N007P049(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A( 7)='0' AND A(14)='1' )then
          cVar1S13S110P011P029P005P010(0) <='1';
          else
          cVar1S13S110P011P029P005P010(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A( 7)='0' AND A(14)='1' )then
          cVar1S14S110P011P029P005P010(0) <='1';
          else
          cVar1S14S110P011P029P005P010(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A( 7)='0' AND A(14)='0' )then
          cVar1S15S110P011P029P005N010(0) <='1';
          else
          cVar1S15S110P011P029P005N010(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A( 7)='0' AND A(14)='0' )then
          cVar1S16S110P011P029P005N010(0) <='1';
          else
          cVar1S16S110P011P029P005N010(0) <='0';
          end if;
        if(A( 4)='0' AND B( 5)='1' AND A( 7)='0' AND A(14)='0' )then
          cVar1S17S110P011P029P005N010(0) <='1';
          else
          cVar1S17S110P011P029P005N010(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND E( 4)='1' AND D(11)='0' )then
          cVar1S18S110P011P029P054P057(0) <='1';
          else
          cVar1S18S110P011P029P054P057(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND E( 4)='1' AND D(11)='0' )then
          cVar1S19S110P011P029P054P057(0) <='1';
          else
          cVar1S19S110P011P029P054P057(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND E( 4)='0' AND D(12)='1' )then
          cVar1S20S110P011P029N054P053nsss(0) <='1';
          else
          cVar1S20S110P011P029N054P053nsss(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND E( 4)='0' AND D(12)='0' )then
          cVar1S21S110P011P029N054N053(0) <='1';
          else
          cVar1S21S110P011P029N054N053(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='1' AND E( 4)='0' AND D(12)='0' )then
          cVar1S22S110P011P029N054N053(0) <='1';
          else
          cVar1S22S110P011P029N054N053(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='0' )then
          cVar1S23S110P011N029P069P030(0) <='1';
          else
          cVar1S23S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='0' )then
          cVar1S24S110P011N029P069P030(0) <='1';
          else
          cVar1S24S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='0' )then
          cVar1S25S110P011N029P069P030(0) <='1';
          else
          cVar1S25S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='0' )then
          cVar1S26S110P011N029P069P030(0) <='1';
          else
          cVar1S26S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='1' )then
          cVar1S27S110P011N029P069P030(0) <='1';
          else
          cVar1S27S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='0' AND B(14)='1' )then
          cVar1S28S110P011N029P069P030(0) <='1';
          else
          cVar1S28S110P011N029P069P030(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='1' AND D( 0)='1' )then
          cVar1S29S110P011N029P069P068(0) <='1';
          else
          cVar1S29S110P011N029P069P068(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='1' AND D( 0)='1' )then
          cVar1S30S110P011N029P069P068(0) <='1';
          else
          cVar1S30S110P011N029P069P068(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S31S110P011N029P069N068(0) <='1';
          else
          cVar1S31S110P011N029P069N068(0) <='0';
          end if;
        if(A( 4)='1' AND B( 5)='0' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S32S110P011N029P069N068(0) <='1';
          else
          cVar1S32S110P011N029P069N068(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND B( 7)='1' )then
          cVar1S0S111P009P049P025nsss(0) <='1';
          else
          cVar1S0S111P009P049P025nsss(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND B( 7)='0' AND E( 9)='0' )then
          cVar1S1S111P009P049N025P067(0) <='1';
          else
          cVar1S1S111P009P049N025P067(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='1' AND B( 5)='1' )then
          cVar1S2S111P009N049P053P029nsss(0) <='1';
          else
          cVar1S2S111P009N049P053P029nsss(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='1' AND B( 5)='0' )then
          cVar1S3S111P009N049P053N029(0) <='1';
          else
          cVar1S3S111P009N049P053N029(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S4S111P009N049N053P050(0) <='1';
          else
          cVar1S4S111P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S5S111P009N049N053P050(0) <='1';
          else
          cVar1S5S111P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='1' )then
          cVar1S6S111P009N049N053P050(0) <='1';
          else
          cVar1S6S111P009N049N053P050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S7S111P009N049N053N050(0) <='1';
          else
          cVar1S7S111P009N049N053N050(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND D(12)='0' AND E( 5)='0' )then
          cVar1S8S111P009N049N053N050(0) <='1';
          else
          cVar1S8S111P009N049N053N050(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='1' AND A(17)='1' )then
          cVar1S9S111N009P044P004nsss(0) <='1';
          else
          cVar1S9S111N009P044P004nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='1' AND A(17)='0' AND E(13)='1' )then
          cVar1S10S111N009P044N004P051nsss(0) <='1';
          else
          cVar1S10S111N009P044N004P051nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='1' AND A(17)='0' AND E(13)='0' )then
          cVar1S11S111N009P044N004N051(0) <='1';
          else
          cVar1S11S111N009P044N004N051(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='1' AND A(17)='0' AND E(13)='0' )then
          cVar1S12S111N009P044N004N051(0) <='1';
          else
          cVar1S12S111N009P044N004N051(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='1' AND A(17)='0' AND E(13)='0' )then
          cVar1S13S111N009P044N004N051(0) <='1';
          else
          cVar1S13S111N009P044N004N051(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='0' AND B( 8)='0' )then
          cVar1S14S111N009N044P042P023(0) <='1';
          else
          cVar1S14S111N009N044P042P023(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='0' AND B( 8)='0' )then
          cVar1S15S111N009N044P042P023(0) <='1';
          else
          cVar1S15S111N009N044P042P023(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='0' AND B( 8)='1' )then
          cVar1S16S111N009N044P042P023(0) <='1';
          else
          cVar1S16S111N009N044P042P023(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='0' AND B( 8)='1' )then
          cVar1S17S111N009N044P042P023(0) <='1';
          else
          cVar1S17S111N009N044P042P023(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='1' )then
          cVar1S18S111N009N044P042P058nsss(0) <='1';
          else
          cVar1S18S111N009N044P042P058nsss(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='0' )then
          cVar1S19S111N009N044P042N058(0) <='1';
          else
          cVar1S19S111N009N044P042N058(0) <='0';
          end if;
        if(A( 5)='0' AND D( 6)='0' AND E( 7)='1' AND E( 3)='0' )then
          cVar1S20S111N009N044P042N058(0) <='1';
          else
          cVar1S20S111N009N044P042N058(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND B( 7)='1' )then
          cVar1S0S112P009P049P025nsss(0) <='1';
          else
          cVar1S0S112P009P049P025nsss(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='1' AND B( 7)='0' AND E( 9)='0' )then
          cVar1S1S112P009P049N025P067(0) <='1';
          else
          cVar1S1S112P009P049N025P067(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='1' AND B( 6)='1' )then
          cVar1S2S112P009N049P050P027(0) <='1';
          else
          cVar1S2S112P009N049P050P027(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S3S112P009N049P050N027(0) <='1';
          else
          cVar1S3S112P009N049P050N027(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S4S112P009N049P050N027(0) <='1';
          else
          cVar1S4S112P009N049P050N027(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='1' AND B( 6)='0' )then
          cVar1S5S112P009N049P050N027(0) <='1';
          else
          cVar1S5S112P009N049P050N027(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='0' AND D(12)='1' )then
          cVar1S6S112P009N049N050P053(0) <='1';
          else
          cVar1S6S112P009N049N050P053(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='0' AND D(12)='1' )then
          cVar1S7S112P009N049N050P053(0) <='1';
          else
          cVar1S7S112P009N049N050P053(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='0' AND D(12)='1' )then
          cVar1S8S112P009N049N050P053(0) <='1';
          else
          cVar1S8S112P009N049N050P053(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='0' AND D(12)='0' )then
          cVar1S9S112P009N049N050N053(0) <='1';
          else
          cVar1S9S112P009N049N050N053(0) <='0';
          end if;
        if(A( 5)='1' AND D(13)='0' AND E( 5)='0' AND D(12)='0' )then
          cVar1S10S112P009N049N050N053(0) <='1';
          else
          cVar1S10S112P009N049N050N053(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='0' AND D( 1)='1' )then
          cVar1S11S112N009P011P053P064(0) <='1';
          else
          cVar1S11S112N009P011P053P064(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='0' AND D( 1)='1' )then
          cVar1S12S112N009P011P053P064(0) <='1';
          else
          cVar1S12S112N009P011P053P064(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='0' AND D( 1)='1' )then
          cVar1S13S112N009P011P053P064(0) <='1';
          else
          cVar1S13S112N009P011P053P064(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='0' AND D( 1)='0' )then
          cVar1S14S112N009P011P053N064(0) <='1';
          else
          cVar1S14S112N009P011P053N064(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='0' AND D( 1)='0' )then
          cVar1S15S112N009P011P053N064(0) <='1';
          else
          cVar1S15S112N009P011P053N064(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='1' AND B(11)='0' )then
          cVar1S16S112N009P011P053P036(0) <='1';
          else
          cVar1S16S112N009P011P053P036(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='1' AND B(11)='0' )then
          cVar1S17S112N009P011P053P036(0) <='1';
          else
          cVar1S17S112N009P011P053P036(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='1' AND B(11)='0' )then
          cVar1S18S112N009P011P053P036(0) <='1';
          else
          cVar1S18S112N009P011P053P036(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='0' AND D(12)='1' AND B(11)='1' )then
          cVar1S19S112N009P011P053P036(0) <='1';
          else
          cVar1S19S112N009P011P053P036(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='1' AND E( 4)='1' )then
          cVar1S20S112N009P011P029P054(0) <='1';
          else
          cVar1S20S112N009P011P029P054(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='1' AND E( 4)='1' )then
          cVar1S21S112N009P011P029P054(0) <='1';
          else
          cVar1S21S112N009P011P029P054(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='1' AND E( 4)='0' )then
          cVar1S22S112N009P011P029N054(0) <='1';
          else
          cVar1S22S112N009P011P029N054(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='1' AND E( 4)='0' )then
          cVar1S23S112N009P011P029N054(0) <='1';
          else
          cVar1S23S112N009P011P029N054(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='1' AND E( 4)='0' )then
          cVar1S24S112N009P011P029N054(0) <='1';
          else
          cVar1S24S112N009P011P029N054(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='1' )then
          cVar1S25S112N009P011N029P047(0) <='1';
          else
          cVar1S25S112N009P011N029P047(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='1' )then
          cVar1S26S112N009P011N029P047(0) <='1';
          else
          cVar1S26S112N009P011N029P047(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='1' )then
          cVar1S27S112N009P011N029P047(0) <='1';
          else
          cVar1S27S112N009P011N029P047(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='0' )then
          cVar1S28S112N009P011N029N047(0) <='1';
          else
          cVar1S28S112N009P011N029N047(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='0' )then
          cVar1S29S112N009P011N029N047(0) <='1';
          else
          cVar1S29S112N009P011N029N047(0) <='0';
          end if;
        if(A( 5)='0' AND A( 4)='1' AND B( 5)='0' AND E(14)='0' )then
          cVar1S30S112N009P011N029N047(0) <='1';
          else
          cVar1S30S112N009P011N029N047(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND B( 6)='0' AND E(14)='1' )then
          cVar1S0S113P037P066P027P047nsss(0) <='1';
          else
          cVar1S0S113P037P066P027P047nsss(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND B( 6)='0' AND E(14)='0' )then
          cVar1S1S113P037P066P027N047(0) <='1';
          else
          cVar1S1S113P037P066P027N047(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND B( 6)='0' AND E(14)='0' )then
          cVar1S2S113P037P066P027N047(0) <='1';
          else
          cVar1S2S113P037P066P027N047(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='1' AND B( 6)='1' AND D( 0)='1' )then
          cVar1S3S113P037P066P027P068(0) <='1';
          else
          cVar1S3S113P037P066P027P068(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S4S113P037N066P069P068(0) <='1';
          else
          cVar1S4S113P037N066P069P068(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='1' AND D( 0)='0' )then
          cVar1S5S113P037N066P069P068(0) <='1';
          else
          cVar1S5S113P037N066P069P068(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='0' AND B( 2)='1' )then
          cVar1S6S113P037N066N069P035(0) <='1';
          else
          cVar1S6S113P037N066N069P035(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='0' AND B( 2)='1' )then
          cVar1S7S113P037N066N069P035(0) <='1';
          else
          cVar1S7S113P037N066N069P035(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='0' AND B( 2)='0' )then
          cVar1S8S113P037N066N069N035(0) <='1';
          else
          cVar1S8S113P037N066N069N035(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='0' AND B( 2)='0' )then
          cVar1S9S113P037N066N069N035(0) <='1';
          else
          cVar1S9S113P037N066N069N035(0) <='0';
          end if;
        if(B( 1)='1' AND E( 1)='0' AND D( 8)='0' AND B( 2)='0' )then
          cVar1S10S113P037N066N069N035(0) <='1';
          else
          cVar1S10S113P037N066N069N035(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='1' AND E(15)='1' )then
          cVar1S11S113N037P059P043nsss(0) <='1';
          else
          cVar1S11S113N037P059P043nsss(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='1' AND E(15)='0' AND E( 3)='0' )then
          cVar1S12S113N037P059N043P058(0) <='1';
          else
          cVar1S12S113N037P059N043P058(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='1' AND E(15)='0' AND E( 3)='1' )then
          cVar1S13S113N037P059N043P058(0) <='1';
          else
          cVar1S13S113N037P059N043P058(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='1' AND E(15)='0' AND E( 3)='1' )then
          cVar1S14S113N037P059N043P058(0) <='1';
          else
          cVar1S14S113N037P059N043P058(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='1' )then
          cVar1S15S113N037N059P009P049(0) <='1';
          else
          cVar1S15S113N037N059P009P049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='1' )then
          cVar1S16S113N037N059P009P049(0) <='1';
          else
          cVar1S16S113N037N059P009P049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='1' )then
          cVar1S17S113N037N059P009P049(0) <='1';
          else
          cVar1S17S113N037N059P009P049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='0' )then
          cVar1S18S113N037N059P009N049(0) <='1';
          else
          cVar1S18S113N037N059P009N049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='0' )then
          cVar1S19S113N037N059P009N049(0) <='1';
          else
          cVar1S19S113N037N059P009N049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='0' )then
          cVar1S20S113N037N059P009N049(0) <='1';
          else
          cVar1S20S113N037N059P009N049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='1' AND D(13)='0' )then
          cVar1S21S113N037N059P009N049(0) <='1';
          else
          cVar1S21S113N037N059P009N049(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='1' )then
          cVar1S22S113N037N059N009P054(0) <='1';
          else
          cVar1S22S113N037N059N009P054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='1' )then
          cVar1S23S113N037N059N009P054(0) <='1';
          else
          cVar1S23S113N037N059N009P054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='1' )then
          cVar1S24S113N037N059N009P054(0) <='1';
          else
          cVar1S24S113N037N059N009P054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='1' )then
          cVar1S25S113N037N059N009P054(0) <='1';
          else
          cVar1S25S113N037N059N009P054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='0' )then
          cVar1S26S113N037N059N009N054(0) <='1';
          else
          cVar1S26S113N037N059N009N054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='0' )then
          cVar1S27S113N037N059N009N054(0) <='1';
          else
          cVar1S27S113N037N059N009N054(0) <='0';
          end if;
        if(B( 1)='0' AND E(11)='0' AND A( 5)='0' AND E( 4)='0' )then
          cVar1S28S113N037N059N009N054(0) <='1';
          else
          cVar1S28S113N037N059N009N054(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='1' AND E(15)='1' )then
          cVar1S0S114P064P037P005P043(0) <='1';
          else
          cVar1S0S114P064P037P005P043(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='1' AND E(15)='0' )then
          cVar1S1S114P064P037P005N043(0) <='1';
          else
          cVar1S1S114P064P037P005N043(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='1' AND E(15)='0' )then
          cVar1S2S114P064P037P005N043(0) <='1';
          else
          cVar1S2S114P064P037P005N043(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='1' AND E(15)='0' )then
          cVar1S3S114P064P037P005N043(0) <='1';
          else
          cVar1S3S114P064P037P005N043(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='1' )then
          cVar1S4S114P064P037N005P028(0) <='1';
          else
          cVar1S4S114P064P037N005P028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='1' )then
          cVar1S5S114P064P037N005P028(0) <='1';
          else
          cVar1S5S114P064P037N005P028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='1' )then
          cVar1S6S114P064P037N005P028(0) <='1';
          else
          cVar1S6S114P064P037N005P028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='1' )then
          cVar1S7S114P064P037N005P028(0) <='1';
          else
          cVar1S7S114P064P037N005P028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='0' )then
          cVar1S8S114P064P037N005N028(0) <='1';
          else
          cVar1S8S114P064P037N005N028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='0' )then
          cVar1S9S114P064P037N005N028(0) <='1';
          else
          cVar1S9S114P064P037N005N028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='0' )then
          cVar1S10S114P064P037N005N028(0) <='1';
          else
          cVar1S10S114P064P037N005N028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='0' AND A( 7)='0' AND B(15)='0' )then
          cVar1S11S114P064P037N005N028(0) <='1';
          else
          cVar1S11S114P064P037N005N028(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='1' )then
          cVar1S12S114P064P037P061P012(0) <='1';
          else
          cVar1S12S114P064P037P061P012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='1' )then
          cVar1S13S114P064P037P061P012(0) <='1';
          else
          cVar1S13S114P064P037P061P012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='1' )then
          cVar1S14S114P064P037P061P012(0) <='1';
          else
          cVar1S14S114P064P037P061P012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='1' )then
          cVar1S15S114P064P037P061P012(0) <='1';
          else
          cVar1S15S114P064P037P061P012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='0' )then
          cVar1S16S114P064P037P061N012(0) <='1';
          else
          cVar1S16S114P064P037P061N012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='0' AND A(13)='0' )then
          cVar1S17S114P064P037P061N012(0) <='1';
          else
          cVar1S17S114P064P037P061N012(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='1' AND E( 2)='1' )then
          cVar1S18S114P064P037P061P062nsss(0) <='1';
          else
          cVar1S18S114P064P037P061P062nsss(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='1' AND E( 2)='0' )then
          cVar1S19S114P064P037P061N062(0) <='1';
          else
          cVar1S19S114P064P037P061N062(0) <='0';
          end if;
        if(D( 1)='0' AND B( 1)='1' AND D(10)='1' AND E( 2)='0' )then
          cVar1S20S114P064P037P061N062(0) <='1';
          else
          cVar1S20S114P064P037P061N062(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='1' )then
          cVar1S21S114P064P046nsss(0) <='1';
          else
          cVar1S21S114P064P046nsss(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='0' AND E( 7)='1' )then
          cVar1S22S114P064N046P042nsss(0) <='1';
          else
          cVar1S22S114P064N046P042nsss(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='0' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S23S114P064N046N042P003(0) <='1';
          else
          cVar1S23S114P064N046N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='0' AND E( 7)='0' AND A( 8)='0' )then
          cVar1S24S114P064N046N042P003(0) <='1';
          else
          cVar1S24S114P064N046N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='0' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S25S114P064N046N042P003(0) <='1';
          else
          cVar1S25S114P064N046N042P003(0) <='0';
          end if;
        if(D( 1)='1' AND E( 6)='0' AND E( 7)='0' AND A( 8)='1' )then
          cVar1S26S114P064N046N042P003(0) <='1';
          else
          cVar1S26S114P064N046N042P003(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='1' AND B( 3)='0' AND A( 6)='1' )then
          cVar1S0S115P049P026P033P007nsss(0) <='1';
          else
          cVar1S0S115P049P026P033P007nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='1' AND B( 3)='0' AND A( 6)='0' )then
          cVar1S1S115P049P026P033N007(0) <='1';
          else
          cVar1S1S115P049P026P033N007(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='1' AND B( 3)='0' AND A( 6)='0' )then
          cVar1S2S115P049P026P033N007(0) <='1';
          else
          cVar1S2S115P049P026P033N007(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='1' AND A(17)='1' )then
          cVar1S3S115P049N026P024P004nsss(0) <='1';
          else
          cVar1S3S115P049N026P024P004nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S4S115P049N026P024N004(0) <='1';
          else
          cVar1S4S115P049N026P024N004(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S5S115P049N026P024N004(0) <='1';
          else
          cVar1S5S115P049N026P024N004(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S6S115P049N026P024N004(0) <='1';
          else
          cVar1S6S115P049N026P024N004(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='1' )then
          cVar1S7S115P049N026N024P027(0) <='1';
          else
          cVar1S7S115P049N026N024P027(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='1' )then
          cVar1S8S115P049N026N024P027(0) <='1';
          else
          cVar1S8S115P049N026N024P027(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='1' )then
          cVar1S9S115P049N026N024P027(0) <='1';
          else
          cVar1S9S115P049N026N024P027(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='0' )then
          cVar1S10S115P049N026N024N027(0) <='1';
          else
          cVar1S10S115P049N026N024N027(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='0' )then
          cVar1S11S115P049N026N024N027(0) <='1';
          else
          cVar1S11S115P049N026N024N027(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(17)='0' AND B( 6)='0' )then
          cVar1S12S115P049N026N024N027(0) <='1';
          else
          cVar1S12S115P049N026N024N027(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='1' AND D( 9)='1' )then
          cVar1S13S115N049P064P050P065nsss(0) <='1';
          else
          cVar1S13S115N049P064P050P065nsss(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='1' AND D( 9)='0' )then
          cVar1S14S115N049P064P050N065(0) <='1';
          else
          cVar1S14S115N049P064P050N065(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='1' AND D( 9)='0' )then
          cVar1S15S115N049P064P050N065(0) <='1';
          else
          cVar1S15S115N049P064P050N065(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='0' AND A(15)='0' )then
          cVar1S16S115N049P064N050P008(0) <='1';
          else
          cVar1S16S115N049P064N050P008(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='0' AND A(15)='0' )then
          cVar1S17S115N049P064N050P008(0) <='1';
          else
          cVar1S17S115N049P064N050P008(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='0' AND A(15)='0' )then
          cVar1S18S115N049P064N050P008(0) <='1';
          else
          cVar1S18S115N049P064N050P008(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='0' AND A(15)='1' )then
          cVar1S19S115N049P064N050P008(0) <='1';
          else
          cVar1S19S115N049P064N050P008(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='1' AND E( 5)='0' AND A(15)='1' )then
          cVar1S20S115N049P064N050P008(0) <='1';
          else
          cVar1S20S115N049P064N050P008(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='1' )then
          cVar1S21S115N049N064P047P028(0) <='1';
          else
          cVar1S21S115N049N064P047P028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='1' )then
          cVar1S22S115N049N064P047P028(0) <='1';
          else
          cVar1S22S115N049N064P047P028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='1' )then
          cVar1S23S115N049N064P047P028(0) <='1';
          else
          cVar1S23S115N049N064P047P028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='0' )then
          cVar1S24S115N049N064P047N028(0) <='1';
          else
          cVar1S24S115N049N064P047N028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='0' )then
          cVar1S25S115N049N064P047N028(0) <='1';
          else
          cVar1S25S115N049N064P047N028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='0' AND B(15)='0' )then
          cVar1S26S115N049N064P047N028(0) <='1';
          else
          cVar1S26S115N049N064P047N028(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='1' AND D( 8)='1' )then
          cVar1S27S115N049N064P047P069nsss(0) <='1';
          else
          cVar1S27S115N049N064P047P069nsss(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='1' AND D( 8)='0' )then
          cVar1S28S115N049N064P047N069(0) <='1';
          else
          cVar1S28S115N049N064P047N069(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='1' AND D( 8)='0' )then
          cVar1S29S115N049N064P047N069(0) <='1';
          else
          cVar1S29S115N049N064P047N069(0) <='0';
          end if;
        if(D(13)='0' AND D( 1)='0' AND E(14)='1' AND D( 8)='0' )then
          cVar1S30S115N049N064P047N069(0) <='1';
          else
          cVar1S30S115N049N064P047N069(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S0S116P060P062P049P024(0) <='1';
          else
          cVar1S0S116P060P062P049P024(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S1S116P060P062P049P024(0) <='1';
          else
          cVar1S1S116P060P062P049P024(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S2S116P060P062P049P024(0) <='1';
          else
          cVar1S2S116P060P062P049P024(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S3S116P060P062P049N024(0) <='1';
          else
          cVar1S3S116P060P062P049N024(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S4S116P060P062P049N024(0) <='1';
          else
          cVar1S4S116P060P062P049N024(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S5S116P060P062N049P047(0) <='1';
          else
          cVar1S5S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S6S116P060P062N049P047(0) <='1';
          else
          cVar1S6S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S7S116P060P062N049P047(0) <='1';
          else
          cVar1S7S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='1' )then
          cVar1S8S116P060P062N049P047(0) <='1';
          else
          cVar1S8S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='1' )then
          cVar1S9S116P060P062N049P047(0) <='1';
          else
          cVar1S9S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='0' AND D(13)='0' AND E(14)='1' )then
          cVar1S10S116P060P062N049P047(0) <='1';
          else
          cVar1S10S116P060P062N049P047(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='1' AND A(12)='0' )then
          cVar1S11S116P060P062P050P014nsss(0) <='1';
          else
          cVar1S11S116P060P062P050P014nsss(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='0' AND D( 0)='0' )then
          cVar1S12S116P060P062N050P068(0) <='1';
          else
          cVar1S12S116P060P062N050P068(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='0' AND D( 0)='0' )then
          cVar1S13S116P060P062N050P068(0) <='1';
          else
          cVar1S13S116P060P062N050P068(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='0' AND D( 0)='1' )then
          cVar1S14S116P060P062N050P068(0) <='1';
          else
          cVar1S14S116P060P062N050P068(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='0' AND D( 0)='1' )then
          cVar1S15S116P060P062N050P068(0) <='1';
          else
          cVar1S15S116P060P062N050P068(0) <='0';
          end if;
        if(D( 2)='0' AND E( 2)='1' AND E( 5)='0' AND D( 0)='1' )then
          cVar1S16S116P060P062N050P068(0) <='1';
          else
          cVar1S16S116P060P062N050P068(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='1' AND A(15)='0' AND B(13)='1' )then
          cVar1S17S116P060P014P008P032nsss(0) <='1';
          else
          cVar1S17S116P060P014P008P032nsss(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='1' AND A(15)='0' AND B(13)='0' )then
          cVar1S18S116P060P014P008N032(0) <='1';
          else
          cVar1S18S116P060P014P008N032(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='1' AND A(15)='0' AND B(13)='0' )then
          cVar1S19S116P060P014P008N032(0) <='1';
          else
          cVar1S19S116P060P014P008N032(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='1' )then
          cVar1S20S116P060N014P033P013(0) <='1';
          else
          cVar1S20S116P060N014P033P013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='1' )then
          cVar1S21S116P060N014P033P013(0) <='1';
          else
          cVar1S21S116P060N014P033P013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='1' )then
          cVar1S22S116P060N014P033P013(0) <='1';
          else
          cVar1S22S116P060N014P033P013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='0' )then
          cVar1S23S116P060N014P033N013(0) <='1';
          else
          cVar1S23S116P060N014P033N013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='0' )then
          cVar1S24S116P060N014P033N013(0) <='1';
          else
          cVar1S24S116P060N014P033N013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='1' AND A( 3)='0' )then
          cVar1S25S116P060N014P033N013(0) <='1';
          else
          cVar1S25S116P060N014P033N013(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='1' )then
          cVar1S26S116P060N014N033P066(0) <='1';
          else
          cVar1S26S116P060N014N033P066(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='1' )then
          cVar1S27S116P060N014N033P066(0) <='1';
          else
          cVar1S27S116P060N014N033P066(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='0' )then
          cVar1S28S116P060N014N033N066(0) <='1';
          else
          cVar1S28S116P060N014N033N066(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='0' )then
          cVar1S29S116P060N014N033N066(0) <='1';
          else
          cVar1S29S116P060N014N033N066(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='0' )then
          cVar1S30S116P060N014N033N066(0) <='1';
          else
          cVar1S30S116P060N014N033N066(0) <='0';
          end if;
        if(D( 2)='1' AND A(12)='0' AND B( 3)='0' AND E( 1)='0' )then
          cVar1S31S116P060N014N033N066(0) <='1';
          else
          cVar1S31S116P060N014N033N066(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='1' )then
          cVar1S0S117P049P005nsss(0) <='1';
          else
          cVar1S0S117P049P005nsss(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='1' AND B( 3)='0' )then
          cVar1S1S117P049N005P026P033nsss(0) <='1';
          else
          cVar1S1S117P049N005P026P033nsss(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='1' )then
          cVar1S2S117P049N005N026P024(0) <='1';
          else
          cVar1S2S117P049N005N026P024(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='1' )then
          cVar1S3S117P049N005N026P024(0) <='1';
          else
          cVar1S3S117P049N005N026P024(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='1' )then
          cVar1S4S117P049N005N026P024(0) <='1';
          else
          cVar1S4S117P049N005N026P024(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='0' )then
          cVar1S5S117P049N005N026N024(0) <='1';
          else
          cVar1S5S117P049N005N026N024(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='0' )then
          cVar1S6S117P049N005N026N024(0) <='1';
          else
          cVar1S6S117P049N005N026N024(0) <='0';
          end if;
        if(D(13)='1' AND A( 7)='0' AND B(16)='0' AND B(17)='0' )then
          cVar1S7S117P049N005N026N024(0) <='1';
          else
          cVar1S7S117P049N005N026N024(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='1' AND B(15)='1' )then
          cVar1S8S117N049P024P053P028(0) <='1';
          else
          cVar1S8S117N049P024P053P028(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='1' AND B(15)='1' )then
          cVar1S9S117N049P024P053P028(0) <='1';
          else
          cVar1S9S117N049P024P053P028(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='1' AND B(15)='0' )then
          cVar1S10S117N049P024P053N028(0) <='1';
          else
          cVar1S10S117N049P024P053N028(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='1' AND B(15)='0' )then
          cVar1S11S117N049P024P053N028(0) <='1';
          else
          cVar1S11S117N049P024P053N028(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='1' AND B(15)='0' )then
          cVar1S12S117N049P024P053N028(0) <='1';
          else
          cVar1S12S117N049P024P053N028(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='0' )then
          cVar1S13S117N049P024N053P051(0) <='1';
          else
          cVar1S13S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='0' )then
          cVar1S14S117N049P024N053P051(0) <='1';
          else
          cVar1S14S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='0' )then
          cVar1S15S117N049P024N053P051(0) <='1';
          else
          cVar1S15S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='0' )then
          cVar1S16S117N049P024N053P051(0) <='1';
          else
          cVar1S16S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='1' )then
          cVar1S17S117N049P024N053P051(0) <='1';
          else
          cVar1S17S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='0' AND D(12)='0' AND E(13)='1' )then
          cVar1S18S117N049P024N053P051(0) <='1';
          else
          cVar1S18S117N049P024N053P051(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='1' AND B(16)='0' AND A(18)='1' )then
          cVar1S19S117N049P024P026P002nsss(0) <='1';
          else
          cVar1S19S117N049P024P026P002nsss(0) <='0';
          end if;
        if(D(13)='0' AND B(17)='1' AND B(16)='0' AND A(18)='0' )then
          cVar1S20S117N049P024P026N002(0) <='1';
          else
          cVar1S20S117N049P024P026N002(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='1' AND B(17)='1' )then
          cVar1S0S118P049P006P024nsss(0) <='1';
          else
          cVar1S0S118P049P006P024nsss(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S118P049P006N024P026nsss(0) <='1';
          else
          cVar1S1S118P049P006N024P026nsss(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='1' AND A( 0)='0' )then
          cVar1S2S118P049N006P007P019(0) <='1';
          else
          cVar1S2S118P049N006P007P019(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='1' AND A( 0)='1' )then
          cVar1S3S118P049N006P007P019(0) <='1';
          else
          cVar1S3S118P049N006P007P019(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S4S118P049N006N007P009(0) <='1';
          else
          cVar1S4S118P049N006N007P009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S5S118P049N006N007P009(0) <='1';
          else
          cVar1S5S118P049N006N007P009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S6S118P049N006N007N009(0) <='1';
          else
          cVar1S6S118P049N006N007N009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S7S118P049N006N007N009(0) <='1';
          else
          cVar1S7S118P049N006N007N009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S8S118P049N006N007N009(0) <='1';
          else
          cVar1S8S118P049N006N007N009(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='1' )then
          cVar1S9S118N049P052P024P042(0) <='1';
          else
          cVar1S9S118N049P052P024P042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='1' )then
          cVar1S10S118N049P052P024P042(0) <='1';
          else
          cVar1S10S118N049P052P024P042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='1' )then
          cVar1S11S118N049P052P024P042(0) <='1';
          else
          cVar1S11S118N049P052P024P042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='0' )then
          cVar1S12S118N049P052P024N042(0) <='1';
          else
          cVar1S12S118N049P052P024N042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='0' )then
          cVar1S13S118N049P052P024N042(0) <='1';
          else
          cVar1S13S118N049P052P024N042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='0' AND E( 7)='0' )then
          cVar1S14S118N049P052P024N042(0) <='1';
          else
          cVar1S14S118N049P052P024N042(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='1' AND D( 0)='0' )then
          cVar1S15S118N049P052P024P068(0) <='1';
          else
          cVar1S15S118N049P052P024P068(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='1' AND D( 0)='0' )then
          cVar1S16S118N049P052P024P068(0) <='1';
          else
          cVar1S16S118N049P052P024P068(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='0' AND B(17)='1' AND D( 0)='1' )then
          cVar1S17S118N049P052P024P068(0) <='1';
          else
          cVar1S17S118N049P052P024P068(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='1' AND E( 1)='0' )then
          cVar1S18S118N049P052P065P066nsss(0) <='1';
          else
          cVar1S18S118N049P052P065P066nsss(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='0' AND E( 9)='1' )then
          cVar1S19S118N049P052N065P067(0) <='1';
          else
          cVar1S19S118N049P052N065P067(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='0' AND E( 9)='1' )then
          cVar1S20S118N049P052N065P067(0) <='1';
          else
          cVar1S20S118N049P052N065P067(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='0' AND E( 9)='0' )then
          cVar1S21S118N049P052N065N067(0) <='1';
          else
          cVar1S21S118N049P052N065N067(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='0' AND E( 9)='0' )then
          cVar1S22S118N049P052N065N067(0) <='1';
          else
          cVar1S22S118N049P052N065N067(0) <='0';
          end if;
        if(D(13)='0' AND D( 4)='1' AND D( 9)='0' AND E( 9)='0' )then
          cVar1S23S118N049P052N065N067(0) <='1';
          else
          cVar1S23S118N049P052N065N067(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='1' AND A( 6)='0' AND A(10)='0' )then
          cVar1S0S119P049P006P007P018nsss(0) <='1';
          else
          cVar1S0S119P049P006P007P018nsss(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='1' AND A( 6)='0' AND A(10)='1' )then
          cVar1S1S119P049P006P007P018(0) <='1';
          else
          cVar1S1S119P049P006P007P018(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar1S2S119P049N006P007P025nsss(0) <='1';
          else
          cVar1S2S119P049N006P007P025nsss(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='1' AND B( 7)='0' )then
          cVar1S3S119P049N006P007N025(0) <='1';
          else
          cVar1S3S119P049N006P007N025(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S4S119P049N006N007P009(0) <='1';
          else
          cVar1S4S119P049N006N007P009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S5S119P049N006N007P009(0) <='1';
          else
          cVar1S5S119P049N006N007P009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='1' )then
          cVar1S6S119P049N006N007P009(0) <='1';
          else
          cVar1S6S119P049N006N007P009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S7S119P049N006N007N009(0) <='1';
          else
          cVar1S7S119P049N006N007N009(0) <='0';
          end if;
        if(D(13)='1' AND A(16)='0' AND A( 6)='0' AND A( 5)='0' )then
          cVar1S8S119P049N006N007N009(0) <='1';
          else
          cVar1S8S119P049N006N007N009(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='1' )then
          cVar1S9S119N049P042P051nsss(0) <='1';
          else
          cVar1S9S119N049P042P051nsss(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='0' AND E( 5)='0' )then
          cVar1S10S119N049P042N051P050(0) <='1';
          else
          cVar1S10S119N049P042N051P050(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='0' AND E( 5)='0' )then
          cVar1S11S119N049P042N051P050(0) <='1';
          else
          cVar1S11S119N049P042N051P050(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='0' AND E( 5)='0' )then
          cVar1S12S119N049P042N051P050(0) <='1';
          else
          cVar1S12S119N049P042N051P050(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='1' )then
          cVar1S13S119N049N042P045P022nsss(0) <='1';
          else
          cVar1S13S119N049N042P045P022nsss(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S14S119N049N042P045N022(0) <='1';
          else
          cVar1S14S119N049N042P045N022(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S15S119N049N042P045N022(0) <='1';
          else
          cVar1S15S119N049N042P045N022(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S16S119N049N042P045N022(0) <='1';
          else
          cVar1S16S119N049N042P045N022(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S17S119N049N042N045P047(0) <='1';
          else
          cVar1S17S119N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S18S119N049N042N045P047(0) <='1';
          else
          cVar1S18S119N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S19S119N049N042N045P047(0) <='1';
          else
          cVar1S19S119N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S20S119N049N042N045P047(0) <='1';
          else
          cVar1S20S119N049N042N045P047(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='1' AND A(14)='0' AND A(16)='1' )then
          cVar1S0S120P049P024P010P006(0) <='1';
          else
          cVar1S0S120P049P024P010P006(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='1' AND A(14)='0' AND A(16)='1' )then
          cVar1S1S120P049P024P010P006(0) <='1';
          else
          cVar1S1S120P049P024P010P006(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='1' AND A(14)='0' AND A(16)='0' )then
          cVar1S2S120P049P024P010N006(0) <='1';
          else
          cVar1S2S120P049P024P010N006(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='1' )then
          cVar1S3S120P049N024P026P007nsss(0) <='1';
          else
          cVar1S3S120P049N024P026P007nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S4S120P049N024P026N007(0) <='1';
          else
          cVar1S4S120P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S5S120P049N024P026N007(0) <='1';
          else
          cVar1S5S120P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S6S120P049N024P026N007(0) <='1';
          else
          cVar1S6S120P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='1' )then
          cVar1S7S120P049N024N026P027nsss(0) <='1';
          else
          cVar1S7S120P049N024N026P027nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S8S120P049N024N026N027(0) <='1';
          else
          cVar1S8S120P049N024N026N027(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S9S120P049N024N026N027(0) <='1';
          else
          cVar1S9S120P049N024N026N027(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S10S120P049N024N026N027(0) <='1';
          else
          cVar1S10S120P049N024N026N027(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='1' )then
          cVar1S11S120N049P042P050P004(0) <='1';
          else
          cVar1S11S120N049P042P050P004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='1' )then
          cVar1S12S120N049P042P050P004(0) <='1';
          else
          cVar1S12S120N049P042P050P004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='1' )then
          cVar1S13S120N049P042P050P004(0) <='1';
          else
          cVar1S13S120N049P042P050P004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='0' )then
          cVar1S14S120N049P042P050N004(0) <='1';
          else
          cVar1S14S120N049P042P050N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='0' )then
          cVar1S15S120N049P042P050N004(0) <='1';
          else
          cVar1S15S120N049P042P050N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E( 5)='0' AND A(17)='0' )then
          cVar1S16S120N049P042P050N004(0) <='1';
          else
          cVar1S16S120N049P042P050N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='1' )then
          cVar1S17S120N049N042P045P022nsss(0) <='1';
          else
          cVar1S17S120N049N042P045P022nsss(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S18S120N049N042P045N022(0) <='1';
          else
          cVar1S18S120N049N042P045N022(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND B(18)='0' )then
          cVar1S19S120N049N042P045N022(0) <='1';
          else
          cVar1S19S120N049N042P045N022(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S20S120N049N042N045P047(0) <='1';
          else
          cVar1S20S120N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S21S120N049N042N045P047(0) <='1';
          else
          cVar1S21S120N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S22S120N049N042N045P047(0) <='1';
          else
          cVar1S22S120N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S23S120N049N042N045P047(0) <='1';
          else
          cVar1S23S120N049N042N045P047(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='1' AND A(14)='0' AND A(16)='1' )then
          cVar1S0S121P049P024P010P006nsss(0) <='1';
          else
          cVar1S0S121P049P024P010P006nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='1' AND A(14)='0' AND A(16)='0' )then
          cVar1S1S121P049P024P010N006(0) <='1';
          else
          cVar1S1S121P049P024P010N006(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='1' )then
          cVar1S2S121P049N024P026P007nsss(0) <='1';
          else
          cVar1S2S121P049N024P026P007nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S3S121P049N024P026N007(0) <='1';
          else
          cVar1S3S121P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S4S121P049N024P026N007(0) <='1';
          else
          cVar1S4S121P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='1' AND A( 6)='0' )then
          cVar1S5S121P049N024P026N007(0) <='1';
          else
          cVar1S5S121P049N024P026N007(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='1' )then
          cVar1S6S121P049N024N026P027nsss(0) <='1';
          else
          cVar1S6S121P049N024N026P027nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S7S121P049N024N026N027(0) <='1';
          else
          cVar1S7S121P049N024N026N027(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S8S121P049N024N026N027(0) <='1';
          else
          cVar1S8S121P049N024N026N027(0) <='0';
          end if;
        if(D(13)='1' AND B(17)='0' AND B(16)='0' AND B( 6)='0' )then
          cVar1S9S121P049N024N026N027(0) <='1';
          else
          cVar1S9S121P049N024N026N027(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='1' )then
          cVar1S10S121N049P042P051nsss(0) <='1';
          else
          cVar1S10S121N049P042P051nsss(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='1' AND E(13)='0' AND E( 5)='0' )then
          cVar1S11S121N049P042N051P050nsss(0) <='1';
          else
          cVar1S11S121N049P042N051P050nsss(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND A(17)='1' )then
          cVar1S12S121N049N042P045P004(0) <='1';
          else
          cVar1S12S121N049N042P045P004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S13S121N049N042P045N004(0) <='1';
          else
          cVar1S13S121N049N042P045N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S14S121N049N042P045N004(0) <='1';
          else
          cVar1S14S121N049N042P045N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S15S121N049N042P045N004(0) <='1';
          else
          cVar1S15S121N049N042P045N004(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S16S121N049N042N045P047(0) <='1';
          else
          cVar1S16S121N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S17S121N049N042N045P047(0) <='1';
          else
          cVar1S17S121N049N042N045P047(0) <='0';
          end if;
        if(D(13)='0' AND E( 7)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S18S121N049N042N045P047(0) <='1';
          else
          cVar1S18S121N049N042N045P047(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='1' AND A( 3)='1' )then
          cVar1S0S122P045P027P024P013nsss(0) <='1';
          else
          cVar1S0S122P045P027P024P013nsss(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='1' AND A( 3)='0' )then
          cVar1S1S122P045P027P024N013(0) <='1';
          else
          cVar1S1S122P045P027P024N013(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='1' AND A( 3)='0' )then
          cVar1S2S122P045P027P024N013(0) <='1';
          else
          cVar1S2S122P045P027P024N013(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='1' AND A( 3)='0' )then
          cVar1S3S122P045P027P024N013(0) <='1';
          else
          cVar1S3S122P045P027P024N013(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='0' AND B( 7)='1' )then
          cVar1S4S122P045P027N024P025(0) <='1';
          else
          cVar1S4S122P045P027N024P025(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='0' AND B( 7)='1' )then
          cVar1S5S122P045P027N024P025(0) <='1';
          else
          cVar1S5S122P045P027N024P025(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='0' AND B( 7)='0' )then
          cVar1S6S122P045P027N024N025(0) <='1';
          else
          cVar1S6S122P045P027N024N025(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='0' AND B( 7)='0' )then
          cVar1S7S122P045P027N024N025(0) <='1';
          else
          cVar1S7S122P045P027N024N025(0) <='0';
          end if;
        if(D(14)='1' AND B( 6)='0' AND B(17)='0' AND B( 7)='0' )then
          cVar1S8S122P045P027N024N025(0) <='1';
          else
          cVar1S8S122P045P027N024N025(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='1' AND B(16)='0' )then
          cVar1S9S122N045P049P024P026(0) <='1';
          else
          cVar1S9S122N045P049P024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='1' AND B(16)='0' )then
          cVar1S10S122N045P049P024P026(0) <='1';
          else
          cVar1S10S122N045P049P024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='1' AND B(16)='0' )then
          cVar1S11S122N045P049P024P026(0) <='1';
          else
          cVar1S11S122N045P049P024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S12S122N045P049N024P026(0) <='1';
          else
          cVar1S12S122N045P049N024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S13S122N045P049N024P026(0) <='1';
          else
          cVar1S13S122N045P049N024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S14S122N045P049N024P026(0) <='1';
          else
          cVar1S14S122N045P049N024P026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S15S122N045P049N024N026(0) <='1';
          else
          cVar1S15S122N045P049N024N026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S16S122N045P049N024N026(0) <='1';
          else
          cVar1S16S122N045P049N024N026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S17S122N045P049N024N026(0) <='1';
          else
          cVar1S17S122N045P049N024N026(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='1' )then
          cVar1S18S122N045N049P047P042(0) <='1';
          else
          cVar1S18S122N045N049P047P042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='1' )then
          cVar1S19S122N045N049P047P042(0) <='1';
          else
          cVar1S19S122N045N049P047P042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='1' )then
          cVar1S20S122N045N049P047P042(0) <='1';
          else
          cVar1S20S122N045N049P047P042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='0' )then
          cVar1S21S122N045N049P047N042(0) <='1';
          else
          cVar1S21S122N045N049P047N042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='0' )then
          cVar1S22S122N045N049P047N042(0) <='1';
          else
          cVar1S22S122N045N049P047N042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='0' )then
          cVar1S23S122N045N049P047N042(0) <='1';
          else
          cVar1S23S122N045N049P047N042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='0' AND E( 7)='0' )then
          cVar1S24S122N045N049P047N042(0) <='1';
          else
          cVar1S24S122N045N049P047N042(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='1' AND D( 1)='1' )then
          cVar1S25S122N045N049P047P064nsss(0) <='1';
          else
          cVar1S25S122N045N049P047P064nsss(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='1' AND D( 1)='0' )then
          cVar1S26S122N045N049P047N064(0) <='1';
          else
          cVar1S26S122N045N049P047N064(0) <='0';
          end if;
        if(D(14)='0' AND D(13)='0' AND E(14)='1' AND D( 1)='0' )then
          cVar1S27S122N045N049P047N064(0) <='1';
          else
          cVar1S27S122N045N049P047N064(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='1' )then
          cVar1S0S123P042P051nsss(0) <='1';
          else
          cVar1S0S123P042P051nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND E( 5)='0' AND B( 0)='1' )then
          cVar1S1S123P042N051P050P039nsss(0) <='1';
          else
          cVar1S1S123P042N051P050P039nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND E( 5)='0' AND B( 0)='0' )then
          cVar1S2S123P042N051P050N039(0) <='1';
          else
          cVar1S2S123P042N051P050N039(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND E( 5)='0' AND B( 0)='0' )then
          cVar1S3S123P042N051P050N039(0) <='1';
          else
          cVar1S3S123P042N051P050N039(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND E( 5)='0' AND B( 0)='0' )then
          cVar1S4S123P042N051P050N039(0) <='1';
          else
          cVar1S4S123P042N051P050N039(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='1' )then
          cVar1S5S123N042P049P024P004nsss(0) <='1';
          else
          cVar1S5S123N042P049P024P004nsss(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S6S123N042P049P024N004(0) <='1';
          else
          cVar1S6S123N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S7S123N042P049P024N004(0) <='1';
          else
          cVar1S7S123N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S8S123N042P049P024N004(0) <='1';
          else
          cVar1S8S123N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S9S123N042P049N024P026(0) <='1';
          else
          cVar1S9S123N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S10S123N042P049N024P026(0) <='1';
          else
          cVar1S10S123N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S11S123N042P049N024P026(0) <='1';
          else
          cVar1S11S123N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S12S123N042P049N024N026(0) <='1';
          else
          cVar1S12S123N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S13S123N042P049N024N026(0) <='1';
          else
          cVar1S13S123N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S14S123N042P049N024N026(0) <='1';
          else
          cVar1S14S123N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND A( 6)='1' )then
          cVar1S15S123N042N049P045P007(0) <='1';
          else
          cVar1S15S123N042N049P045P007(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND A( 6)='1' )then
          cVar1S16S123N042N049P045P007(0) <='1';
          else
          cVar1S16S123N042N049P045P007(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND A( 6)='0' )then
          cVar1S17S123N042N049P045N007(0) <='1';
          else
          cVar1S17S123N042N049P045N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND A( 6)='0' )then
          cVar1S18S123N042N049P045N007(0) <='1';
          else
          cVar1S18S123N042N049P045N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND A( 6)='0' )then
          cVar1S19S123N042N049P045N007(0) <='1';
          else
          cVar1S19S123N042N049P045N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S20S123N042N049N045P047(0) <='1';
          else
          cVar1S20S123N042N049N045P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND E(14)='0' )then
          cVar1S21S123N042N049N045P047(0) <='1';
          else
          cVar1S21S123N042N049N045P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND E(14)='1' )then
          cVar1S22S123N042N049N045P047(0) <='1';
          else
          cVar1S22S123N042N049N045P047(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND B( 9)='1' )then
          cVar1S0S124P042P050P021nsss(0) <='1';
          else
          cVar1S0S124P042P050P021nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND B( 9)='0' AND E(13)='1' )then
          cVar1S1S124P042P050N021P051nsss(0) <='1';
          else
          cVar1S1S124P042P050N021P051nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND B( 9)='0' AND E(13)='0' )then
          cVar1S2S124P042P050N021N051(0) <='1';
          else
          cVar1S2S124P042P050N021N051(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND B( 9)='0' AND E(13)='0' )then
          cVar1S3S124P042P050N021N051(0) <='1';
          else
          cVar1S3S124P042P050N021N051(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND B( 9)='0' AND E(13)='0' )then
          cVar1S4S124P042P050N021N051(0) <='1';
          else
          cVar1S4S124P042P050N021N051(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S5S124N042P045P027P024(0) <='1';
          else
          cVar1S5S124N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S6S124N042P045P027P024(0) <='1';
          else
          cVar1S6S124N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S7S124N042P045P027P024(0) <='1';
          else
          cVar1S7S124N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S8S124N042P045P027N024(0) <='1';
          else
          cVar1S8S124N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S9S124N042P045P027N024(0) <='1';
          else
          cVar1S9S124N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S10S124N042P045P027N024(0) <='1';
          else
          cVar1S10S124N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S11S124N042P045P027N024(0) <='1';
          else
          cVar1S11S124N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S12S124N042N045P049P024(0) <='1';
          else
          cVar1S12S124N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S13S124N042N045P049P024(0) <='1';
          else
          cVar1S13S124N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S14S124N042N045P049P024(0) <='1';
          else
          cVar1S14S124N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S15S124N042N045P049N024(0) <='1';
          else
          cVar1S15S124N042N045P049N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S16S124N042N045P049N024(0) <='1';
          else
          cVar1S16S124N042N045P049N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S17S124N042N045P049N024(0) <='1';
          else
          cVar1S17S124N042N045P049N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S18S124N042N045N049P047(0) <='1';
          else
          cVar1S18S124N042N045N049P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S19S124N042N045N049P047(0) <='1';
          else
          cVar1S19S124N042N045N049P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S20S124N042N045N049P047(0) <='1';
          else
          cVar1S20S124N042N045N049P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(14)='0' )then
          cVar1S21S124N042N045N049P047(0) <='1';
          else
          cVar1S21S124N042N045N049P047(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(14)='1' )then
          cVar1S22S124N042N045N049P047(0) <='1';
          else
          cVar1S22S124N042N045N049P047(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' )then
          cVar1S0S125P042P050nsss(0) <='1';
          else
          cVar1S0S125P042P050nsss(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S1S125N042P045P027P024(0) <='1';
          else
          cVar1S1S125N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S2S125N042P045P027P024(0) <='1';
          else
          cVar1S2S125N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S3S125N042P045P027P024(0) <='1';
          else
          cVar1S3S125N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S4S125N042P045P027N024psss(0) <='1';
          else
          cVar1S4S125N042P045P027N024psss(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S5S125N042N045P049P024(0) <='1';
          else
          cVar1S5S125N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S6S125N042N045P049P024(0) <='1';
          else
          cVar1S6S125N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='1' )then
          cVar1S7S125N042N045P049P024(0) <='1';
          else
          cVar1S7S125N042N045P049P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S8S125N042N045P049N024(0) <='1';
          else
          cVar1S8S125N042N045P049N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND B(17)='0' )then
          cVar1S9S125N042N045P049N024(0) <='1';
          else
          cVar1S9S125N042N045P049N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND B(13)='1' )then
          cVar1S10S125N042N045N049P032(0) <='1';
          else
          cVar1S10S125N042N045N049P032(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND B(13)='1' )then
          cVar1S11S125N042N045N049P032(0) <='1';
          else
          cVar1S11S125N042N045N049P032(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND B(13)='0' )then
          cVar1S12S125N042N045N049N032(0) <='1';
          else
          cVar1S12S125N042N045N049N032(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND B(13)='0' )then
          cVar1S13S125N042N045N049N032(0) <='1';
          else
          cVar1S13S125N042N045N049N032(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='1' )then
          cVar1S0S126P042P051nsss(0) <='1';
          else
          cVar1S0S126P042P051nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='1' AND A( 7)='1' )then
          cVar1S1S126P042N051P023P005nsss(0) <='1';
          else
          cVar1S1S126P042N051P023P005nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S2S126P042N051P023N005(0) <='1';
          else
          cVar1S2S126P042N051P023N005(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S3S126P042N051P023N005(0) <='1';
          else
          cVar1S3S126P042N051P023N005(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='1' AND A( 7)='0' )then
          cVar1S4S126P042N051P023N005(0) <='1';
          else
          cVar1S4S126P042N051P023N005(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='0' AND A(19)='1' )then
          cVar1S5S126P042N051N023P000nsss(0) <='1';
          else
          cVar1S5S126P042N051N023P000nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='0' AND A(19)='0' )then
          cVar1S6S126P042N051N023N000(0) <='1';
          else
          cVar1S6S126P042N051N023N000(0) <='0';
          end if;
        if(E( 7)='1' AND E(13)='0' AND B( 8)='0' AND A(19)='0' )then
          cVar1S7S126P042N051N023N000(0) <='1';
          else
          cVar1S7S126P042N051N023N000(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S8S126N042P045P027P024(0) <='1';
          else
          cVar1S8S126N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S9S126N042P045P027P024(0) <='1';
          else
          cVar1S9S126N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='1' )then
          cVar1S10S126N042P045P027P024(0) <='1';
          else
          cVar1S10S126N042P045P027P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S11S126N042P045P027N024(0) <='1';
          else
          cVar1S11S126N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S12S126N042P045P027N024(0) <='1';
          else
          cVar1S12S126N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S13S126N042P045P027N024(0) <='1';
          else
          cVar1S13S126N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='1' AND B( 6)='0' AND B(17)='0' )then
          cVar1S14S126N042P045P027N024(0) <='1';
          else
          cVar1S14S126N042P045P027N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND A( 6)='1' )then
          cVar1S15S126N042N045P049P007(0) <='1';
          else
          cVar1S15S126N042N045P049P007(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND A( 6)='0' )then
          cVar1S16S126N042N045P049N007(0) <='1';
          else
          cVar1S16S126N042N045P049N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND A( 6)='0' )then
          cVar1S17S126N042N045P049N007(0) <='1';
          else
          cVar1S17S126N042N045P049N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND A( 6)='0' )then
          cVar1S18S126N042N045P049N007(0) <='1';
          else
          cVar1S18S126N042N045P049N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='1' AND A( 6)='0' )then
          cVar1S19S126N042N045P049N007(0) <='1';
          else
          cVar1S19S126N042N045P049N007(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(11)='0' )then
          cVar1S20S126N042N045N049P059(0) <='1';
          else
          cVar1S20S126N042N045N049P059(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(11)='0' )then
          cVar1S21S126N042N045N049P059(0) <='1';
          else
          cVar1S21S126N042N045N049P059(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(11)='0' )then
          cVar1S22S126N042N045N049P059(0) <='1';
          else
          cVar1S22S126N042N045N049P059(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(11)='1' )then
          cVar1S23S126N042N045N049P059(0) <='1';
          else
          cVar1S23S126N042N045N049P059(0) <='0';
          end if;
        if(E( 7)='0' AND D(14)='0' AND D(13)='0' AND E(11)='1' )then
          cVar1S24S126N042N045N049P059(0) <='1';
          else
          cVar1S24S126N042N045N049P059(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='1' AND D( 7)='1' )then
          cVar1S0S127P042P050P004P040nsss(0) <='1';
          else
          cVar1S0S127P042P050P004P040nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='1' AND D( 7)='0' )then
          cVar1S1S127P042P050P004N040(0) <='1';
          else
          cVar1S1S127P042P050P004N040(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar1S2S127P042P050N004P005nsss(0) <='1';
          else
          cVar1S2S127P042P050N004P005nsss(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='0' AND A( 7)='0' )then
          cVar1S3S127P042P050N004N005(0) <='1';
          else
          cVar1S3S127P042P050N004N005(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='0' AND A( 7)='0' )then
          cVar1S4S127P042P050N004N005(0) <='1';
          else
          cVar1S4S127P042P050N004N005(0) <='0';
          end if;
        if(E( 7)='1' AND E( 5)='0' AND A(17)='0' AND A( 7)='0' )then
          cVar1S5S127P042P050N004N005(0) <='1';
          else
          cVar1S5S127P042P050N004N005(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='1' )then
          cVar1S6S127N042P049P024P004nsss(0) <='1';
          else
          cVar1S6S127N042P049P024P004nsss(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S7S127N042P049P024N004(0) <='1';
          else
          cVar1S7S127N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S8S127N042P049P024N004(0) <='1';
          else
          cVar1S8S127N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='1' AND A(17)='0' )then
          cVar1S9S127N042P049P024N004(0) <='1';
          else
          cVar1S9S127N042P049P024N004(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S10S127N042P049N024P026(0) <='1';
          else
          cVar1S10S127N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S11S127N042P049N024P026(0) <='1';
          else
          cVar1S11S127N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S12S127N042P049N024P026(0) <='1';
          else
          cVar1S12S127N042P049N024P026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S13S127N042P049N024N026(0) <='1';
          else
          cVar1S13S127N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S14S127N042P049N024N026(0) <='1';
          else
          cVar1S14S127N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S15S127N042P049N024N026(0) <='1';
          else
          cVar1S15S127N042P049N024N026(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='1' )then
          cVar1S16S127N042N049P045P024(0) <='1';
          else
          cVar1S16S127N042N049P045P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='1' )then
          cVar1S17S127N042N049P045P024(0) <='1';
          else
          cVar1S17S127N042N049P045P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='1' )then
          cVar1S18S127N042N049P045P024(0) <='1';
          else
          cVar1S18S127N042N049P045P024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='0' )then
          cVar1S19S127N042N049P045N024(0) <='1';
          else
          cVar1S19S127N042N049P045N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='0' )then
          cVar1S20S127N042N049P045N024(0) <='1';
          else
          cVar1S20S127N042N049P045N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='0' )then
          cVar1S21S127N042N049P045N024(0) <='1';
          else
          cVar1S21S127N042N049P045N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='1' AND B(17)='0' )then
          cVar1S22S127N042N049P045N024(0) <='1';
          else
          cVar1S22S127N042N049P045N024(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S23S127N042N049N045P020(0) <='1';
          else
          cVar1S23S127N042N049N045P020(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S24S127N042N049N045P020(0) <='1';
          else
          cVar1S24S127N042N049N045P020(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='1' )then
          cVar1S25S127N042N049N045P020(0) <='1';
          else
          cVar1S25S127N042N049N045P020(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S26S127N042N049N045N020(0) <='1';
          else
          cVar1S26S127N042N049N045N020(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S27S127N042N049N045N020(0) <='1';
          else
          cVar1S27S127N042N049N045N020(0) <='0';
          end if;
        if(E( 7)='0' AND D(13)='0' AND D(14)='0' AND B(19)='0' )then
          cVar1S28S127N042N049N045N020(0) <='1';
          else
          cVar1S28S127N042N049N045N020(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV2 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar1S3S0P055N030N031N028(0)='1' AND  B( 5)='1' )then
          cVar2S3S0P029nsss(0) <='1';
          else
          cVar2S3S0P029nsss(0) <='0';
          end if;
        if(cVar1S4S0P055N030N031N028(0)='1' AND  B( 5)='0' AND D(10)='1' )then
          cVar2S4S0N029P061nsss(0) <='1';
          else
          cVar2S4S0N029P061nsss(0) <='0';
          end if;
        if(cVar1S5S0P055N030N031N028(0)='1' AND  B( 5)='0' AND D(10)='0' AND D(13)='1' )then
          cVar2S5S0N029N061P049nsss(0) <='1';
          else
          cVar2S5S0N029N061P049nsss(0) <='0';
          end if;
        if(cVar1S7S0N055P059P061N032(0)='1' AND  D( 2)='1' )then
          cVar2S7S0P060nsss(0) <='1';
          else
          cVar2S7S0P060nsss(0) <='0';
          end if;
        if(cVar1S8S0N055P059P061N032(0)='1' AND  D( 2)='0' AND B( 3)='1' )then
          cVar2S8S0N060P033nsss(0) <='1';
          else
          cVar2S8S0N060P033nsss(0) <='0';
          end if;
        if(cVar1S9S0N055P059P061N032(0)='1' AND  D( 2)='0' AND B( 3)='0' AND B(12)='1' )then
          cVar2S9S0N060N033P034nsss(0) <='1';
          else
          cVar2S9S0N060N033P034nsss(0) <='0';
          end if;
        if(cVar1S11S0N055P059N061N058(0)='1' AND  E(10)='1' )then
          cVar2S11S0P063nsss(0) <='1';
          else
          cVar2S11S0P063nsss(0) <='0';
          end if;
        if(cVar1S12S0N055P059N061N058(0)='1' AND  E(10)='0' AND B(14)='1' )then
          cVar2S12S0N063P030nsss(0) <='1';
          else
          cVar2S12S0N063P030nsss(0) <='0';
          end if;
        if(cVar1S13S0N055P059N061N058(0)='1' AND  E(10)='0' AND B(14)='0' AND E( 9)='1' )then
          cVar2S13S0N063N030P067nsss(0) <='1';
          else
          cVar2S13S0N063N030P067nsss(0) <='0';
          end if;
        if(cVar1S15S0N055N059P052N029(0)='1' AND  B( 6)='1' )then
          cVar2S15S0P027nsss(0) <='1';
          else
          cVar2S15S0P027nsss(0) <='0';
          end if;
        if(cVar1S16S0N055N059P052N029(0)='1' AND  B( 6)='0' AND E(13)='1' )then
          cVar2S16S0N027P051nsss(0) <='1';
          else
          cVar2S16S0N027P051nsss(0) <='0';
          end if;
        if(cVar1S17S0N055N059P052N029(0)='1' AND  B( 6)='0' AND E(13)='0' AND B(15)='1' )then
          cVar2S17S0N027N051P028nsss(0) <='1';
          else
          cVar2S17S0N027N051P028nsss(0) <='0';
          end if;
        if(cVar1S18S0N055N059N052P047(0)='1' AND  D(13)='1' )then
          cVar2S18S0P049nsss(0) <='1';
          else
          cVar2S18S0P049nsss(0) <='0';
          end if;
        if(cVar1S19S0N055N059N052P047(0)='1' AND  D(13)='0' AND B(17)='1' )then
          cVar2S19S0N049P024nsss(0) <='1';
          else
          cVar2S19S0N049P024nsss(0) <='0';
          end if;
        if(cVar1S20S0N055N059N052P047(0)='1' AND  D(13)='0' AND B(17)='0' AND B( 7)='1' )then
          cVar2S20S0N049N024P025nsss(0) <='1';
          else
          cVar2S20S0N049N024P025nsss(0) <='0';
          end if;
        if(cVar1S21S0N055N059N052N047(0)='1' AND  D( 9)='1' AND E(10)='1' )then
          cVar2S21S0P065P063nsss(0) <='1';
          else
          cVar2S21S0P065P063nsss(0) <='0';
          end if;
        if(cVar1S22S0N055N059N052N047(0)='1' AND  D( 9)='0' AND E(15)='1' )then
          cVar2S22S0N065P043nsss(0) <='1';
          else
          cVar2S22S0N065P043nsss(0) <='0';
          end if;
        if(cVar1S23S0N055N059N052N047(0)='1' AND  D( 9)='0' AND E(15)='0' AND E( 9)='1' )then
          cVar2S23S0N065N043P067nsss(0) <='1';
          else
          cVar2S23S0N065N043P067nsss(0) <='0';
          end if;
        if(cVar1S1S1P058P033N060P018(0)='1' AND  D( 3)='1' )then
          cVar2S1S1P056nsss(0) <='1';
          else
          cVar2S1S1P056nsss(0) <='0';
          end if;
        if(cVar1S2S1P058P033N060P018(0)='1' AND  D( 3)='0' AND E(11)='1' )then
          cVar2S2S1N056P059nsss(0) <='1';
          else
          cVar2S2S1N056P059nsss(0) <='0';
          end if;
        if(cVar1S5S1P058N033N031N032(0)='1' AND  B(14)='1' )then
          cVar2S5S1P030nsss(0) <='1';
          else
          cVar2S5S1P030nsss(0) <='0';
          end if;
        if(cVar1S6S1P058N033N031N032(0)='1' AND  B(14)='0' AND B( 2)='1' )then
          cVar2S6S1N030P035nsss(0) <='1';
          else
          cVar2S6S1N030P035nsss(0) <='0';
          end if;
        if(cVar1S7S1P058N033N031N032(0)='1' AND  B(14)='0' AND B( 2)='0' AND D(12)='1' )then
          cVar2S7S1N030N035P053nsss(0) <='1';
          else
          cVar2S7S1N030N035P053nsss(0) <='0';
          end if;
        if(cVar1S9S1N058P051P053N028(0)='1' AND  B(16)='1' )then
          cVar2S9S1P026nsss(0) <='1';
          else
          cVar2S9S1P026nsss(0) <='0';
          end if;
        if(cVar1S10S1N058P051P053N028(0)='1' AND  B(16)='0' AND B( 5)='1' )then
          cVar2S10S1N026P029nsss(0) <='1';
          else
          cVar2S10S1N026P029nsss(0) <='0';
          end if;
        if(cVar1S11S1N058P051P053N028(0)='1' AND  B(16)='0' AND B( 5)='0' AND B( 6)='1' )then
          cVar2S11S1N026N029P027nsss(0) <='1';
          else
          cVar2S11S1N026N029P027nsss(0) <='0';
          end if;
        if(cVar1S13S1N058P051N053N026(0)='1' AND  B( 6)='1' )then
          cVar2S13S1P027nsss(0) <='1';
          else
          cVar2S13S1P027nsss(0) <='0';
          end if;
        if(cVar1S14S1N058P051N053N026(0)='1' AND  B( 6)='0' AND E( 4)='1' )then
          cVar2S14S1N027P054nsss(0) <='1';
          else
          cVar2S14S1N027P054nsss(0) <='0';
          end if;
        if(cVar1S15S1N058P051N053N026(0)='1' AND  B( 6)='0' AND E( 4)='0' AND B(13)='1' )then
          cVar2S15S1N027N054P032nsss(0) <='1';
          else
          cVar2S15S1N027N054P032nsss(0) <='0';
          end if;
        if(cVar1S17S1N058N051P046N025(0)='1' AND  B( 6)='1' )then
          cVar2S17S1P027nsss(0) <='1';
          else
          cVar2S17S1P027nsss(0) <='0';
          end if;
        if(cVar1S18S1N058N051P046N025(0)='1' AND  B( 6)='0' AND B(17)='1' )then
          cVar2S18S1N027P024nsss(0) <='1';
          else
          cVar2S18S1N027P024nsss(0) <='0';
          end if;
        if(cVar1S19S1N058N051P046N025(0)='1' AND  B( 6)='0' AND B(17)='0' AND B(16)='1' )then
          cVar2S19S1N027N024P026nsss(0) <='1';
          else
          cVar2S19S1N027N024P026nsss(0) <='0';
          end if;
        if(cVar1S20S1N058N051N046P064(0)='1' AND  B( 2)='1' AND E( 2)='1' )then
          cVar2S20S1P035P062nsss(0) <='1';
          else
          cVar2S20S1P035P062nsss(0) <='0';
          end if;
        if(cVar1S21S1N058N051N046P064(0)='1' AND  B( 2)='0' AND B( 1)='1' )then
          cVar2S21S1N035P037nsss(0) <='1';
          else
          cVar2S21S1N035P037nsss(0) <='0';
          end if;
        if(cVar1S22S1N058N051N046P064(0)='1' AND  B( 2)='0' AND B( 1)='0' AND B(12)='1' )then
          cVar2S22S1N035N037P034nsss(0) <='1';
          else
          cVar2S22S1N035N037P034nsss(0) <='0';
          end if;
        if(cVar1S23S1N058N051N046N064(0)='1' AND  E( 4)='1' AND D( 3)='1' )then
          cVar2S23S1P054P056nsss(0) <='1';
          else
          cVar2S23S1P054P056nsss(0) <='0';
          end if;
        if(cVar1S24S1N058N051N046N064(0)='1' AND  E( 4)='1' AND D( 3)='0' AND B( 5)='1' )then
          cVar2S24S1P054N056P029nsss(0) <='1';
          else
          cVar2S24S1P054N056P029nsss(0) <='0';
          end if;
        if(cVar1S25S1N058N051N046N064(0)='1' AND  E( 4)='0' AND E( 7)='1' )then
          cVar2S25S1N054P042nsss(0) <='1';
          else
          cVar2S25S1N054P042nsss(0) <='0';
          end if;
        if(cVar1S26S1N058N051N046N064(0)='1' AND  E( 4)='0' AND E( 7)='0' AND B( 0)='1' )then
          cVar2S26S1N054N042P039nsss(0) <='1';
          else
          cVar2S26S1N054N042P039nsss(0) <='0';
          end if;
        if(cVar1S1S2P068P019P015N066(0)='1' AND  A( 3)='0' AND E( 9)='0' )then
          cVar2S1S2P013P067nsss(0) <='1';
          else
          cVar2S1S2P013P067nsss(0) <='0';
          end if;
        if(cVar1S2S2P068P019P015P064(0)='1' AND  E( 1)='1' )then
          cVar2S2S2P066nsss(0) <='1';
          else
          cVar2S2S2P066nsss(0) <='0';
          end if;
        if(cVar1S3S2P068P019P015P064(0)='1' AND  E( 1)='0' AND A(11)='0' )then
          cVar2S3S2N066P016nsss(0) <='1';
          else
          cVar2S3S2N066P016nsss(0) <='0';
          end if;
        if(cVar1S4S2P068P019P015P064(0)='1' AND  E( 2)='1' )then
          cVar2S4S2P062nsss(0) <='1';
          else
          cVar2S4S2P062nsss(0) <='0';
          end if;
        if(cVar1S6S2P068N019P011N018(0)='1' AND  A( 1)='1' )then
          cVar2S6S2P017nsss(0) <='1';
          else
          cVar2S6S2P017nsss(0) <='0';
          end if;
        if(cVar1S7S2P068N019P011N018(0)='1' AND  A( 1)='0' AND E( 9)='0' AND D( 1)='0' )then
          cVar2S7S2N017P067P064nsss(0) <='1';
          else
          cVar2S7S2N017P067P064nsss(0) <='0';
          end if;
        if(cVar1S8S2P068N019P011P067(0)='1' AND  D( 9)='0' AND D( 4)='1' )then
          cVar2S8S2P065P052nsss(0) <='1';
          else
          cVar2S8S2P065P052nsss(0) <='0';
          end if;
        if(cVar1S9S2P068N019P011P067(0)='1' AND  D( 9)='0' AND D( 4)='0' AND A( 1)='1' )then
          cVar2S9S2P065N052P017nsss(0) <='1';
          else
          cVar2S9S2P065N052P017nsss(0) <='0';
          end if;
        if(cVar1S10S2P068N019P011P067(0)='1' AND  B( 1)='0' AND A(10)='1' )then
          cVar2S10S2P037P018nsss(0) <='1';
          else
          cVar2S10S2P037P018nsss(0) <='0';
          end if;
        if(cVar1S13S2N068P040N038N023(0)='1' AND  B( 9)='1' )then
          cVar2S13S2P021nsss(0) <='1';
          else
          cVar2S13S2P021nsss(0) <='0';
          end if;
        if(cVar1S14S2N068P040N038N023(0)='1' AND  B( 9)='0' AND A(17)='1' )then
          cVar2S14S2N021P004nsss(0) <='1';
          else
          cVar2S14S2N021P004nsss(0) <='0';
          end if;
        if(cVar1S15S2N068P040N038N023(0)='1' AND  B( 9)='0' AND A(17)='0' AND E( 6)='1' )then
          cVar2S15S2N021N004P046nsss(0) <='1';
          else
          cVar2S15S2N021N004P046nsss(0) <='0';
          end if;
        if(cVar1S17S2N068N040P050N027(0)='1' AND  D( 4)='1' )then
          cVar2S17S2P052nsss(0) <='1';
          else
          cVar2S17S2P052nsss(0) <='0';
          end if;
        if(cVar1S18S2N068N040P050N027(0)='1' AND  D( 4)='0' AND B(16)='1' )then
          cVar2S18S2N052P026nsss(0) <='1';
          else
          cVar2S18S2N052P026nsss(0) <='0';
          end if;
        if(cVar1S19S2N068N040P050N027(0)='1' AND  D( 4)='0' AND B(16)='0' AND E(13)='1' )then
          cVar2S19S2N052N026P051nsss(0) <='1';
          else
          cVar2S19S2N052N026P051nsss(0) <='0';
          end if;
        if(cVar1S20S2N068N040N050P046(0)='1' AND  B( 7)='1' )then
          cVar2S20S2P025nsss(0) <='1';
          else
          cVar2S20S2P025nsss(0) <='0';
          end if;
        if(cVar1S21S2N068N040N050P046(0)='1' AND  B( 7)='0' AND B(11)='0' )then
          cVar2S21S2N025P036nsss(0) <='1';
          else
          cVar2S21S2N025P036nsss(0) <='0';
          end if;
        if(cVar1S22S2N068N040N050N046(0)='1' AND  D( 2)='1' AND B( 3)='1' )then
          cVar2S22S2P060P033nsss(0) <='1';
          else
          cVar2S22S2P060P033nsss(0) <='0';
          end if;
        if(cVar1S23S2N068N040N050N046(0)='1' AND  D( 2)='1' AND B( 3)='0' AND E( 9)='0' )then
          cVar2S23S2P060N033P067nsss(0) <='1';
          else
          cVar2S23S2P060N033P067nsss(0) <='0';
          end if;
        if(cVar1S24S2N068N040N050N046(0)='1' AND  D( 2)='0' )then
          cVar2S24S2N060psss(0) <='1';
          else
          cVar2S24S2N060psss(0) <='0';
          end if;
        if(cVar1S0S3P068P019P015P017(0)='1' AND  A( 3)='0' )then
          cVar2S0S3P013nsss(0) <='1';
          else
          cVar2S0S3P013nsss(0) <='0';
          end if;
        if(cVar1S1S3P068P019P015P017(0)='1' AND  A( 3)='1' AND B( 1)='1' )then
          cVar2S1S3P013P037nsss(0) <='1';
          else
          cVar2S1S3P013P037nsss(0) <='0';
          end if;
        if(cVar1S2S3P068P019P015P017(0)='1' AND  A( 3)='1' AND B( 1)='0' AND A(11)='0' )then
          cVar2S2S3P013N037P016nsss(0) <='1';
          else
          cVar2S2S3P013N037P016nsss(0) <='0';
          end if;
        if(cVar1S3S3P068P019P015P017(0)='1' AND  E( 1)='1' AND A(10)='0' )then
          cVar2S3S3P066P018nsss(0) <='1';
          else
          cVar2S3S3P066P018nsss(0) <='0';
          end if;
        if(cVar1S4S3P068P019P015P017(0)='1' AND  E( 1)='1' AND A(10)='1' AND A(12)='0' )then
          cVar2S4S3P066P018P014nsss(0) <='1';
          else
          cVar2S4S3P066P018P014nsss(0) <='0';
          end if;
        if(cVar1S5S3P068P019P015P017(0)='1' AND  E( 1)='0' AND A(11)='0' )then
          cVar2S5S3N066P016nsss(0) <='1';
          else
          cVar2S5S3N066P016nsss(0) <='0';
          end if;
        if(cVar1S6S3P068P019P015P064(0)='1' AND  E( 1)='1' AND D( 3)='0' )then
          cVar2S6S3P066P056nsss(0) <='1';
          else
          cVar2S6S3P066P056nsss(0) <='0';
          end if;
        if(cVar1S7S3P068P019P015P064(0)='1' AND  E( 1)='0' AND A(12)='0' AND A(10)='0' )then
          cVar2S7S3N066P014P018nsss(0) <='1';
          else
          cVar2S7S3N066P014P018nsss(0) <='0';
          end if;
        if(cVar1S8S3P068P019P015P064(0)='1' AND  A( 5)='0' AND A( 1)='0' )then
          cVar2S8S3P009P017nsss(0) <='1';
          else
          cVar2S8S3P009P017nsss(0) <='0';
          end if;
        if(cVar1S9S3P068N019P018P001(0)='1' AND  A( 2)='0' AND E( 1)='1' )then
          cVar2S9S3P015P066nsss(0) <='1';
          else
          cVar2S9S3P015P066nsss(0) <='0';
          end if;
        if(cVar1S10S3P068N019P018P001(0)='1' AND  A( 2)='0' AND E( 1)='0' AND A(12)='0' )then
          cVar2S10S3P015N066P014nsss(0) <='1';
          else
          cVar2S10S3P015N066P014nsss(0) <='0';
          end if;
        if(cVar1S11S3P068N019P018P001(0)='1' AND  A( 2)='1' AND A(11)='0' )then
          cVar2S11S3P015P016nsss(0) <='1';
          else
          cVar2S11S3P015P016nsss(0) <='0';
          end if;
        if(cVar1S12S3P068N019P018P001(0)='1' AND  A( 2)='1' AND A(11)='1' AND A( 3)='0' )then
          cVar2S12S3P015P016P013nsss(0) <='1';
          else
          cVar2S12S3P015P016P013nsss(0) <='0';
          end if;
        if(cVar1S13S3P068N019N018P010(0)='1' AND  A( 1)='1' AND B( 1)='1' AND A( 3)='0' )then
          cVar2S13S3P017P037P013nsss(0) <='1';
          else
          cVar2S13S3P017P037P013nsss(0) <='0';
          end if;
        if(cVar1S14S3P068N019N018P010(0)='1' AND  A( 1)='1' AND B( 1)='0' AND B( 2)='1' )then
          cVar2S14S3P017N037P035nsss(0) <='1';
          else
          cVar2S14S3P017N037P035nsss(0) <='0';
          end if;
        if(cVar1S15S3P068N019N018P010(0)='1' AND  A( 1)='0' AND A(11)='1' AND A(12)='0' )then
          cVar2S15S3N017P016P014nsss(0) <='1';
          else
          cVar2S15S3N017P016P014nsss(0) <='0';
          end if;
        if(cVar1S16S3P068N019N018P010(0)='1' AND  A( 1)='0' AND A(11)='0' AND B( 1)='0' )then
          cVar2S16S3N017N016P037nsss(0) <='1';
          else
          cVar2S16S3N017N016P037nsss(0) <='0';
          end if;
        if(cVar1S17S3P068N019N018P010(0)='1' AND  B(11)='0' AND E(12)='1' )then
          cVar2S17S3P036P055nsss(0) <='1';
          else
          cVar2S17S3P036P055nsss(0) <='0';
          end if;
        if(cVar1S18S3P068N019N018P010(0)='1' AND  B(11)='0' AND E(12)='0' AND A( 1)='1' )then
          cVar2S18S3P036N055P017nsss(0) <='1';
          else
          cVar2S18S3P036N055P017nsss(0) <='0';
          end if;
        if(cVar1S21S3N068P040N021N020(0)='1' AND  B( 8)='1' )then
          cVar2S21S3P023nsss(0) <='1';
          else
          cVar2S21S3P023nsss(0) <='0';
          end if;
        if(cVar1S22S3N068P040N021N020(0)='1' AND  B( 8)='0' AND B(18)='1' )then
          cVar2S22S3N023P022nsss(0) <='1';
          else
          cVar2S22S3N023P022nsss(0) <='0';
          end if;
        if(cVar1S23S3N068P040N021N020(0)='1' AND  B( 8)='0' AND B(18)='0' AND E( 6)='1' )then
          cVar2S23S3N023N022P046nsss(0) <='1';
          else
          cVar2S23S3N023N022P046nsss(0) <='0';
          end if;
        if(cVar1S26S3N068N040N050N046(0)='1' AND  D( 2)='1' )then
          cVar2S26S3P060nsss(0) <='1';
          else
          cVar2S26S3P060nsss(0) <='0';
          end if;
        if(cVar1S27S3N068N040N050N046(0)='1' AND  D( 2)='0' AND E(13)='1' AND D(12)='1' )then
          cVar2S27S3N060P051P053nsss(0) <='1';
          else
          cVar2S27S3N060P051P053nsss(0) <='0';
          end if;
        if(cVar1S28S3N068N040N050N046(0)='1' AND  D( 2)='0' AND E(13)='0' AND D(11)='1' )then
          cVar2S28S3N060N051P057nsss(0) <='1';
          else
          cVar2S28S3N060N051P057nsss(0) <='0';
          end if;
        if(cVar1S2S4P040N038P067N023(0)='1' AND  D( 0)='0' )then
          cVar2S2S4P068nsss(0) <='1';
          else
          cVar2S2S4P068nsss(0) <='0';
          end if;
        if(cVar1S5S4N040P044N023N022(0)='1' AND  B( 7)='1' )then
          cVar2S5S4P025nsss(0) <='1';
          else
          cVar2S5S4P025nsss(0) <='0';
          end if;
        if(cVar1S6S4N040P044N023N022(0)='1' AND  B( 7)='0' AND B(17)='1' )then
          cVar2S6S4N025P024nsss(0) <='1';
          else
          cVar2S6S4N025P024nsss(0) <='0';
          end if;
        if(cVar1S7S4N040P044N023N022(0)='1' AND  B( 7)='0' AND B(17)='0' AND E( 5)='1' )then
          cVar2S7S4N025N024P050nsss(0) <='1';
          else
          cVar2S7S4N025N024P050nsss(0) <='0';
          end if;
        if(cVar1S9S4N040N044P047N024(0)='1' AND  B(16)='1' )then
          cVar2S9S4P026nsss(0) <='1';
          else
          cVar2S9S4P026nsss(0) <='0';
          end if;
        if(cVar1S10S4N040N044P047N024(0)='1' AND  B(16)='0' AND B( 7)='1' )then
          cVar2S10S4N026P025nsss(0) <='1';
          else
          cVar2S10S4N026P025nsss(0) <='0';
          end if;
        if(cVar1S11S4N040N044P047N024(0)='1' AND  B(16)='0' AND B( 7)='0' AND B( 6)='1' )then
          cVar2S11S4N026N025P027nsss(0) <='1';
          else
          cVar2S11S4N026N025P027nsss(0) <='0';
          end if;
        if(cVar1S12S4N040N044N047P061(0)='1' AND  E(11)='1' AND E( 3)='0' )then
          cVar2S12S4P059P058nsss(0) <='1';
          else
          cVar2S12S4P059P058nsss(0) <='0';
          end if;
        if(cVar1S13S4N040N044N047P061(0)='1' AND  E(11)='1' AND E( 3)='1' AND A(13)='0' )then
          cVar2S13S4P059P058P012nsss(0) <='1';
          else
          cVar2S13S4P059P058P012nsss(0) <='0';
          end if;
        if(cVar1S14S4N040N044N047P061(0)='1' AND  E(11)='0' AND E(10)='1' AND D( 9)='0' )then
          cVar2S14S4N059P063P065nsss(0) <='1';
          else
          cVar2S14S4N059P063P065nsss(0) <='0';
          end if;
        if(cVar1S15S4N040N044N047P061(0)='1' AND  E(11)='0' AND E(10)='0' AND E( 4)='1' )then
          cVar2S15S4N059N063P054nsss(0) <='1';
          else
          cVar2S15S4N059N063P054nsss(0) <='0';
          end if;
        if(cVar1S16S4N040N044N047N061(0)='1' AND  D( 3)='1' AND B( 4)='1' )then
          cVar2S16S4P056P031nsss(0) <='1';
          else
          cVar2S16S4P056P031nsss(0) <='0';
          end if;
        if(cVar1S17S4N040N044N047N061(0)='1' AND  D( 3)='1' AND B( 4)='0' AND B( 5)='1' )then
          cVar2S17S4P056N031P029nsss(0) <='1';
          else
          cVar2S17S4P056N031P029nsss(0) <='0';
          end if;
        if(cVar1S18S4N040N044N047N061(0)='1' AND  D( 3)='0' )then
          cVar2S18S4N056psss(0) <='1';
          else
          cVar2S18S4N056psss(0) <='0';
          end if;
        if(cVar1S3S5P044N023N022N025(0)='1' AND  B(17)='1' )then
          cVar2S3S5P024nsss(0) <='1';
          else
          cVar2S3S5P024nsss(0) <='0';
          end if;
        if(cVar1S4S5P044N023N022N025(0)='1' AND  B(17)='0' AND E( 4)='1' )then
          cVar2S4S5N024P054nsss(0) <='1';
          else
          cVar2S4S5N024P054nsss(0) <='0';
          end if;
        if(cVar1S7S5N044P040N021N020(0)='1' AND  B( 8)='1' )then
          cVar2S7S5P023nsss(0) <='1';
          else
          cVar2S7S5P023nsss(0) <='0';
          end if;
        if(cVar1S8S5N044P040N021N020(0)='1' AND  B( 8)='0' AND A(19)='1' )then
          cVar2S8S5N023P000nsss(0) <='1';
          else
          cVar2S8S5N023P000nsss(0) <='0';
          end if;
        if(cVar1S9S5N044P040N021N020(0)='1' AND  B( 8)='0' AND A(19)='0' AND A( 2)='0' )then
          cVar2S9S5N023N000P015nsss(0) <='1';
          else
          cVar2S9S5N023N000P015nsss(0) <='0';
          end if;
        if(cVar1S11S5N044N040P047N006(0)='1' AND  E( 1)='0' )then
          cVar2S11S5P066nsss(0) <='1';
          else
          cVar2S11S5P066nsss(0) <='0';
          end if;
        if(cVar1S12S5N044N040P047N006(0)='1' AND  E( 1)='1' AND D( 1)='0' AND E( 9)='1' )then
          cVar2S12S5P066P064P067nsss(0) <='1';
          else
          cVar2S12S5P066P064P067nsss(0) <='0';
          end if;
        if(cVar1S13S5N044N040N047P056(0)='1' AND  B( 4)='1' AND A( 3)='1' )then
          cVar2S13S5P031P013nsss(0) <='1';
          else
          cVar2S13S5P031P013nsss(0) <='0';
          end if;
        if(cVar1S14S5N044N040N047P056(0)='1' AND  B( 4)='1' AND A( 3)='0' AND E(12)='0' )then
          cVar2S14S5P031N013P055nsss(0) <='1';
          else
          cVar2S14S5P031N013P055nsss(0) <='0';
          end if;
        if(cVar1S15S5N044N040N047P056(0)='1' AND  B( 4)='0' AND B(14)='1' )then
          cVar2S15S5N031P030nsss(0) <='1';
          else
          cVar2S15S5N031P030nsss(0) <='0';
          end if;
        if(cVar1S16S5N044N040N047P056(0)='1' AND  B( 4)='0' AND B(14)='0' AND B( 5)='1' )then
          cVar2S16S5N031N030P029nsss(0) <='1';
          else
          cVar2S16S5N031N030P029nsss(0) <='0';
          end if;
        if(cVar1S17S5N044N040N047N056(0)='1' AND  D(10)='1' AND B(13)='1' AND E( 3)='0' )then
          cVar2S17S5P061P032P058nsss(0) <='1';
          else
          cVar2S17S5P061P032P058nsss(0) <='0';
          end if;
        if(cVar1S18S5N044N040N047N056(0)='1' AND  D(10)='1' AND B(13)='0' AND E(11)='1' )then
          cVar2S18S5P061N032P059nsss(0) <='1';
          else
          cVar2S18S5P061N032P059nsss(0) <='0';
          end if;
        if(cVar1S19S5N044N040N047N056(0)='1' AND  D(10)='0' AND D(15)='1' )then
          cVar2S19S5N061P041nsss(0) <='1';
          else
          cVar2S19S5N061P041nsss(0) <='0';
          end if;
        if(cVar1S20S5N044N040N047N056(0)='1' AND  D(10)='0' AND D(15)='0' AND D(14)='1' )then
          cVar2S20S5N061N041P045nsss(0) <='1';
          else
          cVar2S20S5N061N041P045nsss(0) <='0';
          end if;
        if(cVar1S3S6P044N023N004N006(0)='1' AND  A( 6)='1' AND B( 7)='1' )then
          cVar2S3S6P007P025nsss(0) <='1';
          else
          cVar2S3S6P007P025nsss(0) <='0';
          end if;
        if(cVar1S4S6P044N023N004N006(0)='1' AND  A( 6)='0' AND A(12)='0' )then
          cVar2S4S6N007P014nsss(0) <='1';
          else
          cVar2S4S6N007P014nsss(0) <='0';
          end if;
        if(cVar1S6S6N044P015P050N027(0)='1' AND  B(16)='1' )then
          cVar2S6S6P026nsss(0) <='1';
          else
          cVar2S6S6P026nsss(0) <='0';
          end if;
        if(cVar1S7S6N044P015P050N027(0)='1' AND  B(16)='0' AND B( 5)='1' AND D( 5)='0' )then
          cVar2S7S6N026P029P048nsss(0) <='1';
          else
          cVar2S7S6N026P029P048nsss(0) <='0';
          end if;
        if(cVar1S8S6N044P015P050N027(0)='1' AND  B(16)='0' AND B( 5)='0' AND A(14)='1' )then
          cVar2S8S6N026N029P010nsss(0) <='1';
          else
          cVar2S8S6N026N029P010nsss(0) <='0';
          end if;
        if(cVar1S9S6N044P015N050P056(0)='1' AND  B( 4)='1' AND A( 5)='0' )then
          cVar2S9S6P031P009nsss(0) <='1';
          else
          cVar2S9S6P031P009nsss(0) <='0';
          end if;
        if(cVar1S10S6N044P015N050P056(0)='1' AND  B( 4)='0' AND A( 3)='0' )then
          cVar2S10S6N031P013nsss(0) <='1';
          else
          cVar2S10S6N031P013nsss(0) <='0';
          end if;
        if(cVar1S11S6N044P015N050P056(0)='1' AND  B( 4)='0' AND A( 3)='1' AND B( 5)='1' )then
          cVar2S11S6N031P013P029nsss(0) <='1';
          else
          cVar2S11S6N031P013P029nsss(0) <='0';
          end if;
        if(cVar1S12S6N044P015N050N056(0)='1' AND  D( 7)='1' )then
          cVar2S12S6P040nsss(0) <='1';
          else
          cVar2S12S6P040nsss(0) <='0';
          end if;
        if(cVar1S13S6N044P015N050N056(0)='1' AND  D( 7)='0' AND E( 7)='0' )then
          cVar2S13S6N040P042nsss(0) <='1';
          else
          cVar2S13S6N040P042nsss(0) <='0';
          end if;
        if(cVar1S14S6N044P015P062P035(0)='1' AND  A(13)='0' AND B( 1)='0' )then
          cVar2S14S6P012P037nsss(0) <='1';
          else
          cVar2S14S6P012P037nsss(0) <='0';
          end if;
        if(cVar1S15S6N044P015P062P035(0)='1' AND  A(13)='0' AND B( 1)='1' AND A(12)='0' )then
          cVar2S15S6P012P037P014nsss(0) <='1';
          else
          cVar2S15S6P012P037P014nsss(0) <='0';
          end if;
        if(cVar1S16S6N044P015P062P035(0)='1' AND  A(13)='1' AND E(10)='0' AND A( 1)='1' )then
          cVar2S16S6P012P063P017nsss(0) <='1';
          else
          cVar2S16S6P012P063P017nsss(0) <='0';
          end if;
        if(cVar1S17S6N044P015P062N035(0)='1' AND  E( 3)='1' AND A(13)='0' )then
          cVar2S17S6P058P012nsss(0) <='1';
          else
          cVar2S17S6P058P012nsss(0) <='0';
          end if;
        if(cVar1S18S6N044P015P062N035(0)='1' AND  E( 3)='0' AND B( 1)='0' AND B( 3)='1' )then
          cVar2S18S6N058P037P033nsss(0) <='1';
          else
          cVar2S18S6N058P037P033nsss(0) <='0';
          end if;
        if(cVar1S19S6N044P015N062P058(0)='1' AND  B( 3)='1' AND A( 1)='0' )then
          cVar2S19S6P033P017nsss(0) <='1';
          else
          cVar2S19S6P033P017nsss(0) <='0';
          end if;
        if(cVar1S20S6N044P015N062P058(0)='1' AND  B( 3)='1' AND A( 1)='1' AND A(11)='0' )then
          cVar2S20S6P033P017P016nsss(0) <='1';
          else
          cVar2S20S6P033P017P016nsss(0) <='0';
          end if;
        if(cVar1S21S6N044P015N062N058(0)='1' AND  D(10)='1' AND E(11)='1' )then
          cVar2S21S6P061P059nsss(0) <='1';
          else
          cVar2S21S6P061P059nsss(0) <='0';
          end if;
        if(cVar1S22S6N044P015N062N058(0)='1' AND  D(10)='1' AND E(11)='0' AND A(10)='1' )then
          cVar2S22S6P061N059P018nsss(0) <='1';
          else
          cVar2S22S6P061N059P018nsss(0) <='0';
          end if;
        if(cVar1S23S6N044P015N062N058(0)='1' AND  D(10)='0' AND D( 7)='1' )then
          cVar2S23S6N061P040nsss(0) <='1';
          else
          cVar2S23S6N061P040nsss(0) <='0';
          end if;
        if(cVar1S24S6N044P015N062N058(0)='1' AND  D(10)='0' AND D( 7)='0' AND D( 9)='1' )then
          cVar2S24S6N061N040P065nsss(0) <='1';
          else
          cVar2S24S6N061N040P065nsss(0) <='0';
          end if;
        if(cVar1S2S7P050P027N048N009(0)='1' AND  A(15)='1' )then
          cVar2S2S7P008nsss(0) <='1';
          else
          cVar2S2S7P008nsss(0) <='0';
          end if;
        if(cVar1S3S7P050P027N048N009(0)='1' AND  A(15)='0' AND A( 4)='1' )then
          cVar2S3S7N008P011nsss(0) <='1';
          else
          cVar2S3S7N008P011nsss(0) <='0';
          end if;
        if(cVar1S5S7P050N027P052N008(0)='1' AND  B( 5)='1' )then
          cVar2S5S7P029nsss(0) <='1';
          else
          cVar2S5S7P029nsss(0) <='0';
          end if;
        if(cVar1S6S7P050N027P052N008(0)='1' AND  B( 5)='0' AND A(14)='1' )then
          cVar2S6S7N029P010nsss(0) <='1';
          else
          cVar2S6S7N029P010nsss(0) <='0';
          end if;
        if(cVar1S7S7P050N027P052N008(0)='1' AND  B( 5)='0' AND A(14)='0' AND A(16)='1' )then
          cVar2S7S7N029N010P006nsss(0) <='1';
          else
          cVar2S7S7N029N010P006nsss(0) <='0';
          end if;
        if(cVar1S8S7P050N027N052P048(0)='1' AND  B(16)='1' )then
          cVar2S8S7P026nsss(0) <='1';
          else
          cVar2S8S7P026nsss(0) <='0';
          end if;
        if(cVar1S9S7P050N027N052P048(0)='1' AND  B(16)='0' AND A( 2)='0' )then
          cVar2S9S7N026P015nsss(0) <='1';
          else
          cVar2S9S7N026P015nsss(0) <='0';
          end if;
        if(cVar1S10S7P050N027N052N048(0)='1' AND  D(11)='1' )then
          cVar2S10S7P057nsss(0) <='1';
          else
          cVar2S10S7P057nsss(0) <='0';
          end if;
        if(cVar1S13S7N050P044N023N004(0)='1' AND  A(16)='1' )then
          cVar2S13S7P006nsss(0) <='1';
          else
          cVar2S13S7P006nsss(0) <='0';
          end if;
        if(cVar1S14S7N050P044N023N004(0)='1' AND  A(16)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar2S14S7N006P007P025nsss(0) <='1';
          else
          cVar2S14S7N006P007P025nsss(0) <='0';
          end if;
        if(cVar1S15S7N050P044N023N004(0)='1' AND  A(16)='0' AND A( 6)='0' AND A(18)='1' )then
          cVar2S15S7N006N007P002nsss(0) <='1';
          else
          cVar2S15S7N006N007P002nsss(0) <='0';
          end if;
        if(cVar1S16S7N050N044P056P031(0)='1' AND  A( 3)='1' )then
          cVar2S16S7P013nsss(0) <='1';
          else
          cVar2S16S7P013nsss(0) <='0';
          end if;
        if(cVar1S17S7N050N044P056P031(0)='1' AND  A( 3)='0' AND E( 9)='0' )then
          cVar2S17S7N013P067nsss(0) <='1';
          else
          cVar2S17S7N013P067nsss(0) <='0';
          end if;
        if(cVar1S18S7N050N044P056N031(0)='1' AND  E( 9)='0' )then
          cVar2S18S7P067nsss(0) <='1';
          else
          cVar2S18S7P067nsss(0) <='0';
          end if;
        if(cVar1S19S7N050N044P056N031(0)='1' AND  E( 9)='1' AND D( 9)='1' )then
          cVar2S19S7P067P065nsss(0) <='1';
          else
          cVar2S19S7P067P065nsss(0) <='0';
          end if;
        if(cVar1S20S7N050N044N056P038(0)='1' AND  B( 9)='1' )then
          cVar2S20S7P021nsss(0) <='1';
          else
          cVar2S20S7P021nsss(0) <='0';
          end if;
        if(cVar1S21S7N050N044N056P038(0)='1' AND  B( 9)='0' AND B(19)='1' )then
          cVar2S21S7N021P020nsss(0) <='1';
          else
          cVar2S21S7N021P020nsss(0) <='0';
          end if;
        if(cVar1S22S7N050N044N056N038(0)='1' AND  E( 2)='1' AND E( 9)='0' )then
          cVar2S22S7P062P067nsss(0) <='1';
          else
          cVar2S22S7P062P067nsss(0) <='0';
          end if;
        if(cVar1S23S7N050N044N056N038(0)='1' AND  E( 2)='1' AND E( 9)='1' AND D( 9)='1' )then
          cVar2S23S7P062P067P065nsss(0) <='1';
          else
          cVar2S23S7P062P067P065nsss(0) <='0';
          end if;
        if(cVar1S24S7N050N044N056N038(0)='1' AND  E( 2)='0' AND E( 1)='1' AND D( 0)='1' )then
          cVar2S24S7N062P066P068nsss(0) <='1';
          else
          cVar2S24S7N062P066P068nsss(0) <='0';
          end if;
        if(cVar1S25S7N050N044N056N038(0)='1' AND  E( 2)='0' AND E( 1)='0' AND E(14)='1' )then
          cVar2S25S7N062N066P047nsss(0) <='1';
          else
          cVar2S25S7N062N066P047nsss(0) <='0';
          end if;
        if(cVar1S2S8P044P023N005N004(0)='1' AND  A( 2)='0' )then
          cVar2S2S8P015nsss(0) <='1';
          else
          cVar2S2S8P015nsss(0) <='0';
          end if;
        if(cVar1S5S8P044N023N004N006(0)='1' AND  A( 6)='1' )then
          cVar2S5S8P007nsss(0) <='1';
          else
          cVar2S5S8P007nsss(0) <='0';
          end if;
        if(cVar1S6S8P044N023N004N006(0)='1' AND  A( 6)='0' AND E( 7)='0' AND E( 6)='0' )then
          cVar2S6S8N007P042P046nsss(0) <='1';
          else
          cVar2S6S8N007P042P046nsss(0) <='0';
          end if;
        if(cVar1S7S8P044N023N004N006(0)='1' AND  A( 6)='0' AND E( 7)='1' AND A(18)='1' )then
          cVar2S7S8N007P042P002nsss(0) <='1';
          else
          cVar2S7S8N007P042P002nsss(0) <='0';
          end if;
        if(cVar1S9S8N044P050P027N009(0)='1' AND  D( 5)='1' )then
          cVar2S9S8P048nsss(0) <='1';
          else
          cVar2S9S8P048nsss(0) <='0';
          end if;
        if(cVar1S10S8N044P050P027N009(0)='1' AND  D( 5)='0' AND A(16)='1' )then
          cVar2S10S8N048P006nsss(0) <='1';
          else
          cVar2S10S8N048P006nsss(0) <='0';
          end if;
        if(cVar1S11S8N044P050P027N009(0)='1' AND  D( 5)='0' AND A(16)='0' AND A(15)='1' )then
          cVar2S11S8N048N006P008nsss(0) <='1';
          else
          cVar2S11S8N048N006P008nsss(0) <='0';
          end if;
        if(cVar1S12S8N044P050N027P026(0)='1' AND  A(15)='1' )then
          cVar2S12S8P008nsss(0) <='1';
          else
          cVar2S12S8P008nsss(0) <='0';
          end if;
        if(cVar1S13S8N044P050N027P026(0)='1' AND  A(15)='0' AND A(14)='1' )then
          cVar2S13S8N008P010nsss(0) <='1';
          else
          cVar2S13S8N008P010nsss(0) <='0';
          end if;
        if(cVar1S14S8N044P050N027P026(0)='1' AND  A(15)='0' AND A(14)='0' AND A(16)='1' )then
          cVar2S14S8N008N010P006nsss(0) <='1';
          else
          cVar2S14S8N008N010P006nsss(0) <='0';
          end if;
        if(cVar1S15S8N044P050N027N026(0)='1' AND  B( 5)='1' )then
          cVar2S15S8P029nsss(0) <='1';
          else
          cVar2S15S8P029nsss(0) <='0';
          end if;
        if(cVar1S16S8N044P050N027N026(0)='1' AND  B( 5)='0' AND A( 5)='0' )then
          cVar2S16S8N029P009nsss(0) <='1';
          else
          cVar2S16S8N029P009nsss(0) <='0';
          end if;
        if(cVar1S17S8N044N050P014P051(0)='1' AND  B(15)='1' AND E( 4)='0' )then
          cVar2S17S8P028P054nsss(0) <='1';
          else
          cVar2S17S8P028P054nsss(0) <='0';
          end if;
        if(cVar1S18S8N044N050P014P051(0)='1' AND  B(15)='0' AND A(15)='1' AND B(16)='1' )then
          cVar2S18S8N028P008P026nsss(0) <='1';
          else
          cVar2S18S8N028P008P026nsss(0) <='0';
          end if;
        if(cVar1S19S8N044N050P014P051(0)='1' AND  B(15)='0' AND A(15)='0' AND A( 5)='1' )then
          cVar2S19S8N028N008P009nsss(0) <='1';
          else
          cVar2S19S8N028N008P009nsss(0) <='0';
          end if;
        if(cVar1S20S8N044N050P014N051(0)='1' AND  B(18)='1' AND E(15)='1' )then
          cVar2S20S8P022P043nsss(0) <='1';
          else
          cVar2S20S8P022P043nsss(0) <='0';
          end if;
        if(cVar1S21S8N044N050P014N051(0)='1' AND  B(18)='1' AND E(15)='0' AND B( 0)='1' )then
          cVar2S21S8P022N043P039nsss(0) <='1';
          else
          cVar2S21S8P022N043P039nsss(0) <='0';
          end if;
        if(cVar1S22S8N044N050P014N051(0)='1' AND  B(18)='0' )then
          cVar2S22S8N022psss(0) <='1';
          else
          cVar2S22S8N022psss(0) <='0';
          end if;
        if(cVar1S23S8N044N050P014P032(0)='1' AND  D(10)='1' AND A( 3)='0' )then
          cVar2S23S8P061P013nsss(0) <='1';
          else
          cVar2S23S8P061P013nsss(0) <='0';
          end if;
        if(cVar1S24S8N044N050P014P032(0)='1' AND  D(10)='1' AND A( 3)='1' AND D( 0)='0' )then
          cVar2S24S8P061P013P068nsss(0) <='1';
          else
          cVar2S24S8P061P013P068nsss(0) <='0';
          end if;
        if(cVar1S25S8N044N050P014P032(0)='1' AND  D(10)='0' AND B(14)='0' )then
          cVar2S25S8N061P030nsss(0) <='1';
          else
          cVar2S25S8N061P030nsss(0) <='0';
          end if;
        if(cVar1S26S8N044N050P014N032(0)='1' AND  D( 9)='1' AND B(12)='1' )then
          cVar2S26S8P065P034nsss(0) <='1';
          else
          cVar2S26S8P065P034nsss(0) <='0';
          end if;
        if(cVar1S27S8N044N050P014N032(0)='1' AND  D( 9)='1' AND B(12)='0' AND E(10)='0' )then
          cVar2S27S8P065N034P063nsss(0) <='1';
          else
          cVar2S27S8P065N034P063nsss(0) <='0';
          end if;
        if(cVar1S28S8N044N050P014N032(0)='1' AND  D( 9)='0' AND E( 9)='0' AND A( 2)='1' )then
          cVar2S28S8N065P067P015nsss(0) <='1';
          else
          cVar2S28S8N065P067P015nsss(0) <='0';
          end if;
        if(cVar1S3S9P051N028N029P026(0)='1' AND  A(15)='1' AND A( 3)='0' )then
          cVar2S3S9P008P013nsss(0) <='1';
          else
          cVar2S3S9P008P013nsss(0) <='0';
          end if;
        if(cVar1S4S9P051N028N029P026(0)='1' AND  A(15)='0' AND A( 5)='1' )then
          cVar2S4S9N008P009nsss(0) <='1';
          else
          cVar2S4S9N008P009nsss(0) <='0';
          end if;
        if(cVar1S5S9P051N028N029P026(0)='1' AND  A(15)='0' AND A( 5)='0' AND A( 6)='1' )then
          cVar2S5S9N008N009P007nsss(0) <='1';
          else
          cVar2S5S9N008N009P007nsss(0) <='0';
          end if;
        if(cVar1S6S9P051N028N029N026(0)='1' AND  B( 6)='1' AND A( 5)='1' )then
          cVar2S6S9P027P009nsss(0) <='1';
          else
          cVar2S6S9P027P009nsss(0) <='0';
          end if;
        if(cVar1S7S9P051N028N029N026(0)='1' AND  B( 6)='0' AND D(11)='1' AND B(14)='1' )then
          cVar2S7S9N027P057P030nsss(0) <='1';
          else
          cVar2S7S9N027P057P030nsss(0) <='0';
          end if;
        if(cVar1S10S9N051P022N043N004(0)='1' AND  A(14)='0' AND B( 8)='0' )then
          cVar2S10S9P010P023nsss(0) <='1';
          else
          cVar2S10S9P010P023nsss(0) <='0';
          end if;
        if(cVar1S12S9N051N022P044N023(0)='1' AND  B( 7)='1' AND A(12)='0' )then
          cVar2S12S9P025P014nsss(0) <='1';
          else
          cVar2S12S9P025P014nsss(0) <='0';
          end if;
        if(cVar1S13S9N051N022P044N023(0)='1' AND  B( 7)='0' AND E(14)='1' )then
          cVar2S13S9N025P047nsss(0) <='1';
          else
          cVar2S13S9N025P047nsss(0) <='0';
          end if;
        if(cVar1S14S9N051N022P044N023(0)='1' AND  B( 7)='0' AND E(14)='0' AND A( 0)='0' )then
          cVar2S14S9N025N047P019nsss(0) <='1';
          else
          cVar2S14S9N025N047P019nsss(0) <='0';
          end if;
        if(cVar1S15S9N051N022N044P050(0)='1' AND  B( 6)='1' )then
          cVar2S15S9P027nsss(0) <='1';
          else
          cVar2S15S9P027nsss(0) <='0';
          end if;
        if(cVar1S16S9N051N022N044P050(0)='1' AND  B( 6)='0' AND B(16)='1' )then
          cVar2S16S9N027P026nsss(0) <='1';
          else
          cVar2S16S9N027P026nsss(0) <='0';
          end if;
        if(cVar1S17S9N051N022N044P050(0)='1' AND  B( 6)='0' AND B(16)='0' AND B( 5)='1' )then
          cVar2S17S9N027N026P029nsss(0) <='1';
          else
          cVar2S17S9N027N026P029nsss(0) <='0';
          end if;
        if(cVar1S18S9N051N022N044N050(0)='1' AND  B(10)='1' AND B( 9)='1' )then
          cVar2S18S9P038P021nsss(0) <='1';
          else
          cVar2S18S9P038P021nsss(0) <='0';
          end if;
        if(cVar1S19S9N051N022N044N050(0)='1' AND  B(10)='1' AND B( 9)='0' AND A(18)='1' )then
          cVar2S19S9P038N021P002nsss(0) <='1';
          else
          cVar2S19S9P038N021P002nsss(0) <='0';
          end if;
        if(cVar1S20S9N051N022N044N050(0)='1' AND  B(10)='0' AND A( 5)='0' AND D( 9)='1' )then
          cVar2S20S9N038P009P065nsss(0) <='1';
          else
          cVar2S20S9N038P009P065nsss(0) <='0';
          end if;
        if(cVar1S21S9N051N022N044N050(0)='1' AND  B(10)='0' AND A( 5)='1' AND E( 6)='1' )then
          cVar2S21S9N038P009P046nsss(0) <='1';
          else
          cVar2S21S9N038P009P046nsss(0) <='0';
          end if;
        if(cVar1S0S10P017P037P051P063(0)='1' AND  E( 9)='0' AND A(15)='1' )then
          cVar2S0S10P067P008nsss(0) <='1';
          else
          cVar2S0S10P067P008nsss(0) <='0';
          end if;
        if(cVar1S1S10P017P037P051P063(0)='1' AND  E( 9)='0' AND A(15)='0' AND E(14)='0' )then
          cVar2S1S10P067N008P047nsss(0) <='1';
          else
          cVar2S1S10P067N008P047nsss(0) <='0';
          end if;
        if(cVar1S2S10P017P037P051P063(0)='1' AND  E( 9)='1' AND A( 3)='1' )then
          cVar2S2S10P067P013nsss(0) <='1';
          else
          cVar2S2S10P067P013nsss(0) <='0';
          end if;
        if(cVar1S3S10P017P037N051P048(0)='1' AND  B( 6)='1' )then
          cVar2S3S10P027nsss(0) <='1';
          else
          cVar2S3S10P027nsss(0) <='0';
          end if;
        if(cVar1S4S10P017P037N051P048(0)='1' AND  B( 6)='0' AND B( 7)='1' )then
          cVar2S4S10N027P025nsss(0) <='1';
          else
          cVar2S4S10N027P025nsss(0) <='0';
          end if;
        if(cVar1S5S10P017P037N051P048(0)='1' AND  B( 6)='0' AND B( 7)='0' AND A(16)='1' )then
          cVar2S5S10N027N025P006nsss(0) <='1';
          else
          cVar2S5S10N027N025P006nsss(0) <='0';
          end if;
        if(cVar1S6S10P017P037N051N048(0)='1' AND  B(18)='1' AND E(15)='1' )then
          cVar2S6S10P022P043nsss(0) <='1';
          else
          cVar2S6S10P022P043nsss(0) <='0';
          end if;
        if(cVar1S7S10P017P037N051N048(0)='1' AND  B(18)='1' AND E(15)='0' AND A(17)='1' )then
          cVar2S7S10P022N043P004nsss(0) <='1';
          else
          cVar2S7S10P022N043P004nsss(0) <='0';
          end if;
        if(cVar1S8S10P017P037N051N048(0)='1' AND  B(18)='0' )then
          cVar2S8S10N022psss(0) <='1';
          else
          cVar2S8S10N022psss(0) <='0';
          end if;
        if(cVar1S9S10P017P037P019P064(0)='1' AND  E( 1)='1' AND A(10)='0' AND A(14)='0' )then
          cVar2S9S10P066P018P010nsss(0) <='1';
          else
          cVar2S9S10P066P018P010nsss(0) <='0';
          end if;
        if(cVar1S10S10P017P037P019P064(0)='1' AND  E( 1)='1' AND A(10)='1' AND B( 3)='0' )then
          cVar2S10S10P066P018P033nsss(0) <='1';
          else
          cVar2S10S10P066P018P033nsss(0) <='0';
          end if;
        if(cVar1S11S10P017P037P019P064(0)='1' AND  E( 1)='0' AND D( 8)='1' )then
          cVar2S11S10N066P069nsss(0) <='1';
          else
          cVar2S11S10N066P069nsss(0) <='0';
          end if;
        if(cVar1S12S10P017P037P019P064(0)='1' AND  D( 0)='0' AND E( 1)='1' )then
          cVar2S12S10P068P066nsss(0) <='1';
          else
          cVar2S12S10P068P066nsss(0) <='0';
          end if;
        if(cVar1S13S10P017P037P019P064(0)='1' AND  D( 0)='1' AND D( 9)='0' AND A(12)='1' )then
          cVar2S13S10P068P065P014nsss(0) <='1';
          else
          cVar2S13S10P068P065P014nsss(0) <='0';
          end if;
        if(cVar1S14S10P017P037N019P063(0)='1' AND  D( 0)='1' AND E( 9)='0' AND A( 2)='1' )then
          cVar2S14S10P068P067P015nsss(0) <='1';
          else
          cVar2S14S10P068P067P015nsss(0) <='0';
          end if;
        if(cVar1S15S10P017P037N019P063(0)='1' AND  A(11)='1' AND A(13)='0' AND B(12)='1' )then
          cVar2S15S10P016P012P034nsss(0) <='1';
          else
          cVar2S15S10P016P012P034nsss(0) <='0';
          end if;
        if(cVar1S16S10P017P064P019P068(0)='1' AND  A( 8)='0' AND B( 2)='1' )then
          cVar2S16S10P003P035nsss(0) <='1';
          else
          cVar2S16S10P003P035nsss(0) <='0';
          end if;
        if(cVar1S17S10P017P064P019P068(0)='1' AND  A( 8)='0' AND B( 2)='0' AND B( 1)='1' )then
          cVar2S17S10P003N035P037nsss(0) <='1';
          else
          cVar2S17S10P003N035P037nsss(0) <='0';
          end if;
        if(cVar1S18S10P017P064P019P068(0)='1' AND  E( 1)='1' AND E( 9)='0' AND A( 2)='1' )then
          cVar2S18S10P066P067P015nsss(0) <='1';
          else
          cVar2S18S10P066P067P015nsss(0) <='0';
          end if;
        if(cVar1S19S10P017P064P019P015(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S19S10P016P018nsss(0) <='1';
          else
          cVar2S19S10P016P018nsss(0) <='0';
          end if;
        if(cVar1S20S10P017P064P019P015(0)='1' AND  A(11)='0' AND A(10)='0' AND B( 1)='0' )then
          cVar2S20S10P016N018P037nsss(0) <='1';
          else
          cVar2S20S10P016N018P037nsss(0) <='0';
          end if;
        if(cVar1S21S10P017P064P019P015(0)='1' AND  A(11)='1' AND D( 0)='1' )then
          cVar2S21S10P016P068nsss(0) <='1';
          else
          cVar2S21S10P016P068nsss(0) <='0';
          end if;
        if(cVar1S22S10P017P064P019N015(0)='1' AND  A( 8)='0' AND B( 2)='1' AND E( 9)='0' )then
          cVar2S22S10P003P035P067nsss(0) <='1';
          else
          cVar2S22S10P003P035P067nsss(0) <='0';
          end if;
        if(cVar1S23S10P017N064P015P065(0)='1' AND  E( 9)='0' AND E(13)='1' )then
          cVar2S23S10P067P051nsss(0) <='1';
          else
          cVar2S23S10P067P051nsss(0) <='0';
          end if;
        if(cVar1S24S10P017N064P015P065(0)='1' AND  E( 9)='0' AND E(13)='0' AND E(15)='0' )then
          cVar2S24S10P067N051P043nsss(0) <='1';
          else
          cVar2S24S10P067N051P043nsss(0) <='0';
          end if;
        if(cVar1S25S10P017N064P015P065(0)='1' AND  E( 9)='1' AND D( 8)='1' AND A( 4)='0' )then
          cVar2S25S10P067P069P011nsss(0) <='1';
          else
          cVar2S25S10P067P069P011nsss(0) <='0';
          end if;
        if(cVar1S26S10P017N064P015P065(0)='1' AND  B(12)='1' AND E( 1)='0' AND A( 0)='0' )then
          cVar2S26S10P034P066P019nsss(0) <='1';
          else
          cVar2S26S10P034P066P019nsss(0) <='0';
          end if;
        if(cVar1S27S10P017N064N015P037(0)='1' AND  E( 1)='1' AND A(13)='0' AND A(15)='0' )then
          cVar2S27S10P066P012P008nsss(0) <='1';
          else
          cVar2S27S10P066P012P008nsss(0) <='0';
          end if;
        if(cVar1S28S10P017N064N015P037(0)='1' AND  E( 1)='1' AND A(13)='1' AND A(10)='0' )then
          cVar2S28S10P066P012P018nsss(0) <='1';
          else
          cVar2S28S10P066P012P018nsss(0) <='0';
          end if;
        if(cVar1S29S10P017N064N015P037(0)='1' AND  E( 1)='0' AND D( 8)='1' AND A(11)='0' )then
          cVar2S29S10N066P069P016nsss(0) <='1';
          else
          cVar2S29S10N066P069P016nsss(0) <='0';
          end if;
        if(cVar1S30S10P017N064N015P037(0)='1' AND  E( 1)='0' AND D( 8)='0' AND A(15)='1' )then
          cVar2S30S10N066N069P008nsss(0) <='1';
          else
          cVar2S30S10N066N069P008nsss(0) <='0';
          end if;
        if(cVar1S31S10P017N064N015N037(0)='1' AND  B(12)='1' AND E(10)='1' AND A(13)='0' )then
          cVar2S31S10P034P063P012nsss(0) <='1';
          else
          cVar2S31S10P034P063P012nsss(0) <='0';
          end if;
        if(cVar1S32S10P017N064N015N037(0)='1' AND  B(12)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar2S32S10N034P031P013nsss(0) <='1';
          else
          cVar2S32S10N034P031P013nsss(0) <='0';
          end if;
        if(cVar1S33S10P017N064N015N037(0)='1' AND  B(12)='0' AND B( 4)='0' AND B(10)='1' )then
          cVar2S33S10N034N031P038nsss(0) <='1';
          else
          cVar2S33S10N034N031P038nsss(0) <='0';
          end if;
        if(cVar1S2S11P048P025N007N006(0)='1' AND  A( 5)='1' )then
          cVar2S2S11P009nsss(0) <='1';
          else
          cVar2S2S11P009nsss(0) <='0';
          end if;
        if(cVar1S3S11P048P025N007N006(0)='1' AND  A( 5)='0' AND A( 7)='1' )then
          cVar2S3S11N009P005nsss(0) <='1';
          else
          cVar2S3S11N009P005nsss(0) <='0';
          end if;
        if(cVar1S4S11P048P025N007N006(0)='1' AND  A( 5)='0' AND A( 7)='0' AND A(15)='1' )then
          cVar2S4S11N009N005P008nsss(0) <='1';
          else
          cVar2S4S11N009N005P008nsss(0) <='0';
          end if;
        if(cVar1S5S11P048N025P027P011(0)='1' AND  A( 5)='1' )then
          cVar2S5S11P009nsss(0) <='1';
          else
          cVar2S5S11P009nsss(0) <='0';
          end if;
        if(cVar1S6S11P048N025P027P011(0)='1' AND  A( 5)='0' AND A( 6)='1' )then
          cVar2S6S11N009P007nsss(0) <='1';
          else
          cVar2S6S11N009P007nsss(0) <='0';
          end if;
        if(cVar1S7S11P048N025P027P011(0)='1' AND  A( 5)='0' AND A( 6)='0' AND A(15)='1' )then
          cVar2S7S11N009N007P008nsss(0) <='1';
          else
          cVar2S7S11N009N007P008nsss(0) <='0';
          end if;
        if(cVar1S8S11P048N025P027P011(0)='1' AND  E( 6)='0' )then
          cVar2S8S11P046nsss(0) <='1';
          else
          cVar2S8S11P046nsss(0) <='0';
          end if;
        if(cVar1S9S11P048N025N027P007(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S9S11P006P024nsss(0) <='1';
          else
          cVar2S9S11P006P024nsss(0) <='0';
          end if;
        if(cVar1S10S11P048N025N027P007(0)='1' AND  A(16)='1' AND B(17)='0' AND B(16)='1' )then
          cVar2S10S11P006N024P026nsss(0) <='1';
          else
          cVar2S10S11P006N024P026nsss(0) <='0';
          end if;
        if(cVar1S11S11P048N025N027P007(0)='1' AND  A(16)='0' AND B(16)='1' AND A(15)='1' )then
          cVar2S11S11N006P026P008nsss(0) <='1';
          else
          cVar2S11S11N006P026P008nsss(0) <='0';
          end if;
        if(cVar1S12S11P048N025N027P007(0)='1' AND  A(16)='0' AND B(16)='0' AND E( 3)='1' )then
          cVar2S12S11N006N026P058nsss(0) <='1';
          else
          cVar2S12S11N006N026P058nsss(0) <='0';
          end if;
        if(cVar1S15S11N048P051N028N029(0)='1' AND  B(16)='1' AND A(15)='1' )then
          cVar2S15S11P026P008nsss(0) <='1';
          else
          cVar2S15S11P026P008nsss(0) <='0';
          end if;
        if(cVar1S16S11N048P051N028N029(0)='1' AND  B(16)='1' AND A(15)='0' AND E(14)='0' )then
          cVar2S16S11P026N008P047nsss(0) <='1';
          else
          cVar2S16S11P026N008P047nsss(0) <='0';
          end if;
        if(cVar1S17S11N048P051N028N029(0)='1' AND  B(16)='0' AND B( 6)='1' )then
          cVar2S17S11N026P027nsss(0) <='1';
          else
          cVar2S17S11N026P027nsss(0) <='0';
          end if;
        if(cVar1S18S11N048N051P022P043(0)='1' AND  B( 2)='0' )then
          cVar2S18S11P035nsss(0) <='1';
          else
          cVar2S18S11P035nsss(0) <='0';
          end if;
        if(cVar1S19S11N048N051P022N043(0)='1' AND  D( 6)='1' )then
          cVar2S19S11P044nsss(0) <='1';
          else
          cVar2S19S11P044nsss(0) <='0';
          end if;
        if(cVar1S20S11N048N051P022N043(0)='1' AND  D( 6)='0' AND D( 7)='1' )then
          cVar2S20S11N044P040nsss(0) <='1';
          else
          cVar2S20S11N044P040nsss(0) <='0';
          end if;
        if(cVar1S21S11N048N051P022N043(0)='1' AND  D( 6)='0' AND D( 7)='0' AND A(12)='0' )then
          cVar2S21S11N044N040P014nsss(0) <='1';
          else
          cVar2S21S11N044N040P014nsss(0) <='0';
          end if;
        if(cVar1S22S11N048N051N022P023(0)='1' AND  E( 7)='1' AND A(15)='0' )then
          cVar2S22S11P042P008nsss(0) <='1';
          else
          cVar2S22S11P042P008nsss(0) <='0';
          end if;
        if(cVar1S23S11N048N051N022P023(0)='1' AND  E( 7)='0' AND E(15)='1' )then
          cVar2S23S11N042P043nsss(0) <='1';
          else
          cVar2S23S11N042P043nsss(0) <='0';
          end if;
        if(cVar1S24S11N048N051N022P023(0)='1' AND  E( 7)='0' AND E(15)='0' AND D( 1)='1' )then
          cVar2S24S11N042N043P064nsss(0) <='1';
          else
          cVar2S24S11N042N043P064nsss(0) <='0';
          end if;
        if(cVar1S25S11N048N051N022N023(0)='1' AND  E(15)='0' AND A( 6)='0' AND B( 4)='1' )then
          cVar2S25S11P043P007P031nsss(0) <='1';
          else
          cVar2S25S11P043P007P031nsss(0) <='0';
          end if;
        if(cVar1S26S11N048N051N022N023(0)='1' AND  E(15)='0' AND A( 6)='1' AND E(14)='1' )then
          cVar2S26S11P043P007P047nsss(0) <='1';
          else
          cVar2S26S11P043P007P047nsss(0) <='0';
          end if;
        if(cVar1S27S11N048N051N022N023(0)='1' AND  E(15)='1' AND B(17)='1' )then
          cVar2S27S11P043P024nsss(0) <='1';
          else
          cVar2S27S11P043P024nsss(0) <='0';
          end if;
        if(cVar1S28S11N048N051N022N023(0)='1' AND  E(15)='1' AND B(17)='0' AND B( 7)='1' )then
          cVar2S28S11P043N024P025nsss(0) <='1';
          else
          cVar2S28S11P043N024P025nsss(0) <='0';
          end if;
        if(cVar1S2S12P048P025N007N006(0)='1' AND  A( 5)='1' )then
          cVar2S2S12P009nsss(0) <='1';
          else
          cVar2S2S12P009nsss(0) <='0';
          end if;
        if(cVar1S3S12P048P025N007N006(0)='1' AND  A( 5)='0' AND A( 7)='1' )then
          cVar2S3S12N009P005nsss(0) <='1';
          else
          cVar2S3S12N009P005nsss(0) <='0';
          end if;
        if(cVar1S4S12P048P025N007N006(0)='1' AND  A( 5)='0' AND A( 7)='0' AND A(15)='1' )then
          cVar2S4S12N009N005P008nsss(0) <='1';
          else
          cVar2S4S12N009N005P008nsss(0) <='0';
          end if;
        if(cVar1S6S12P048N025N027P067(0)='1' AND  B(17)='1' )then
          cVar2S6S12P024nsss(0) <='1';
          else
          cVar2S6S12P024nsss(0) <='0';
          end if;
        if(cVar1S7S12P048N025N027P067(0)='1' AND  B(17)='0' AND B(16)='1' )then
          cVar2S7S12N024P026nsss(0) <='1';
          else
          cVar2S7S12N024P026nsss(0) <='0';
          end if;
        if(cVar1S8S12P048N025N027P067(0)='1' AND  B(17)='0' AND B(16)='0' AND A(15)='0' )then
          cVar2S8S12N024N026P008nsss(0) <='1';
          else
          cVar2S8S12N024N026P008nsss(0) <='0';
          end if;
        if(cVar1S9S12N048P001P051P013(0)='1' AND  A(15)='1' AND B(16)='1' )then
          cVar2S9S12P008P026nsss(0) <='1';
          else
          cVar2S9S12P008P026nsss(0) <='0';
          end if;
        if(cVar1S10S12N048P001P051P013(0)='1' AND  A(15)='1' AND B(16)='0' AND B(15)='1' )then
          cVar2S10S12P008N026P028nsss(0) <='1';
          else
          cVar2S10S12P008N026P028nsss(0) <='0';
          end if;
        if(cVar1S11S12N048P001P051P013(0)='1' AND  A(15)='0' )then
          cVar2S11S12N008psss(0) <='1';
          else
          cVar2S11S12N008psss(0) <='0';
          end if;
        if(cVar1S12S12N048P001P051P013(0)='1' AND  A( 8)='0' AND A(11)='0' )then
          cVar2S12S12P003P016nsss(0) <='1';
          else
          cVar2S12S12P003P016nsss(0) <='0';
          end if;
        if(cVar1S13S12N048P001P051P013(0)='1' AND  A( 8)='0' AND A(11)='1' AND A(10)='1' )then
          cVar2S13S12P003P016P018nsss(0) <='1';
          else
          cVar2S13S12P003P016P018nsss(0) <='0';
          end if;
        if(cVar1S14S12N048P001N051P008(0)='1' AND  B(16)='0' )then
          cVar2S14S12P026nsss(0) <='1';
          else
          cVar2S14S12P026nsss(0) <='0';
          end if;
        if(cVar1S15S12N048P001N051P008(0)='1' AND  B(16)='1' AND D(13)='1' )then
          cVar2S15S12P026P049nsss(0) <='1';
          else
          cVar2S15S12P026P049nsss(0) <='0';
          end if;
        if(cVar1S16S12N048P001N051P008(0)='1' AND  E(14)='1' AND B(16)='1' )then
          cVar2S16S12P047P026nsss(0) <='1';
          else
          cVar2S16S12P047P026nsss(0) <='0';
          end if;
        if(cVar1S17S12N048P001N051P008(0)='1' AND  E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar2S17S12P047N026P024nsss(0) <='1';
          else
          cVar2S17S12P047N026P024nsss(0) <='0';
          end if;
        if(cVar1S18S12N048P001N051P008(0)='1' AND  E(14)='0' AND E( 5)='1' AND A( 4)='0' )then
          cVar2S18S12N047P050P011nsss(0) <='1';
          else
          cVar2S18S12N047P050P011nsss(0) <='0';
          end if;
        if(cVar1S20S12N048P001N041P017(0)='1' AND  B( 3)='0' AND A(14)='1' )then
          cVar2S20S12P033P010nsss(0) <='1';
          else
          cVar2S20S12P033P010nsss(0) <='0';
          end if;
        if(cVar1S21S12N048P001N041P017(0)='1' AND  B( 3)='0' AND A(14)='0' AND E( 1)='0' )then
          cVar2S21S12P033N010P066nsss(0) <='1';
          else
          cVar2S21S12P033N010P066nsss(0) <='0';
          end if;
        if(cVar1S22S12N048P001N041N017(0)='1' AND  A( 2)='1' AND A( 3)='0' AND A(10)='1' )then
          cVar2S22S12P015P013P018nsss(0) <='1';
          else
          cVar2S22S12P015P013P018nsss(0) <='0';
          end if;
        if(cVar1S3S13P048N025P027P011(0)='1' AND  E( 5)='1' )then
          cVar2S3S13P050nsss(0) <='1';
          else
          cVar2S3S13P050nsss(0) <='0';
          end if;
        if(cVar1S4S13P048N025N027P007(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S4S13P006P024nsss(0) <='1';
          else
          cVar2S4S13P006P024nsss(0) <='0';
          end if;
        if(cVar1S5S13P048N025N027P007(0)='1' AND  A(16)='1' AND B(17)='0' AND B(16)='1' )then
          cVar2S5S13P006N024P026nsss(0) <='1';
          else
          cVar2S5S13P006N024P026nsss(0) <='0';
          end if;
        if(cVar1S6S13P048N025N027P007(0)='1' AND  A(16)='0' AND A( 1)='0' AND B(16)='1' )then
          cVar2S6S13N006P017P026nsss(0) <='1';
          else
          cVar2S6S13N006P017P026nsss(0) <='0';
          end if;
        if(cVar1S7S13P048N025N027P007(0)='1' AND  A(16)='0' AND A( 1)='1' AND D( 4)='1' )then
          cVar2S7S13N006P017P052nsss(0) <='1';
          else
          cVar2S7S13N006P017P052nsss(0) <='0';
          end if;
        if(cVar1S8S13N048P051P008P013(0)='1' AND  B(15)='1' )then
          cVar2S8S13P028nsss(0) <='1';
          else
          cVar2S8S13P028nsss(0) <='0';
          end if;
        if(cVar1S9S13N048P051P008P013(0)='1' AND  B(15)='0' AND B(16)='1' )then
          cVar2S9S13N028P026nsss(0) <='1';
          else
          cVar2S9S13N028P026nsss(0) <='0';
          end if;
        if(cVar1S10S13N048P051N008P028(0)='1' AND  A(14)='1' AND A(11)='0' AND E( 4)='0' )then
          cVar2S10S13P010P016P054nsss(0) <='1';
          else
          cVar2S10S13P010P016P054nsss(0) <='0';
          end if;
        if(cVar1S11S13N048P051N008P028(0)='1' AND  A(14)='1' AND A(11)='1' )then
          cVar2S11S13P010P016psss(0) <='1';
          else
          cVar2S11S13P010P016psss(0) <='0';
          end if;
        if(cVar1S12S13N048P051N008P028(0)='1' AND  A(14)='0' AND A( 4)='1' )then
          cVar2S12S13N010P011nsss(0) <='1';
          else
          cVar2S12S13N010P011nsss(0) <='0';
          end if;
        if(cVar1S13S13N048P051N008P028(0)='1' AND  A(14)='0' AND A( 4)='0' AND A( 5)='1' )then
          cVar2S13S13N010N011P009nsss(0) <='1';
          else
          cVar2S13S13N010N011P009nsss(0) <='0';
          end if;
        if(cVar1S14S13N048P051N008N028(0)='1' AND  B( 5)='1' AND A( 4)='1' )then
          cVar2S14S13P029P011nsss(0) <='1';
          else
          cVar2S14S13P029P011nsss(0) <='0';
          end if;
        if(cVar1S15S13N048P051N008N028(0)='1' AND  B( 5)='1' AND A( 4)='0' AND A( 5)='1' )then
          cVar2S15S13P029N011P009nsss(0) <='1';
          else
          cVar2S15S13P029N011P009nsss(0) <='0';
          end if;
        if(cVar1S16S13N048P051N008N028(0)='1' AND  B( 5)='0' AND A( 5)='1' AND A( 4)='0' )then
          cVar2S16S13N029P009P011nsss(0) <='1';
          else
          cVar2S16S13N029P009P011nsss(0) <='0';
          end if;
        if(cVar1S18S13N048N051P038N021(0)='1' AND  A(19)='1' )then
          cVar2S18S13P000nsss(0) <='1';
          else
          cVar2S18S13P000nsss(0) <='0';
          end if;
        if(cVar1S19S13N048N051P038N021(0)='1' AND  A(19)='0' AND B(19)='1' AND A(18)='1' )then
          cVar2S19S13N000P020P002nsss(0) <='1';
          else
          cVar2S19S13N000P020P002nsss(0) <='0';
          end if;
        if(cVar1S20S13N048N051P038N021(0)='1' AND  A(19)='0' AND B(19)='0' AND B( 8)='1' )then
          cVar2S20S13N000N020P023nsss(0) <='1';
          else
          cVar2S20S13N000N020P023nsss(0) <='0';
          end if;
        if(cVar1S21S13N048N051N038P061(0)='1' AND  B(13)='1' AND E( 1)='0' AND A(17)='0' )then
          cVar2S21S13P032P066P004nsss(0) <='1';
          else
          cVar2S21S13P032P066P004nsss(0) <='0';
          end if;
        if(cVar1S22S13N048N051N038P061(0)='1' AND  B(13)='1' AND E( 1)='1' AND A(12)='1' )then
          cVar2S22S13P032P066P014nsss(0) <='1';
          else
          cVar2S22S13P032P066P014nsss(0) <='0';
          end if;
        if(cVar1S23S13N048N051N038P061(0)='1' AND  B(13)='0' AND B(14)='1' AND A(13)='1' )then
          cVar2S23S13N032P030P012nsss(0) <='1';
          else
          cVar2S23S13N032P030P012nsss(0) <='0';
          end if;
        if(cVar1S24S13N048N051N038N061(0)='1' AND  E(12)='1' AND B(14)='1' AND B( 2)='0' )then
          cVar2S24S13P055P030P035nsss(0) <='1';
          else
          cVar2S24S13P055P030P035nsss(0) <='0';
          end if;
        if(cVar1S25S13N048N051N038N061(0)='1' AND  E(12)='1' AND B(14)='0' AND B(15)='1' )then
          cVar2S25S13P055N030P028nsss(0) <='1';
          else
          cVar2S25S13P055N030P028nsss(0) <='0';
          end if;
        if(cVar1S26S13N048N051N038N061(0)='1' AND  E(12)='0' AND B(18)='1' AND E(15)='1' )then
          cVar2S26S13N055P022P043nsss(0) <='1';
          else
          cVar2S26S13N055P022P043nsss(0) <='0';
          end if;
        if(cVar1S27S13N048N051N038N061(0)='1' AND  E(12)='0' AND B(18)='0' AND A( 1)='1' )then
          cVar2S27S13N055N022P017nsss(0) <='1';
          else
          cVar2S27S13N055N022P017nsss(0) <='0';
          end if;
        if(cVar1S1S14P017P048N025P027(0)='1' AND  A( 5)='1' )then
          cVar2S1S14P009nsss(0) <='1';
          else
          cVar2S1S14P009nsss(0) <='0';
          end if;
        if(cVar1S2S14P017P048N025P027(0)='1' AND  A( 5)='0' AND A( 6)='1' )then
          cVar2S2S14N009P007nsss(0) <='1';
          else
          cVar2S2S14N009P007nsss(0) <='0';
          end if;
        if(cVar1S3S14P017P048N025P027(0)='1' AND  A( 5)='0' AND A( 6)='0' AND A(15)='1' )then
          cVar2S3S14N009N007P008nsss(0) <='1';
          else
          cVar2S3S14N009N007P008nsss(0) <='0';
          end if;
        if(cVar1S4S14P017P048N025N027(0)='1' AND  A( 6)='0' AND A( 4)='0' AND B( 1)='0' )then
          cVar2S4S14P007P011P037nsss(0) <='1';
          else
          cVar2S4S14P007P011P037nsss(0) <='0';
          end if;
        if(cVar1S5S14P017P048N025N027(0)='1' AND  A( 6)='0' AND A( 4)='1' AND E( 5)='1' )then
          cVar2S5S14P007P011P050nsss(0) <='1';
          else
          cVar2S5S14P007P011P050nsss(0) <='0';
          end if;
        if(cVar1S7S14P017N048P044N023(0)='1' AND  B(18)='1' AND A(16)='1' )then
          cVar2S7S14P022P006nsss(0) <='1';
          else
          cVar2S7S14P022P006nsss(0) <='0';
          end if;
        if(cVar1S8S14P017N048P044N023(0)='1' AND  B(18)='1' AND A(16)='0' AND A(17)='1' )then
          cVar2S8S14P022N006P004nsss(0) <='1';
          else
          cVar2S8S14P022N006P004nsss(0) <='0';
          end if;
        if(cVar1S9S14P017N048P044N023(0)='1' AND  B(18)='0' AND B( 7)='1' )then
          cVar2S9S14N022P025nsss(0) <='1';
          else
          cVar2S9S14N022P025nsss(0) <='0';
          end if;
        if(cVar1S10S14P017N048P044N023(0)='1' AND  B(18)='0' AND B( 7)='0' AND E( 3)='1' )then
          cVar2S10S14N022N025P058nsss(0) <='1';
          else
          cVar2S10S14N022N025P058nsss(0) <='0';
          end if;
        if(cVar1S11S14P017N048N044P038(0)='1' AND  B( 9)='1' )then
          cVar2S11S14P021nsss(0) <='1';
          else
          cVar2S11S14P021nsss(0) <='0';
          end if;
        if(cVar1S12S14P017N048N044P038(0)='1' AND  B( 9)='0' AND B(19)='1' )then
          cVar2S12S14N021P020nsss(0) <='1';
          else
          cVar2S12S14N021P020nsss(0) <='0';
          end if;
        if(cVar1S13S14P017N048N044P038(0)='1' AND  B( 9)='0' AND B(19)='0' AND A( 3)='0' )then
          cVar2S13S14N021N020P013nsss(0) <='1';
          else
          cVar2S13S14N021N020P013nsss(0) <='0';
          end if;
        if(cVar1S14S14P017N048N044N038(0)='1' AND  A( 8)='0' AND E( 6)='0' )then
          cVar2S14S14P003P046nsss(0) <='1';
          else
          cVar2S14S14P003P046nsss(0) <='0';
          end if;
        if(cVar1S15S14P017N048N044N038(0)='1' AND  A( 8)='1' AND B( 0)='1' )then
          cVar2S15S14P003P039nsss(0) <='1';
          else
          cVar2S15S14P003P039nsss(0) <='0';
          end if;
        if(cVar1S16S14P017P064P019P009(0)='1' AND  B( 2)='1' AND D( 0)='0' AND A(13)='0' )then
          cVar2S16S14P035P068P012nsss(0) <='1';
          else
          cVar2S16S14P035P068P012nsss(0) <='0';
          end if;
        if(cVar1S17S14P017P064P019P009(0)='1' AND  B( 2)='1' AND D( 0)='1' AND A(10)='1' )then
          cVar2S17S14P035P068P018nsss(0) <='1';
          else
          cVar2S17S14P035P068P018nsss(0) <='0';
          end if;
        if(cVar1S18S14P017P064P019P009(0)='1' AND  B( 2)='0' AND A( 8)='0' AND A( 4)='0' )then
          cVar2S18S14N035P003P011nsss(0) <='1';
          else
          cVar2S18S14N035P003P011nsss(0) <='0';
          end if;
        if(cVar1S20S14P017P064P019N050(0)='1' AND  D( 3)='1' )then
          cVar2S20S14P056nsss(0) <='1';
          else
          cVar2S20S14P056nsss(0) <='0';
          end if;
        if(cVar1S21S14P017P064P019N050(0)='1' AND  D( 3)='0' AND A( 2)='1' AND A(15)='1' )then
          cVar2S21S14N056P015P008nsss(0) <='1';
          else
          cVar2S21S14N056P015P008nsss(0) <='0';
          end if;
        if(cVar1S22S14P017N064P061P003(0)='1' AND  A( 0)='0' AND E(11)='1' )then
          cVar2S22S14P019P059nsss(0) <='1';
          else
          cVar2S22S14P019P059nsss(0) <='0';
          end if;
        if(cVar1S23S14P017N064P061P003(0)='1' AND  A( 0)='0' AND E(11)='0' AND E(10)='1' )then
          cVar2S23S14P019N059P063nsss(0) <='1';
          else
          cVar2S23S14P019N059P063nsss(0) <='0';
          end if;
        if(cVar1S24S14P017N064P061P003(0)='1' AND  A( 0)='1' AND A(12)='1' AND A(11)='0' )then
          cVar2S24S14P019P014P016nsss(0) <='1';
          else
          cVar2S24S14P019P014P016nsss(0) <='0';
          end if;
        if(cVar1S25S14P017N064P061P003(0)='1' AND  A( 0)='1' AND A(12)='0' AND A(13)='1' )then
          cVar2S25S14P019N014P012nsss(0) <='1';
          else
          cVar2S25S14P019N014P012nsss(0) <='0';
          end if;
        if(cVar1S26S14P017N064N061P051(0)='1' AND  B(15)='1' )then
          cVar2S26S14P028nsss(0) <='1';
          else
          cVar2S26S14P028nsss(0) <='0';
          end if;
        if(cVar1S27S14P017N064N061P051(0)='1' AND  B(15)='0' AND A(15)='1' )then
          cVar2S27S14N028P008nsss(0) <='1';
          else
          cVar2S27S14N028P008nsss(0) <='0';
          end if;
        if(cVar1S28S14P017N064N061P051(0)='1' AND  B(15)='0' AND A(15)='0' AND B( 5)='1' )then
          cVar2S28S14N028N008P029nsss(0) <='1';
          else
          cVar2S28S14N028N008P029nsss(0) <='0';
          end if;
        if(cVar1S29S14P017N064N061N051(0)='1' AND  E(12)='1' AND B( 5)='0' AND B( 4)='0' )then
          cVar2S29S14P055P029P031nsss(0) <='1';
          else
          cVar2S29S14P055P029P031nsss(0) <='0';
          end if;
        if(cVar1S30S14P017N064N061N051(0)='1' AND  E(12)='0' AND D( 5)='1' AND A( 6)='1' )then
          cVar2S30S14N055P048P007nsss(0) <='1';
          else
          cVar2S30S14N055P048P007nsss(0) <='0';
          end if;
        if(cVar1S2S15P044P023N005N004(0)='1' AND  A( 6)='1' )then
          cVar2S2S15P007nsss(0) <='1';
          else
          cVar2S2S15P007nsss(0) <='0';
          end if;
        if(cVar1S3S15P044P023N005N004(0)='1' AND  A( 6)='0' AND A(16)='1' )then
          cVar2S3S15N007P006nsss(0) <='1';
          else
          cVar2S3S15N007P006nsss(0) <='0';
          end if;
        if(cVar1S5S15P044N023N022P025(0)='1' AND  A( 6)='1' )then
          cVar2S5S15P007nsss(0) <='1';
          else
          cVar2S5S15P007nsss(0) <='0';
          end if;
        if(cVar1S6S15P044N023N022P025(0)='1' AND  A( 6)='0' AND A(16)='1' )then
          cVar2S6S15N007P006nsss(0) <='1';
          else
          cVar2S6S15N007P006nsss(0) <='0';
          end if;
        if(cVar1S7S15P044N023N022P025(0)='1' AND  A( 6)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S7S15N007N006P005nsss(0) <='1';
          else
          cVar2S7S15N007N006P005nsss(0) <='0';
          end if;
        if(cVar1S8S15P044N023N022N025(0)='1' AND  E( 7)='0' )then
          cVar2S8S15P042nsss(0) <='1';
          else
          cVar2S8S15P042nsss(0) <='0';
          end if;
        if(cVar1S9S15P044N023N022N025(0)='1' AND  E( 7)='1' AND A(10)='0' AND A( 1)='0' )then
          cVar2S9S15P042P018P017nsss(0) <='1';
          else
          cVar2S9S15P042P018P017nsss(0) <='0';
          end if;
        if(cVar1S11S15N044P048P025N007(0)='1' AND  A(16)='1' )then
          cVar2S11S15P006nsss(0) <='1';
          else
          cVar2S11S15P006nsss(0) <='0';
          end if;
        if(cVar1S12S15N044P048P025N007(0)='1' AND  A(16)='0' AND A( 5)='1' )then
          cVar2S12S15N006P009nsss(0) <='1';
          else
          cVar2S12S15N006P009nsss(0) <='0';
          end if;
        if(cVar1S13S15N044P048P025N007(0)='1' AND  A(16)='0' AND A( 5)='0' AND A(15)='1' )then
          cVar2S13S15N006N009P008nsss(0) <='1';
          else
          cVar2S13S15N006N009P008nsss(0) <='0';
          end if;
        if(cVar1S14S15N044P048N025P027(0)='1' AND  D( 4)='0' AND E( 5)='1' )then
          cVar2S14S15P052P050nsss(0) <='1';
          else
          cVar2S14S15P052P050nsss(0) <='0';
          end if;
        if(cVar1S15S15N044P048N025P027(0)='1' AND  D( 4)='0' AND E( 5)='0' AND A(10)='0' )then
          cVar2S15S15P052N050P018nsss(0) <='1';
          else
          cVar2S15S15P052N050P018nsss(0) <='0';
          end if;
        if(cVar1S16S15N044P048N025N027(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S16S15P006P024nsss(0) <='1';
          else
          cVar2S16S15P006P024nsss(0) <='0';
          end if;
        if(cVar1S17S15N044P048N025N027(0)='1' AND  A(16)='1' AND B(17)='0' AND A(11)='0' )then
          cVar2S17S15P006N024P016nsss(0) <='1';
          else
          cVar2S17S15P006N024P016nsss(0) <='0';
          end if;
        if(cVar1S18S15N044P048N025N027(0)='1' AND  A(16)='0' AND D( 9)='0' AND A(15)='1' )then
          cVar2S18S15N006P065P008nsss(0) <='1';
          else
          cVar2S18S15N006P065P008nsss(0) <='0';
          end if;
        if(cVar1S19S15N044N048P007P040(0)='1' AND  A(18)='1' )then
          cVar2S19S15P002nsss(0) <='1';
          else
          cVar2S19S15P002nsss(0) <='0';
          end if;
        if(cVar1S20S15N044N048P007P040(0)='1' AND  A(18)='0' AND A(17)='1' )then
          cVar2S20S15N002P004nsss(0) <='1';
          else
          cVar2S20S15N002P004nsss(0) <='0';
          end if;
        if(cVar1S21S15N044N048P007P040(0)='1' AND  A(18)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S21S15N002N004P005nsss(0) <='1';
          else
          cVar2S21S15N002N004P005nsss(0) <='0';
          end if;
        if(cVar1S22S15N044N048P007N040(0)='1' AND  E( 7)='0' AND D( 8)='1' AND B( 2)='0' )then
          cVar2S22S15P042P069P035nsss(0) <='1';
          else
          cVar2S22S15P042P069P035nsss(0) <='0';
          end if;
        if(cVar1S23S15N044N048P007N040(0)='1' AND  E( 7)='1' AND D( 1)='1' )then
          cVar2S23S15P042P064nsss(0) <='1';
          else
          cVar2S23S15P042P064nsss(0) <='0';
          end if;
        if(cVar1S24S15N044N048P007N040(0)='1' AND  E( 7)='1' AND D( 1)='0' AND A( 7)='1' )then
          cVar2S24S15P042N064P005nsss(0) <='1';
          else
          cVar2S24S15P042N064P005nsss(0) <='0';
          end if;
        if(cVar1S25S15N044N048P007P043(0)='1' AND  B(18)='1' )then
          cVar2S25S15P022nsss(0) <='1';
          else
          cVar2S25S15P022nsss(0) <='0';
          end if;
        if(cVar1S26S15N044N048P007P043(0)='1' AND  B(18)='0' AND B( 8)='1' )then
          cVar2S26S15N022P023nsss(0) <='1';
          else
          cVar2S26S15N022P023nsss(0) <='0';
          end if;
        if(cVar1S27S15N044N048P007P043(0)='1' AND  B(18)='0' AND B( 8)='0' AND B( 7)='1' )then
          cVar2S27S15N022N023P025nsss(0) <='1';
          else
          cVar2S27S15N022N023P025nsss(0) <='0';
          end if;
        if(cVar1S28S15N044N048P007N043(0)='1' AND  D(13)='1' AND B( 7)='1' )then
          cVar2S28S15P049P025nsss(0) <='1';
          else
          cVar2S28S15P049P025nsss(0) <='0';
          end if;
        if(cVar1S29S15N044N048P007N043(0)='1' AND  D(13)='1' AND B( 7)='0' AND B(17)='1' )then
          cVar2S29S15P049N025P024nsss(0) <='1';
          else
          cVar2S29S15P049N025P024nsss(0) <='0';
          end if;
        if(cVar1S2S16P067P048N025N027(0)='1' AND  B(17)='1' AND A(16)='1' )then
          cVar2S2S16P024P006nsss(0) <='1';
          else
          cVar2S2S16P024P006nsss(0) <='0';
          end if;
        if(cVar1S3S16P067P048N025N027(0)='1' AND  B(17)='1' AND A(16)='0' AND E( 6)='1' )then
          cVar2S3S16P024N006P046nsss(0) <='1';
          else
          cVar2S3S16P024N006P046nsss(0) <='0';
          end if;
        if(cVar1S4S16P067P048N025N027(0)='1' AND  B(17)='0' AND A( 6)='0' )then
          cVar2S4S16N024P007nsss(0) <='1';
          else
          cVar2S4S16N024P007nsss(0) <='0';
          end if;
        if(cVar1S5S16P067N048P051P008(0)='1' AND  A( 3)='0' AND B(15)='1' )then
          cVar2S5S16P013P028nsss(0) <='1';
          else
          cVar2S5S16P013P028nsss(0) <='0';
          end if;
        if(cVar1S6S16P067N048P051P008(0)='1' AND  A( 3)='0' AND B(15)='0' AND B(16)='1' )then
          cVar2S6S16P013N028P026nsss(0) <='1';
          else
          cVar2S6S16P013N028P026nsss(0) <='0';
          end if;
        if(cVar1S7S16P067N048P051P008(0)='1' AND  A( 3)='1' )then
          cVar2S7S16P013psss(0) <='1';
          else
          cVar2S7S16P013psss(0) <='0';
          end if;
        if(cVar1S8S16P067N048P051N008(0)='1' AND  B(11)='0' )then
          cVar2S8S16P036nsss(0) <='1';
          else
          cVar2S8S16P036nsss(0) <='0';
          end if;
        if(cVar1S9S16P067N048P051N008(0)='1' AND  B(11)='1' AND A( 2)='1' )then
          cVar2S9S16P036P015nsss(0) <='1';
          else
          cVar2S9S16P036P015nsss(0) <='0';
          end if;
        if(cVar1S10S16P067N048N051P022(0)='1' AND  D(14)='1' )then
          cVar2S10S16P045nsss(0) <='1';
          else
          cVar2S10S16P045nsss(0) <='0';
          end if;
        if(cVar1S11S16P067N048N051P022(0)='1' AND  D(14)='0' AND D(15)='1' )then
          cVar2S11S16N045P041nsss(0) <='1';
          else
          cVar2S11S16N045P041nsss(0) <='0';
          end if;
        if(cVar1S12S16P067N048N051P022(0)='1' AND  D(14)='0' AND D(15)='0' AND D( 6)='1' )then
          cVar2S12S16N045N041P044nsss(0) <='1';
          else
          cVar2S12S16N045N041P044nsss(0) <='0';
          end if;
        if(cVar1S13S16P067N048N051N022(0)='1' AND  B(10)='1' AND D( 7)='1' )then
          cVar2S13S16P038P040nsss(0) <='1';
          else
          cVar2S13S16P038P040nsss(0) <='0';
          end if;
        if(cVar1S14S16P067N048N051N022(0)='1' AND  B(10)='1' AND D( 7)='0' AND A(13)='1' )then
          cVar2S14S16P038N040P012nsss(0) <='1';
          else
          cVar2S14S16P038N040P012nsss(0) <='0';
          end if;
        if(cVar1S15S16P067N048N051N022(0)='1' AND  B(10)='0' AND E(15)='0' )then
          cVar2S15S16N038P043nsss(0) <='1';
          else
          cVar2S15S16N038P043nsss(0) <='0';
          end if;
        if(cVar1S16S16P067N048N051N022(0)='1' AND  B(10)='0' AND E(15)='1' AND D(14)='1' )then
          cVar2S16S16N038P043P045nsss(0) <='1';
          else
          cVar2S16S16N038P043P045nsss(0) <='0';
          end if;
        if(cVar1S17S16P067P069P018P010(0)='1' AND  B( 3)='0' AND A(11)='0' AND B(12)='0' )then
          cVar2S17S16P033P016P034nsss(0) <='1';
          else
          cVar2S17S16P033P016P034nsss(0) <='0';
          end if;
        if(cVar1S18S16P067P069P018P010(0)='1' AND  B( 3)='0' AND A(11)='1' AND B(11)='1' )then
          cVar2S18S16P033P016P036nsss(0) <='1';
          else
          cVar2S18S16P033P016P036nsss(0) <='0';
          end if;
        if(cVar1S19S16P067P069P018P010(0)='1' AND  B( 3)='1' AND D(10)='1' )then
          cVar2S19S16P033P061nsss(0) <='1';
          else
          cVar2S19S16P033P061nsss(0) <='0';
          end if;
        if(cVar1S20S16P067P069P018P010(0)='1' AND  A(12)='1' AND A( 2)='0' )then
          cVar2S20S16P014P015nsss(0) <='1';
          else
          cVar2S20S16P014P015nsss(0) <='0';
          end if;
        if(cVar1S21S16P067P069N018P019(0)='1' AND  A( 3)='0' AND D( 9)='1' )then
          cVar2S21S16P013P065nsss(0) <='1';
          else
          cVar2S21S16P013P065nsss(0) <='0';
          end if;
        if(cVar1S22S16P067P069N018P019(0)='1' AND  A( 3)='0' AND D( 9)='0' AND B(12)='0' )then
          cVar2S22S16P013N065P034nsss(0) <='1';
          else
          cVar2S22S16P013N065P034nsss(0) <='0';
          end if;
        if(cVar1S23S16P067P069N018P019(0)='1' AND  A( 3)='1' AND A( 2)='1' )then
          cVar2S23S16P013P015nsss(0) <='1';
          else
          cVar2S23S16P013P015nsss(0) <='0';
          end if;
        if(cVar1S24S16P067P069N018N019(0)='1' AND  A(11)='1' AND B(11)='1' AND A(12)='0' )then
          cVar2S24S16P016P036P014nsss(0) <='1';
          else
          cVar2S24S16P016P036P014nsss(0) <='0';
          end if;
        if(cVar1S25S16P067P069N018N019(0)='1' AND  A(11)='1' AND B(11)='0' AND D( 0)='1' )then
          cVar2S25S16P016N036P068nsss(0) <='1';
          else
          cVar2S25S16P016N036P068nsss(0) <='0';
          end if;
        if(cVar1S26S16P067P069N018N019(0)='1' AND  A(11)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar2S26S16N016P017P015nsss(0) <='1';
          else
          cVar2S26S16N016P017P015nsss(0) <='0';
          end if;
        if(cVar1S28S16P067N069N052P065(0)='1' AND  E(10)='0' AND A( 2)='0' )then
          cVar2S28S16P063P015nsss(0) <='1';
          else
          cVar2S28S16P063P015nsss(0) <='0';
          end if;
        if(cVar1S29S16P067N069N052P065(0)='1' AND  E(10)='1' AND B(12)='1' )then
          cVar2S29S16P063P034nsss(0) <='1';
          else
          cVar2S29S16P063P034nsss(0) <='0';
          end if;
        if(cVar1S30S16P067N069N052N065(0)='1' AND  E(12)='1' )then
          cVar2S30S16P055nsss(0) <='1';
          else
          cVar2S30S16P055nsss(0) <='0';
          end if;
        if(cVar1S2S17P022N043P069N004(0)='1' AND  E( 1)='0' AND B(19)='1' )then
          cVar2S2S17P066P020nsss(0) <='1';
          else
          cVar2S2S17P066P020nsss(0) <='0';
          end if;
        if(cVar1S3S17P022N043P069N004(0)='1' AND  E( 1)='0' AND B(19)='0' AND B(17)='0' )then
          cVar2S3S17P066N020P024nsss(0) <='1';
          else
          cVar2S3S17P066N020P024nsss(0) <='0';
          end if;
        if(cVar1S5S17N022P048P025N007(0)='1' AND  A(16)='1' )then
          cVar2S5S17P006nsss(0) <='1';
          else
          cVar2S5S17P006nsss(0) <='0';
          end if;
        if(cVar1S6S17N022P048P025N007(0)='1' AND  A(16)='0' AND A( 5)='1' )then
          cVar2S6S17N006P009nsss(0) <='1';
          else
          cVar2S6S17N006P009nsss(0) <='0';
          end if;
        if(cVar1S7S17N022P048P025N007(0)='1' AND  A(16)='0' AND A( 5)='0' AND A( 7)='1' )then
          cVar2S7S17N006N009P005nsss(0) <='1';
          else
          cVar2S7S17N006N009P005nsss(0) <='0';
          end if;
        if(cVar1S8S17N022P048N025P027(0)='1' AND  A( 3)='0' )then
          cVar2S8S17P013nsss(0) <='1';
          else
          cVar2S8S17P013nsss(0) <='0';
          end if;
        if(cVar1S9S17N022P048N025N027(0)='1' AND  B(17)='1' AND A(13)='0' )then
          cVar2S9S17P024P012nsss(0) <='1';
          else
          cVar2S9S17P024P012nsss(0) <='0';
          end if;
        if(cVar1S10S17N022P048N025N027(0)='1' AND  B(17)='0' AND E( 5)='1' AND B(16)='1' )then
          cVar2S10S17N024P050P026nsss(0) <='1';
          else
          cVar2S10S17N024P050P026nsss(0) <='0';
          end if;
        if(cVar1S11S17N022P048N025N027(0)='1' AND  B(17)='0' AND E( 5)='0' AND A(12)='1' )then
          cVar2S11S17N024N050P014nsss(0) <='1';
          else
          cVar2S11S17N024N050P014nsss(0) <='0';
          end if;
        if(cVar1S12S17N022N048P051P008(0)='1' AND  A( 3)='0' AND B(15)='1' )then
          cVar2S12S17P013P028nsss(0) <='1';
          else
          cVar2S12S17P013P028nsss(0) <='0';
          end if;
        if(cVar1S13S17N022N048P051P008(0)='1' AND  A( 3)='0' AND B(15)='0' AND B(16)='1' )then
          cVar2S13S17P013N028P026nsss(0) <='1';
          else
          cVar2S13S17P013N028P026nsss(0) <='0';
          end if;
        if(cVar1S14S17N022N048P051P008(0)='1' AND  A( 3)='1' AND B(16)='1' )then
          cVar2S14S17P013P026nsss(0) <='1';
          else
          cVar2S14S17P013P026nsss(0) <='0';
          end if;
        if(cVar1S15S17N022N048P051N008(0)='1' AND  A(14)='1' AND B(11)='0' )then
          cVar2S15S17P010P036nsss(0) <='1';
          else
          cVar2S15S17P010P036nsss(0) <='0';
          end if;
        if(cVar1S16S17N022N048P051N008(0)='1' AND  A(14)='0' AND A( 4)='1' )then
          cVar2S16S17N010P011nsss(0) <='1';
          else
          cVar2S16S17N010P011nsss(0) <='0';
          end if;
        if(cVar1S17S17N022N048P051N008(0)='1' AND  A(14)='0' AND A( 4)='0' AND A( 5)='1' )then
          cVar2S17S17N010N011P009nsss(0) <='1';
          else
          cVar2S17S17N010N011P009nsss(0) <='0';
          end if;
        if(cVar1S18S17N022N048N051P038(0)='1' AND  B( 9)='1' AND A( 2)='0' )then
          cVar2S18S17P021P015nsss(0) <='1';
          else
          cVar2S18S17P021P015nsss(0) <='0';
          end if;
        if(cVar1S19S17N022N048N051P038(0)='1' AND  B( 9)='0' AND A(19)='1' )then
          cVar2S19S17N021P000nsss(0) <='1';
          else
          cVar2S19S17N021P000nsss(0) <='0';
          end if;
        if(cVar1S20S17N022N048N051P038(0)='1' AND  B( 9)='0' AND A(19)='0' AND A(17)='1' )then
          cVar2S20S17N021N000P004nsss(0) <='1';
          else
          cVar2S20S17N021N000P004nsss(0) <='0';
          end if;
        if(cVar1S21S17N022N048N051N038(0)='1' AND  D( 4)='1' AND A( 5)='1' AND E( 1)='0' )then
          cVar2S21S17P052P009P066nsss(0) <='1';
          else
          cVar2S21S17P052P009P066nsss(0) <='0';
          end if;
        if(cVar1S22S17N022N048N051N038(0)='1' AND  D( 4)='1' AND A( 5)='0' AND A(14)='1' )then
          cVar2S22S17P052N009P010nsss(0) <='1';
          else
          cVar2S22S17P052N009P010nsss(0) <='0';
          end if;
        if(cVar1S23S17N022N048N051N038(0)='1' AND  D( 4)='0' AND A( 5)='0' AND D(10)='1' )then
          cVar2S23S17N052P009P061nsss(0) <='1';
          else
          cVar2S23S17N052P009P061nsss(0) <='0';
          end if;
        if(cVar1S24S17N022N048N051N038(0)='1' AND  D( 4)='0' AND A( 5)='1' AND E(14)='1' )then
          cVar2S24S17N052P009P047nsss(0) <='1';
          else
          cVar2S24S17N052P009P047nsss(0) <='0';
          end if;
        if(cVar1S2S18P041N020N021P022(0)='1' AND  A(17)='1' )then
          cVar2S2S18P004nsss(0) <='1';
          else
          cVar2S2S18P004nsss(0) <='0';
          end if;
        if(cVar1S3S18P041N020N021P022(0)='1' AND  A(17)='0' AND A( 7)='1' )then
          cVar2S3S18N004P005nsss(0) <='1';
          else
          cVar2S3S18N004P005nsss(0) <='0';
          end if;
        if(cVar1S4S18P041N020N021N022(0)='1' AND  B( 8)='1' )then
          cVar2S4S18P023nsss(0) <='1';
          else
          cVar2S4S18P023nsss(0) <='0';
          end if;
        if(cVar1S5S18P041N020N021N022(0)='1' AND  B( 8)='0' AND D(10)='1' )then
          cVar2S5S18N023P061nsss(0) <='1';
          else
          cVar2S5S18N023P061nsss(0) <='0';
          end if;
        if(cVar1S6S18N041P039P020P044(0)='1' AND  B( 8)='1' )then
          cVar2S6S18P023nsss(0) <='1';
          else
          cVar2S6S18P023nsss(0) <='0';
          end if;
        if(cVar1S7S18N041P039P020P044(0)='1' AND  B( 8)='0' AND A(17)='1' )then
          cVar2S7S18N023P004nsss(0) <='1';
          else
          cVar2S7S18N023P004nsss(0) <='0';
          end if;
        if(cVar1S8S18N041P039P020P044(0)='1' AND  B( 8)='0' AND A(17)='0' AND B( 7)='1' )then
          cVar2S8S18N023N004P025nsss(0) <='1';
          else
          cVar2S8S18N023N004P025nsss(0) <='0';
          end if;
        if(cVar1S9S18N041P039P020N044(0)='1' AND  E( 7)='0' AND E( 5)='1' )then
          cVar2S9S18P042P050nsss(0) <='1';
          else
          cVar2S9S18P042P050nsss(0) <='0';
          end if;
        if(cVar1S10S18N041P039P020N044(0)='1' AND  E( 7)='0' AND E( 5)='0' AND A(18)='0' )then
          cVar2S10S18P042N050P002nsss(0) <='1';
          else
          cVar2S10S18P042N050P002nsss(0) <='0';
          end if;
        if(cVar1S11S18N041P039P020N044(0)='1' AND  E( 7)='1' AND D( 7)='1' )then
          cVar2S11S18P042P040nsss(0) <='1';
          else
          cVar2S11S18P042P040nsss(0) <='0';
          end if;
        if(cVar1S12S18N041P039P020N044(0)='1' AND  E( 7)='1' AND D( 7)='0' AND D( 1)='1' )then
          cVar2S12S18P042N040P064nsss(0) <='1';
          else
          cVar2S12S18P042N040P064nsss(0) <='0';
          end if;
        if(cVar1S13S18N041P039P020P040(0)='1' AND  A(18)='1' )then
          cVar2S13S18P002nsss(0) <='1';
          else
          cVar2S13S18P002nsss(0) <='0';
          end if;
        if(cVar1S14S18N041P039P020N040(0)='1' AND  B(17)='1' )then
          cVar2S14S18P024nsss(0) <='1';
          else
          cVar2S14S18P024nsss(0) <='0';
          end if;
        if(cVar1S15S18N041P039P020N040(0)='1' AND  B(17)='0' AND B( 1)='1' AND A(13)='0' )then
          cVar2S15S18N024P037P012nsss(0) <='1';
          else
          cVar2S15S18N024P037P012nsss(0) <='0';
          end if;
        if(cVar1S18S18N041P039N005N020(0)='1' AND  E(13)='1' )then
          cVar2S18S18P051nsss(0) <='1';
          else
          cVar2S18S18P051nsss(0) <='0';
          end if;
        if(cVar1S2S19P041N020P021N003(0)='1' AND  D( 7)='0' )then
          cVar2S2S19P040nsss(0) <='1';
          else
          cVar2S2S19P040nsss(0) <='0';
          end if;
        if(cVar1S3S19P041N020N021P022(0)='1' AND  A(17)='1' )then
          cVar2S3S19P004nsss(0) <='1';
          else
          cVar2S3S19P004nsss(0) <='0';
          end if;
        if(cVar1S4S19P041N020N021P022(0)='1' AND  A(17)='0' AND A( 7)='1' )then
          cVar2S4S19N004P005nsss(0) <='1';
          else
          cVar2S4S19N004P005nsss(0) <='0';
          end if;
        if(cVar1S5S19P041N020N021N022(0)='1' AND  B( 8)='1' )then
          cVar2S5S19P023nsss(0) <='1';
          else
          cVar2S5S19P023nsss(0) <='0';
          end if;
        if(cVar1S6S19P041N020N021N022(0)='1' AND  B( 8)='0' AND E(14)='1' )then
          cVar2S6S19N023P047nsss(0) <='1';
          else
          cVar2S6S19N023P047nsss(0) <='0';
          end if;
        if(cVar1S7S19P041N020N021N022(0)='1' AND  B( 8)='0' AND E(14)='0' AND D(10)='1' )then
          cVar2S7S19N023N047P061nsss(0) <='1';
          else
          cVar2S7S19N023N047P061nsss(0) <='0';
          end if;
        if(cVar1S8S19N041P039P044P023(0)='1' AND  A( 7)='1' )then
          cVar2S8S19P005nsss(0) <='1';
          else
          cVar2S8S19P005nsss(0) <='0';
          end if;
        if(cVar1S9S19N041P039P044P023(0)='1' AND  A( 7)='0' AND A(17)='1' )then
          cVar2S9S19N005P004nsss(0) <='1';
          else
          cVar2S9S19N005P004nsss(0) <='0';
          end if;
        if(cVar1S10S19N041P039P044P023(0)='1' AND  A( 7)='0' AND A(17)='0' AND A( 2)='0' )then
          cVar2S10S19N005N004P015nsss(0) <='1';
          else
          cVar2S10S19N005N004P015nsss(0) <='0';
          end if;
        if(cVar1S12S19N041P039N044P050(0)='1' AND  A( 5)='1' AND B( 6)='1' )then
          cVar2S12S19P009P027nsss(0) <='1';
          else
          cVar2S12S19P009P027nsss(0) <='0';
          end if;
        if(cVar1S13S19N041P039N044P050(0)='1' AND  A( 5)='1' AND B( 6)='0' AND B( 5)='1' )then
          cVar2S13S19P009N027P029nsss(0) <='1';
          else
          cVar2S13S19P009N027P029nsss(0) <='0';
          end if;
        if(cVar1S14S19N041P039N044P050(0)='1' AND  A( 5)='0' AND A(15)='1' AND A( 4)='0' )then
          cVar2S14S19N009P008P011nsss(0) <='1';
          else
          cVar2S14S19N009P008P011nsss(0) <='0';
          end if;
        if(cVar1S15S19N041P039N044P050(0)='1' AND  A( 5)='0' AND A(15)='0' AND A( 4)='1' )then
          cVar2S15S19N009N008P011nsss(0) <='1';
          else
          cVar2S15S19N009N008P011nsss(0) <='0';
          end if;
        if(cVar1S16S19N041P039N044N050(0)='1' AND  A(19)='0' AND A( 2)='1' AND B( 3)='1' )then
          cVar2S16S19P000P015P033nsss(0) <='1';
          else
          cVar2S16S19P000P015P033nsss(0) <='0';
          end if;
        if(cVar1S17S19N041P039N044N050(0)='1' AND  A(19)='0' AND A( 2)='0' AND E( 4)='1' )then
          cVar2S17S19P000N015P054nsss(0) <='1';
          else
          cVar2S17S19P000N015P054nsss(0) <='0';
          end if;
        if(cVar1S18S19N041P039N044N050(0)='1' AND  A(19)='1' AND D( 7)='1' )then
          cVar2S18S19P000P040nsss(0) <='1';
          else
          cVar2S18S19P000P040nsss(0) <='0';
          end if;
        if(cVar1S20S19N041P039N005N064(0)='1' AND  B(19)='1' )then
          cVar2S20S19P020nsss(0) <='1';
          else
          cVar2S20S19P020nsss(0) <='0';
          end if;
        if(cVar1S0S20P011P029P048P025(0)='1' AND  A( 6)='1' )then
          cVar2S0S20P007nsss(0) <='1';
          else
          cVar2S0S20P007nsss(0) <='0';
          end if;
        if(cVar1S1S20P011P029P048P025(0)='1' AND  A( 6)='0' AND A(17)='1' )then
          cVar2S1S20N007P004nsss(0) <='1';
          else
          cVar2S1S20N007P004nsss(0) <='0';
          end if;
        if(cVar1S2S20P011P029P048P025(0)='1' AND  A( 6)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S2S20N007N004P006nsss(0) <='1';
          else
          cVar2S2S20N007N004P006nsss(0) <='0';
          end if;
        if(cVar1S4S20P011P029N048P041(0)='1' AND  B(19)='1' )then
          cVar2S4S20P020nsss(0) <='1';
          else
          cVar2S4S20P020nsss(0) <='0';
          end if;
        if(cVar1S5S20P011P029N048P041(0)='1' AND  B(19)='0' AND B( 9)='1' )then
          cVar2S5S20N020P021nsss(0) <='1';
          else
          cVar2S5S20N020P021nsss(0) <='0';
          end if;
        if(cVar1S6S20P011P029N048P041(0)='1' AND  B(19)='0' AND B( 9)='0' AND B(18)='1' )then
          cVar2S6S20N020N021P022nsss(0) <='1';
          else
          cVar2S6S20N020N021P022nsss(0) <='0';
          end if;
        if(cVar1S7S20P011P029N048N041(0)='1' AND  B( 0)='0' AND A( 6)='0' )then
          cVar2S7S20P039P007nsss(0) <='1';
          else
          cVar2S7S20P039P007nsss(0) <='0';
          end if;
        if(cVar1S8S20P011P029N048N041(0)='1' AND  B( 0)='0' AND A( 6)='1' AND B( 7)='1' )then
          cVar2S8S20P039P007P025nsss(0) <='1';
          else
          cVar2S8S20P039P007P025nsss(0) <='0';
          end if;
        if(cVar1S9S20P011P029N048N041(0)='1' AND  B( 0)='1' AND D( 1)='1' )then
          cVar2S9S20P039P064nsss(0) <='1';
          else
          cVar2S9S20P039P064nsss(0) <='0';
          end if;
        if(cVar1S10S20P011P029N048N041(0)='1' AND  B( 0)='1' AND D( 1)='0' AND A( 7)='1' )then
          cVar2S10S20P039N064P005nsss(0) <='1';
          else
          cVar2S10S20P039N064P005nsss(0) <='0';
          end if;
        if(cVar1S12S20P011P029P010N052(0)='1' AND  E( 4)='1' )then
          cVar2S12S20P054nsss(0) <='1';
          else
          cVar2S12S20P054nsss(0) <='0';
          end if;
        if(cVar1S13S20P011P029N010P009(0)='1' AND  E( 5)='1' )then
          cVar2S13S20P050nsss(0) <='1';
          else
          cVar2S13S20P050nsss(0) <='0';
          end if;
        if(cVar1S14S20P011P029N010P009(0)='1' AND  E( 5)='0' AND D(12)='1' )then
          cVar2S14S20N050P053nsss(0) <='1';
          else
          cVar2S14S20N050P053nsss(0) <='0';
          end if;
        if(cVar1S15S20P011P029N010N009(0)='1' AND  A(15)='1' AND D( 4)='1' )then
          cVar2S15S20P008P052nsss(0) <='1';
          else
          cVar2S15S20P008P052nsss(0) <='0';
          end if;
        if(cVar1S16S20P011P029P060P014(0)='1' AND  A(11)='0' AND B( 3)='0' )then
          cVar2S16S20P016P033nsss(0) <='1';
          else
          cVar2S16S20P016P033nsss(0) <='0';
          end if;
        if(cVar1S17S20P011P029P060P014(0)='1' AND  A(11)='1' AND A(10)='0' )then
          cVar2S17S20P016P018nsss(0) <='1';
          else
          cVar2S17S20P016P018nsss(0) <='0';
          end if;
        if(cVar1S18S20P011P029P060P014(0)='1' AND  D(12)='1' )then
          cVar2S18S20P053nsss(0) <='1';
          else
          cVar2S18S20P053nsss(0) <='0';
          end if;
        if(cVar1S19S20P011P029P060P014(0)='1' AND  D(12)='0' AND A(10)='0' )then
          cVar2S19S20N053P018nsss(0) <='1';
          else
          cVar2S19S20N053P018nsss(0) <='0';
          end if;
        if(cVar1S20S20P011N029P015P033(0)='1' AND  A( 8)='1' AND A( 5)='0' )then
          cVar2S20S20P003P009nsss(0) <='1';
          else
          cVar2S20S20P003P009nsss(0) <='0';
          end if;
        if(cVar1S21S20P011N029P015P033(0)='1' AND  A( 8)='0' AND E(12)='1' )then
          cVar2S21S20N003P055nsss(0) <='1';
          else
          cVar2S21S20N003P055nsss(0) <='0';
          end if;
        if(cVar1S22S20P011N029P015P033(0)='1' AND  A( 8)='0' AND E(12)='0' AND E(15)='0' )then
          cVar2S22S20N003N055P043nsss(0) <='1';
          else
          cVar2S22S20N003N055P043nsss(0) <='0';
          end if;
        if(cVar1S23S20P011N029P015P033(0)='1' AND  D( 8)='0' AND A( 3)='1' )then
          cVar2S23S20P069P013nsss(0) <='1';
          else
          cVar2S23S20P069P013nsss(0) <='0';
          end if;
        if(cVar1S24S20P011N029N015P017(0)='1' AND  B( 2)='0' AND A(12)='1' AND A(15)='0' )then
          cVar2S24S20P035P014P008nsss(0) <='1';
          else
          cVar2S24S20P035P014P008nsss(0) <='0';
          end if;
        if(cVar1S25S20P011N029N015P017(0)='1' AND  B( 2)='0' AND A(12)='0' AND B( 4)='1' )then
          cVar2S25S20P035N014P031nsss(0) <='1';
          else
          cVar2S25S20P035N014P031nsss(0) <='0';
          end if;
        if(cVar1S26S20P011N029N015P017(0)='1' AND  B( 2)='1' AND A(13)='0' AND E( 2)='1' )then
          cVar2S26S20P035P012P062nsss(0) <='1';
          else
          cVar2S26S20P035P012P062nsss(0) <='0';
          end if;
        if(cVar1S27S20P011N029N015N017(0)='1' AND  E( 4)='1' AND B( 4)='1' )then
          cVar2S27S20P054P031nsss(0) <='1';
          else
          cVar2S27S20P054P031nsss(0) <='0';
          end if;
        if(cVar1S28S20P011N029N015N017(0)='1' AND  E( 4)='0' AND D( 1)='0' AND D(13)='1' )then
          cVar2S28S20N054P064P049nsss(0) <='1';
          else
          cVar2S28S20N054P064P049nsss(0) <='0';
          end if;
        if(cVar1S2S21P041N020P021N003(0)='1' AND  D( 7)='0' )then
          cVar2S2S21P040nsss(0) <='1';
          else
          cVar2S2S21P040nsss(0) <='0';
          end if;
        if(cVar1S4S21P041N020N021N004(0)='1' AND  B( 8)='1' )then
          cVar2S4S21P023nsss(0) <='1';
          else
          cVar2S4S21P023nsss(0) <='0';
          end if;
        if(cVar1S5S21P041N020N021N004(0)='1' AND  B( 8)='0' AND B(18)='1' AND A( 7)='1' )then
          cVar2S5S21N023P022P005nsss(0) <='1';
          else
          cVar2S5S21N023P022P005nsss(0) <='0';
          end if;
        if(cVar1S6S21P041N020N021N004(0)='1' AND  B( 8)='0' AND B(18)='0' AND D(10)='1' )then
          cVar2S6S21N023N022P061nsss(0) <='1';
          else
          cVar2S6S21N023N022P061nsss(0) <='0';
          end if;
        if(cVar1S7S21N041P039P000P048(0)='1' AND  B( 7)='1' )then
          cVar2S7S21P025nsss(0) <='1';
          else
          cVar2S7S21P025nsss(0) <='0';
          end if;
        if(cVar1S8S21N041P039P000P048(0)='1' AND  B( 7)='0' AND B( 6)='1' )then
          cVar2S8S21N025P027nsss(0) <='1';
          else
          cVar2S8S21N025P027nsss(0) <='0';
          end if;
        if(cVar1S9S21N041P039P000P048(0)='1' AND  B( 7)='0' AND B( 6)='0' AND D(13)='1' )then
          cVar2S9S21N025N027P049nsss(0) <='1';
          else
          cVar2S9S21N025N027P049nsss(0) <='0';
          end if;
        if(cVar1S10S21N041P039P000N048(0)='1' AND  E(13)='1' AND A(15)='1' AND A( 3)='0' )then
          cVar2S10S21P051P008P013nsss(0) <='1';
          else
          cVar2S10S21P051P008P013nsss(0) <='0';
          end if;
        if(cVar1S11S21N041P039P000N048(0)='1' AND  E(13)='1' AND A(15)='0' AND A( 0)='0' )then
          cVar2S11S21P051N008P019nsss(0) <='1';
          else
          cVar2S11S21P051N008P019nsss(0) <='0';
          end if;
        if(cVar1S12S21N041P039P000N048(0)='1' AND  E(13)='0' AND E(12)='1' AND B(14)='1' )then
          cVar2S12S21N051P055P030nsss(0) <='1';
          else
          cVar2S12S21N051P055P030nsss(0) <='0';
          end if;
        if(cVar1S14S21N041P039P000N040(0)='1' AND  A( 2)='1' AND A(12)='0' AND E( 2)='0' )then
          cVar2S14S21P015P014P062nsss(0) <='1';
          else
          cVar2S14S21P015P014P062nsss(0) <='0';
          end if;
        if(cVar1S15S21N041P039P000N040(0)='1' AND  A( 2)='0' AND A( 1)='1' AND A(15)='1' )then
          cVar2S15S21N015P017P008nsss(0) <='1';
          else
          cVar2S15S21N015P017P008nsss(0) <='0';
          end if;
        if(cVar1S1S22P000P041N020P005(0)='1' AND  B( 9)='1' )then
          cVar2S1S22P021nsss(0) <='1';
          else
          cVar2S1S22P021nsss(0) <='0';
          end if;
        if(cVar1S2S22P000P041N020P005(0)='1' AND  B( 9)='0' AND A( 1)='0' )then
          cVar2S2S22N021P017nsss(0) <='1';
          else
          cVar2S2S22N021P017nsss(0) <='0';
          end if;
        if(cVar1S3S22P000P041N020N005(0)='1' AND  A( 8)='1' AND B( 9)='1' )then
          cVar2S3S22P003P021nsss(0) <='1';
          else
          cVar2S3S22P003P021nsss(0) <='0';
          end if;
        if(cVar1S4S22P000P041N020N005(0)='1' AND  A( 8)='0' AND B(18)='1' )then
          cVar2S4S22N003P022nsss(0) <='1';
          else
          cVar2S4S22N003P022nsss(0) <='0';
          end if;
        if(cVar1S5S22P000P041N020N005(0)='1' AND  A( 8)='0' AND B(18)='0' AND A(17)='1' )then
          cVar2S5S22N003N022P004nsss(0) <='1';
          else
          cVar2S5S22N003N022P004nsss(0) <='0';
          end if;
        if(cVar1S6S22P000N041P039P012(0)='1' AND  B(14)='0' AND D( 7)='1' )then
          cVar2S6S22P030P040nsss(0) <='1';
          else
          cVar2S6S22P030P040nsss(0) <='0';
          end if;
        if(cVar1S7S22P000N041P039P012(0)='1' AND  B(14)='0' AND D( 7)='0' AND D(11)='0' )then
          cVar2S7S22P030N040P057nsss(0) <='1';
          else
          cVar2S7S22P030N040P057nsss(0) <='0';
          end if;
        if(cVar1S8S22P000N041P039P012(0)='1' AND  B(14)='1' AND A(14)='1' AND A( 5)='0' )then
          cVar2S8S22P030P010P009nsss(0) <='1';
          else
          cVar2S8S22P030P010P009nsss(0) <='0';
          end if;
        if(cVar1S9S22P000N041P039P012(0)='1' AND  B(14)='1' AND B( 4)='0' AND B(11)='0' )then
          cVar2S9S22P030P031P036nsss(0) <='1';
          else
          cVar2S9S22P030P031P036nsss(0) <='0';
          end if;
        if(cVar1S10S22P000N041P039P012(0)='1' AND  B(14)='0' AND B(13)='1' AND A(14)='0' )then
          cVar2S10S22N030P032P010nsss(0) <='1';
          else
          cVar2S10S22N030P032P010nsss(0) <='0';
          end if;
        if(cVar1S11S22P000N041P039P012(0)='1' AND  B(14)='0' AND B(13)='0' AND A( 1)='1' )then
          cVar2S11S22N030N032P017nsss(0) <='1';
          else
          cVar2S11S22N030N032P017nsss(0) <='0';
          end if;
        if(cVar1S13S22P000N041P039N049(0)='1' AND  B(19)='1' )then
          cVar2S13S22P020nsss(0) <='1';
          else
          cVar2S13S22P020nsss(0) <='0';
          end if;
        if(cVar1S14S22P000N041P039N049(0)='1' AND  B(19)='0' AND D( 1)='1' )then
          cVar2S14S22N020P064nsss(0) <='1';
          else
          cVar2S14S22N020P064nsss(0) <='0';
          end if;
        if(cVar1S15S22P000N041P039N049(0)='1' AND  B(19)='0' AND D( 1)='0' AND A( 7)='1' )then
          cVar2S15S22N020N064P005nsss(0) <='1';
          else
          cVar2S15S22N020N064P005nsss(0) <='0';
          end if;
        if(cVar1S18S22P000N040P059N041(0)='1' AND  A(10)='1' AND A(13)='1' AND A(11)='1' )then
          cVar2S18S22P018P012P016nsss(0) <='1';
          else
          cVar2S18S22P018P012P016nsss(0) <='0';
          end if;
        if(cVar1S19S22P000N040P059N041(0)='1' AND  A(10)='0' AND D( 4)='1' )then
          cVar2S19S22N018P052nsss(0) <='1';
          else
          cVar2S19S22N018P052nsss(0) <='0';
          end if;
        if(cVar1S2S23P041N020P005N021(0)='1' AND  B(18)='1' )then
          cVar2S2S23P022nsss(0) <='1';
          else
          cVar2S2S23P022nsss(0) <='0';
          end if;
        if(cVar1S3S23P041N020P005N021(0)='1' AND  B(18)='0' AND E( 7)='1' )then
          cVar2S3S23N022P042nsss(0) <='1';
          else
          cVar2S3S23N022P042nsss(0) <='0';
          end if;
        if(cVar1S4S23P041N020N005P003(0)='1' AND  B( 9)='1' )then
          cVar2S4S23P021nsss(0) <='1';
          else
          cVar2S4S23P021nsss(0) <='0';
          end if;
        if(cVar1S5S23P041N020N005N003(0)='1' AND  A(17)='1' )then
          cVar2S5S23P004nsss(0) <='1';
          else
          cVar2S5S23P004nsss(0) <='0';
          end if;
        if(cVar1S6S23N041P055P061P056(0)='1' AND  A(14)='1' AND B(15)='1' )then
          cVar2S6S23P010P028nsss(0) <='1';
          else
          cVar2S6S23P010P028nsss(0) <='0';
          end if;
        if(cVar1S7S23N041P055P061P056(0)='1' AND  A(14)='1' AND B(15)='0' AND B(14)='1' )then
          cVar2S7S23P010N028P030nsss(0) <='1';
          else
          cVar2S7S23P010N028P030nsss(0) <='0';
          end if;
        if(cVar1S8S23N041P055P061P056(0)='1' AND  A(14)='0' AND E( 3)='0' )then
          cVar2S8S23N010P058nsss(0) <='1';
          else
          cVar2S8S23N010P058nsss(0) <='0';
          end if;
        if(cVar1S9S23N041P055P061P056(0)='1' AND  B( 5)='0' AND B( 3)='1' )then
          cVar2S9S23P029P033nsss(0) <='1';
          else
          cVar2S9S23P029P033nsss(0) <='0';
          end if;
        if(cVar1S11S23N041P055P061N054(0)='1' AND  B(14)='1' )then
          cVar2S11S23P030nsss(0) <='1';
          else
          cVar2S11S23P030nsss(0) <='0';
          end if;
        if(cVar1S12S23N041N055P010P039(0)='1' AND  A(15)='1' AND B(16)='1' )then
          cVar2S12S23P008P026nsss(0) <='1';
          else
          cVar2S12S23P008P026nsss(0) <='0';
          end if;
        if(cVar1S13S23N041N055P010P039(0)='1' AND  A(15)='1' AND B(16)='0' AND B( 6)='1' )then
          cVar2S13S23P008N026P027nsss(0) <='1';
          else
          cVar2S13S23P008N026P027nsss(0) <='0';
          end if;
        if(cVar1S14S23N041N055P010P039(0)='1' AND  A(15)='0' AND B(10)='1' )then
          cVar2S14S23N008P038nsss(0) <='1';
          else
          cVar2S14S23N008P038nsss(0) <='0';
          end if;
        if(cVar1S15S23N041N055P010P039(0)='1' AND  A(15)='0' AND B(10)='0' AND E( 3)='1' )then
          cVar2S15S23N008N038P058nsss(0) <='1';
          else
          cVar2S15S23N008N038P058nsss(0) <='0';
          end if;
        if(cVar1S16S23N041N055P010P039(0)='1' AND  A( 7)='1' )then
          cVar2S16S23P005nsss(0) <='1';
          else
          cVar2S16S23P005nsss(0) <='0';
          end if;
        if(cVar1S17S23N041N055P010P028(0)='1' AND  B( 2)='0' AND D( 8)='0' )then
          cVar2S17S23P035P069nsss(0) <='1';
          else
          cVar2S17S23P035P069nsss(0) <='0';
          end if;
        if(cVar1S18S23N041N055P010N028(0)='1' AND  B( 5)='1' AND E(10)='0' AND A(15)='0' )then
          cVar2S18S23P029P063P008nsss(0) <='1';
          else
          cVar2S18S23P029P063P008nsss(0) <='0';
          end if;
        if(cVar1S19S23N041N055P010N028(0)='1' AND  B( 5)='0' AND B(14)='1' AND A(12)='0' )then
          cVar2S19S23N029P030P014nsss(0) <='1';
          else
          cVar2S19S23N029P030P014nsss(0) <='0';
          end if;
        if(cVar1S2S24P041N020P005N021(0)='1' AND  B(18)='1' )then
          cVar2S2S24P022nsss(0) <='1';
          else
          cVar2S2S24P022nsss(0) <='0';
          end if;
        if(cVar1S3S24P041N020P005N021(0)='1' AND  B(18)='0' AND E( 7)='1' )then
          cVar2S3S24N022P042nsss(0) <='1';
          else
          cVar2S3S24N022P042nsss(0) <='0';
          end if;
        if(cVar1S4S24P041N020N005P003(0)='1' AND  B( 9)='1' )then
          cVar2S4S24P021nsss(0) <='1';
          else
          cVar2S4S24P021nsss(0) <='0';
          end if;
        if(cVar1S5S24P041N020N005N003(0)='1' AND  B(18)='1' AND A(17)='1' )then
          cVar2S5S24P022P004nsss(0) <='1';
          else
          cVar2S5S24P022P004nsss(0) <='0';
          end if;
        if(cVar1S6S24P041N020N005N003(0)='1' AND  B(18)='0' AND D(10)='1' )then
          cVar2S6S24N022P061nsss(0) <='1';
          else
          cVar2S6S24N022P061nsss(0) <='0';
          end if;
        if(cVar1S7S24N041P039P058P033(0)='1' AND  D( 2)='0' AND A( 3)='0' )then
          cVar2S7S24P060P013nsss(0) <='1';
          else
          cVar2S7S24P060P013nsss(0) <='0';
          end if;
        if(cVar1S8S24N041P039P058P033(0)='1' AND  D( 2)='0' AND A( 3)='1' AND B( 4)='1' )then
          cVar2S8S24P060P013P031nsss(0) <='1';
          else
          cVar2S8S24P060P013P031nsss(0) <='0';
          end if;
        if(cVar1S9S24N041P039P058P033(0)='1' AND  D( 2)='1' AND B( 2)='1' AND D( 1)='0' )then
          cVar2S9S24P060P035P064nsss(0) <='1';
          else
          cVar2S9S24P060P035P064nsss(0) <='0';
          end if;
        if(cVar1S10S24N041P039P058P033(0)='1' AND  D( 2)='1' AND B( 2)='0' AND E( 1)='1' )then
          cVar2S10S24P060N035P066nsss(0) <='1';
          else
          cVar2S10S24P060N035P066nsss(0) <='0';
          end if;
        if(cVar1S11S24N041P039P058P033(0)='1' AND  E(10)='0' AND A(12)='1' AND A(11)='0' )then
          cVar2S11S24P063P014P016nsss(0) <='1';
          else
          cVar2S11S24P063P014P016nsss(0) <='0';
          end if;
        if(cVar1S12S24N041P039P058P033(0)='1' AND  E(10)='0' AND A(12)='0' AND E( 2)='1' )then
          cVar2S12S24P063N014P062nsss(0) <='1';
          else
          cVar2S12S24P063N014P062nsss(0) <='0';
          end if;
        if(cVar1S13S24N041P039P058P033(0)='1' AND  E(10)='1' AND B(12)='1' AND A(11)='1' )then
          cVar2S13S24P063P034P016nsss(0) <='1';
          else
          cVar2S13S24P063P034P016nsss(0) <='0';
          end if;
        if(cVar1S14S24N041P039P058P033(0)='1' AND  A( 9)='0' AND A(14)='0' )then
          cVar2S14S24P001P010nsss(0) <='1';
          else
          cVar2S14S24P001P010nsss(0) <='0';
          end if;
        if(cVar1S15S24N041P039P058N033(0)='1' AND  D( 3)='1' AND A( 3)='1' )then
          cVar2S15S24P056P013nsss(0) <='1';
          else
          cVar2S15S24P056P013nsss(0) <='0';
          end if;
        if(cVar1S16S24N041P039P058N033(0)='1' AND  D( 3)='1' AND A( 3)='0' AND A(13)='1' )then
          cVar2S16S24P056N013P012nsss(0) <='1';
          else
          cVar2S16S24P056N013P012nsss(0) <='0';
          end if;
        if(cVar1S17S24N041P039P058N033(0)='1' AND  D( 3)='0' AND A(12)='1' AND B(13)='1' )then
          cVar2S17S24N056P014P032nsss(0) <='1';
          else
          cVar2S17S24N056P014P032nsss(0) <='0';
          end if;
        if(cVar1S20S24N041P039N051N064(0)='1' AND  A(14)='0' AND B(19)='1' )then
          cVar2S20S24P010P020nsss(0) <='1';
          else
          cVar2S20S24P010P020nsss(0) <='0';
          end if;
        if(cVar1S2S25P041N020P005N021(0)='1' AND  A( 1)='0' )then
          cVar2S2S25P017nsss(0) <='1';
          else
          cVar2S2S25P017nsss(0) <='0';
          end if;
        if(cVar1S3S25P041N020N005P003(0)='1' AND  B( 9)='1' )then
          cVar2S3S25P021nsss(0) <='1';
          else
          cVar2S3S25P021nsss(0) <='0';
          end if;
        if(cVar1S4S25P041N020N005N003(0)='1' AND  D( 9)='0' AND B(18)='1' )then
          cVar2S4S25P065P022nsss(0) <='1';
          else
          cVar2S4S25P065P022nsss(0) <='0';
          end if;
        if(cVar1S5S25P041N020N005N003(0)='1' AND  D( 9)='0' AND B(18)='0' AND A(10)='0' )then
          cVar2S5S25P065N022P018nsss(0) <='1';
          else
          cVar2S5S25P065N022P018nsss(0) <='0';
          end if;
        if(cVar1S6S25N041P013P031P056(0)='1' AND  A(11)='0' AND A(14)='0' )then
          cVar2S6S25P016P010nsss(0) <='1';
          else
          cVar2S6S25P016P010nsss(0) <='0';
          end if;
        if(cVar1S7S25N041P013P031P056(0)='1' AND  A(11)='1' AND A( 0)='0' )then
          cVar2S7S25P016P019nsss(0) <='1';
          else
          cVar2S7S25P016P019nsss(0) <='0';
          end if;
        if(cVar1S8S25N041P013P031N056(0)='1' AND  D(11)='1' )then
          cVar2S8S25P057nsss(0) <='1';
          else
          cVar2S8S25P057nsss(0) <='0';
          end if;
        if(cVar1S9S25N041P013P031N056(0)='1' AND  D(11)='0' AND D( 2)='1' AND A( 0)='0' )then
          cVar2S9S25N057P060P019nsss(0) <='1';
          else
          cVar2S9S25N057P060P019nsss(0) <='0';
          end if;
        if(cVar1S10S25N041P013N031P015(0)='1' AND  D( 9)='0' AND A( 0)='1' AND B(19)='0' )then
          cVar2S10S25P065P019P020nsss(0) <='1';
          else
          cVar2S10S25P065P019P020nsss(0) <='0';
          end if;
        if(cVar1S11S25N041P013N031P015(0)='1' AND  D( 9)='0' AND A( 0)='0' )then
          cVar2S11S25P065N019psss(0) <='1';
          else
          cVar2S11S25P065N019psss(0) <='0';
          end if;
        if(cVar1S12S25N041P013N031P015(0)='1' AND  D( 9)='1' AND E(11)='0' AND A( 1)='1' )then
          cVar2S12S25P065P059P017nsss(0) <='1';
          else
          cVar2S12S25P065P059P017nsss(0) <='0';
          end if;
        if(cVar1S13S25N041P013N031N015(0)='1' AND  E( 2)='0' AND A( 1)='1' AND E(14)='0' )then
          cVar2S13S25P062P017P047nsss(0) <='1';
          else
          cVar2S13S25P062P017P047nsss(0) <='0';
          end if;
        if(cVar1S14S25N041P013N031N015(0)='1' AND  E( 2)='0' AND A( 1)='0' AND D(11)='1' )then
          cVar2S14S25P062N017P057nsss(0) <='1';
          else
          cVar2S14S25P062N017P057nsss(0) <='0';
          end if;
        if(cVar1S15S25N041N013P031P044(0)='1' AND  B( 8)='1' )then
          cVar2S15S25P023nsss(0) <='1';
          else
          cVar2S15S25P023nsss(0) <='0';
          end if;
        if(cVar1S16S25N041N013P031P044(0)='1' AND  B( 8)='0' AND B(18)='1' )then
          cVar2S16S25N023P022nsss(0) <='1';
          else
          cVar2S16S25N023P022nsss(0) <='0';
          end if;
        if(cVar1S17S25N041N013P031N044(0)='1' AND  D( 1)='1' AND B( 1)='0' AND E( 2)='1' )then
          cVar2S17S25P064P037P062nsss(0) <='1';
          else
          cVar2S17S25P064P037P062nsss(0) <='0';
          end if;
        if(cVar1S18S25N041N013P031N044(0)='1' AND  D( 1)='0' AND B( 1)='1' AND D( 0)='1' )then
          cVar2S18S25N064P037P068nsss(0) <='1';
          else
          cVar2S18S25N064P037P068nsss(0) <='0';
          end if;
        if(cVar1S19S25N041N013P031N044(0)='1' AND  D( 1)='0' AND B( 1)='0' AND B(18)='1' )then
          cVar2S19S25N064N037P022nsss(0) <='1';
          else
          cVar2S19S25N064N037P022nsss(0) <='0';
          end if;
        if(cVar1S20S25N041N013P031P011(0)='1' AND  A(11)='0' AND E( 4)='1' )then
          cVar2S20S25P016P054nsss(0) <='1';
          else
          cVar2S20S25P016P054nsss(0) <='0';
          end if;
        if(cVar1S21S25N041N013P031P011(0)='1' AND  A(11)='0' AND E( 4)='0' AND D(11)='1' )then
          cVar2S21S25P016N054P057nsss(0) <='1';
          else
          cVar2S21S25P016N054P057nsss(0) <='0';
          end if;
        if(cVar1S22S25N041N013P031N011(0)='1' AND  A(13)='1' AND D( 3)='1' )then
          cVar2S22S25P012P056nsss(0) <='1';
          else
          cVar2S22S25P012P056nsss(0) <='0';
          end if;
        if(cVar1S1S26P068P041N020P005(0)='1' AND  B( 0)='1' )then
          cVar2S1S26P039nsss(0) <='1';
          else
          cVar2S1S26P039nsss(0) <='0';
          end if;
        if(cVar1S2S26P068P041N020P005(0)='1' AND  B( 0)='0' AND B( 8)='1' )then
          cVar2S2S26N039P023nsss(0) <='1';
          else
          cVar2S2S26N039P023nsss(0) <='0';
          end if;
        if(cVar1S3S26P068P041N020N005(0)='1' AND  A( 8)='1' )then
          cVar2S3S26P003nsss(0) <='1';
          else
          cVar2S3S26P003nsss(0) <='0';
          end if;
        if(cVar1S4S26P068P041N020N005(0)='1' AND  A( 8)='0' AND B(18)='1' )then
          cVar2S4S26N003P022nsss(0) <='1';
          else
          cVar2S4S26N003P022nsss(0) <='0';
          end if;
        if(cVar1S5S26P068N041P024P006(0)='1' AND  E(14)='1' )then
          cVar2S5S26P047nsss(0) <='1';
          else
          cVar2S5S26P047nsss(0) <='0';
          end if;
        if(cVar1S6S26P068N041P024P006(0)='1' AND  E(14)='0' AND D(14)='1' )then
          cVar2S6S26N047P045nsss(0) <='1';
          else
          cVar2S6S26N047P045nsss(0) <='0';
          end if;
        if(cVar1S7S26P068N041P024P006(0)='1' AND  E(14)='0' AND D(14)='0' AND E( 6)='1' )then
          cVar2S7S26N047N045P046nsss(0) <='1';
          else
          cVar2S7S26N047N045P046nsss(0) <='0';
          end if;
        if(cVar1S8S26P068N041P024N006(0)='1' AND  A( 6)='1' AND D(14)='1' )then
          cVar2S8S26P007P045nsss(0) <='1';
          else
          cVar2S8S26P007P045nsss(0) <='0';
          end if;
        if(cVar1S9S26P068N041P024N006(0)='1' AND  A( 6)='1' AND D(14)='0' AND D(13)='1' )then
          cVar2S9S26P007N045P049nsss(0) <='1';
          else
          cVar2S9S26P007N045P049nsss(0) <='0';
          end if;
        if(cVar1S10S26P068N041N024P023(0)='1' AND  A( 7)='1' AND E( 7)='1' )then
          cVar2S10S26P005P042nsss(0) <='1';
          else
          cVar2S10S26P005P042nsss(0) <='0';
          end if;
        if(cVar1S11S26P068N041N024P023(0)='1' AND  A( 7)='1' AND E( 7)='0' AND D(14)='1' )then
          cVar2S11S26P005N042P045nsss(0) <='1';
          else
          cVar2S11S26P005N042P045nsss(0) <='0';
          end if;
        if(cVar1S12S26P068N041N024P023(0)='1' AND  A( 7)='0' AND E( 7)='1' )then
          cVar2S12S26N005P042nsss(0) <='1';
          else
          cVar2S12S26N005P042nsss(0) <='0';
          end if;
        if(cVar1S13S26P068N041N024P023(0)='1' AND  A( 7)='0' AND E( 7)='0' AND A( 6)='1' )then
          cVar2S13S26N005N042P007nsss(0) <='1';
          else
          cVar2S13S26N005N042P007nsss(0) <='0';
          end if;
        if(cVar1S14S26P068N041N024N023(0)='1' AND  D(14)='0' AND E(15)='0' AND E( 7)='0' )then
          cVar2S14S26P045P043P042nsss(0) <='1';
          else
          cVar2S14S26P045P043P042nsss(0) <='0';
          end if;
        if(cVar1S15S26P068N041N024N023(0)='1' AND  D(14)='1' AND B(18)='1' )then
          cVar2S15S26P045P022nsss(0) <='1';
          else
          cVar2S15S26P045P022nsss(0) <='0';
          end if;
        if(cVar1S16S26P068N041N024N023(0)='1' AND  D(14)='1' AND B(18)='0' AND B( 7)='1' )then
          cVar2S16S26P045N022P025nsss(0) <='1';
          else
          cVar2S16S26P045N022P025nsss(0) <='0';
          end if;
        if(cVar1S17S26P068P065P019P061(0)='1' AND  D(14)='0' AND B( 6)='0' )then
          cVar2S17S26P045P027nsss(0) <='1';
          else
          cVar2S17S26P045P027nsss(0) <='0';
          end if;
        if(cVar1S18S26P068P065P019P061(0)='1' AND  D(14)='0' AND B( 6)='1' AND A( 2)='1' )then
          cVar2S18S26P045P027P015nsss(0) <='1';
          else
          cVar2S18S26P045P027P015nsss(0) <='0';
          end if;
        if(cVar1S19S26P068P065N019P037(0)='1' AND  E( 9)='0' AND A( 6)='0' AND D(10)='0' )then
          cVar2S19S26P067P007P061nsss(0) <='1';
          else
          cVar2S19S26P067P007P061nsss(0) <='0';
          end if;
        if(cVar1S20S26P068P065N019P037(0)='1' AND  E( 9)='0' AND A( 6)='1' AND A(13)='1' )then
          cVar2S20S26P067P007P012nsss(0) <='1';
          else
          cVar2S20S26P067P007P012nsss(0) <='0';
          end if;
        if(cVar1S21S26P068P065N019P037(0)='1' AND  E( 9)='1' AND E( 2)='1' )then
          cVar2S21S26P067P062nsss(0) <='1';
          else
          cVar2S21S26P067P062nsss(0) <='0';
          end if;
        if(cVar1S22S26P068P065N019N037(0)='1' AND  A(10)='1' AND E( 2)='0' AND A(16)='0' )then
          cVar2S22S26P018P062P006nsss(0) <='1';
          else
          cVar2S22S26P018P062P006nsss(0) <='0';
          end if;
        if(cVar1S23S26P068P065N019N037(0)='1' AND  A(10)='0' AND D( 8)='1' AND A(11)='1' )then
          cVar2S23S26N018P069P016nsss(0) <='1';
          else
          cVar2S23S26N018P069P016nsss(0) <='0';
          end if;
        if(cVar1S24S26P068P065N019N037(0)='1' AND  A(10)='0' AND D( 8)='0' AND D(11)='1' )then
          cVar2S24S26N018N069P057nsss(0) <='1';
          else
          cVar2S24S26N018N069P057nsss(0) <='0';
          end if;
        if(cVar1S25S26P068P065P069P036(0)='1' AND  A( 0)='1' )then
          cVar2S25S26P019nsss(0) <='1';
          else
          cVar2S25S26P019nsss(0) <='0';
          end if;
        if(cVar1S26S26P068P065P069P036(0)='1' AND  A( 0)='0' AND A( 1)='0' )then
          cVar2S26S26N019P017nsss(0) <='1';
          else
          cVar2S26S26N019P017nsss(0) <='0';
          end if;
        if(cVar1S27S26P068P065P069P036(0)='1' AND  D( 1)='0' AND A(11)='1' )then
          cVar2S27S26P064P016nsss(0) <='1';
          else
          cVar2S27S26P064P016nsss(0) <='0';
          end if;
        if(cVar1S28S26P068P065N069P016(0)='1' AND  B(12)='1' AND D( 1)='1' )then
          cVar2S28S26P034P064nsss(0) <='1';
          else
          cVar2S28S26P034P064nsss(0) <='0';
          end if;
        if(cVar1S29S26P068P065N069P016(0)='1' AND  B(12)='1' AND D( 1)='0' AND A( 0)='1' )then
          cVar2S29S26P034N064P019nsss(0) <='1';
          else
          cVar2S29S26P034N064P019nsss(0) <='0';
          end if;
        if(cVar1S30S26P068P065N069N016(0)='1' AND  A(12)='1' AND B(12)='1' )then
          cVar2S30S26P014P034nsss(0) <='1';
          else
          cVar2S30S26P014P034nsss(0) <='0';
          end if;
        if(cVar1S31S26P068P065N069N016(0)='1' AND  A(12)='0' AND E(10)='0' AND A(10)='1' )then
          cVar2S31S26N014P063P018nsss(0) <='1';
          else
          cVar2S31S26N014P063P018nsss(0) <='0';
          end if;
        if(cVar1S2S27P041P020N003N002(0)='1' AND  A(17)='1' )then
          cVar2S2S27P004nsss(0) <='1';
          else
          cVar2S2S27P004nsss(0) <='0';
          end if;
        if(cVar1S3S27P041P020N003N002(0)='1' AND  A(17)='0' AND A( 7)='1' )then
          cVar2S3S27N004P005nsss(0) <='1';
          else
          cVar2S3S27N004P005nsss(0) <='0';
          end if;
        if(cVar1S4S27P041N020P068P005(0)='1' AND  B( 0)='1' )then
          cVar2S4S27P039nsss(0) <='1';
          else
          cVar2S4S27P039nsss(0) <='0';
          end if;
        if(cVar1S5S27P041N020P068P005(0)='1' AND  B( 0)='0' AND B( 8)='1' )then
          cVar2S5S27N039P023nsss(0) <='1';
          else
          cVar2S5S27N039P023nsss(0) <='0';
          end if;
        if(cVar1S6S27P041N020P068N005(0)='1' AND  B(12)='0' AND D( 9)='0' )then
          cVar2S6S27P034P065nsss(0) <='1';
          else
          cVar2S6S27P034P065nsss(0) <='0';
          end if;
        if(cVar1S7S27P041N020P068P039(0)='1' AND  A( 0)='1' )then
          cVar2S7S27P019nsss(0) <='1';
          else
          cVar2S7S27P019nsss(0) <='0';
          end if;
        if(cVar1S9S27N041P024P006N047(0)='1' AND  D(14)='1' )then
          cVar2S9S27P045nsss(0) <='1';
          else
          cVar2S9S27P045nsss(0) <='0';
          end if;
        if(cVar1S10S27N041P024P006N047(0)='1' AND  D(14)='0' AND D( 6)='1' )then
          cVar2S10S27N045P044nsss(0) <='1';
          else
          cVar2S10S27N045P044nsss(0) <='0';
          end if;
        if(cVar1S11S27N041P024P006N047(0)='1' AND  D(14)='0' AND D( 6)='0' AND E( 6)='1' )then
          cVar2S11S27N045N044P046nsss(0) <='1';
          else
          cVar2S11S27N045N044P046nsss(0) <='0';
          end if;
        if(cVar1S12S27N041P024N006P049(0)='1' AND  D( 0)='0' AND A( 6)='1' )then
          cVar2S12S27P068P007nsss(0) <='1';
          else
          cVar2S12S27P068P007nsss(0) <='0';
          end if;
        if(cVar1S13S27N041P024N006P049(0)='1' AND  D( 0)='0' AND A( 6)='0' AND A( 1)='0' )then
          cVar2S13S27P068N007P017nsss(0) <='1';
          else
          cVar2S13S27P068N007P017nsss(0) <='0';
          end if;
        if(cVar1S14S27N041P024N006N049(0)='1' AND  D(14)='1' )then
          cVar2S14S27P045nsss(0) <='1';
          else
          cVar2S14S27P045nsss(0) <='0';
          end if;
        if(cVar1S15S27N041P024N006N049(0)='1' AND  D(14)='0' AND D( 0)='1' AND A( 4)='1' )then
          cVar2S15S27N045P068P011nsss(0) <='1';
          else
          cVar2S15S27N045P068P011nsss(0) <='0';
          end if;
        if(cVar1S16S27N041N024P023P005(0)='1' AND  E( 7)='1' )then
          cVar2S16S27P042nsss(0) <='1';
          else
          cVar2S16S27P042nsss(0) <='0';
          end if;
        if(cVar1S17S27N041N024P023P005(0)='1' AND  E( 7)='0' AND D(14)='1' )then
          cVar2S17S27N042P045nsss(0) <='1';
          else
          cVar2S17S27N042P045nsss(0) <='0';
          end if;
        if(cVar1S18S27N041N024P023N005(0)='1' AND  E( 7)='1' AND A(17)='1' )then
          cVar2S18S27P042P004nsss(0) <='1';
          else
          cVar2S18S27P042P004nsss(0) <='0';
          end if;
        if(cVar1S19S27N041N024P023N005(0)='1' AND  E( 7)='1' AND A(17)='0' AND A( 1)='0' )then
          cVar2S19S27P042N004P017nsss(0) <='1';
          else
          cVar2S19S27P042N004P017nsss(0) <='0';
          end if;
        if(cVar1S20S27N041N024P023N005(0)='1' AND  E( 7)='0' AND A( 6)='1' )then
          cVar2S20S27N042P007nsss(0) <='1';
          else
          cVar2S20S27N042P007nsss(0) <='0';
          end if;
        if(cVar1S21S27N041N024P023N005(0)='1' AND  E( 7)='0' AND A( 6)='0' AND A(15)='1' )then
          cVar2S21S27N042N007P008nsss(0) <='1';
          else
          cVar2S21S27N042N007P008nsss(0) <='0';
          end if;
        if(cVar1S22S27N041N024N023P050(0)='1' AND  A( 5)='1' AND B( 6)='1' AND A( 4)='0' )then
          cVar2S22S27P009P027P011nsss(0) <='1';
          else
          cVar2S22S27P009P027P011nsss(0) <='0';
          end if;
        if(cVar1S23S27N041N024N023P050(0)='1' AND  A( 5)='1' AND B( 6)='0' AND B( 5)='1' )then
          cVar2S23S27P009N027P029nsss(0) <='1';
          else
          cVar2S23S27P009N027P029nsss(0) <='0';
          end if;
        if(cVar1S24S27N041N024N023P050(0)='1' AND  A( 5)='0' AND B(16)='1' )then
          cVar2S24S27N009P026nsss(0) <='1';
          else
          cVar2S24S27N009P026nsss(0) <='0';
          end if;
        if(cVar1S25S27N041N024N023P050(0)='1' AND  A( 5)='0' AND B(16)='0' AND E(12)='1' )then
          cVar2S25S27N009N026P055nsss(0) <='1';
          else
          cVar2S25S27N009N026P055nsss(0) <='0';
          end if;
        if(cVar1S26S27N041N024N023N050(0)='1' AND  A( 7)='0' AND D( 8)='1' AND B(11)='1' )then
          cVar2S26S27P005P069P036nsss(0) <='1';
          else
          cVar2S26S27P005P069P036nsss(0) <='0';
          end if;
        if(cVar1S27S27N041N024N023N050(0)='1' AND  A( 7)='1' AND B(18)='1' )then
          cVar2S27S27P005P022nsss(0) <='1';
          else
          cVar2S27S27P005P022nsss(0) <='0';
          end if;
        if(cVar1S28S27N041N024N023N050(0)='1' AND  A( 7)='1' AND B(18)='0' AND B( 7)='1' )then
          cVar2S28S27P005N022P025nsss(0) <='1';
          else
          cVar2S28S27P005N022P025nsss(0) <='0';
          end if;
        if(cVar1S2S28P024P006N047N045(0)='1' AND  D( 6)='1' )then
          cVar2S2S28P044nsss(0) <='1';
          else
          cVar2S2S28P044nsss(0) <='0';
          end if;
        if(cVar1S3S28P024P006N047N045(0)='1' AND  D( 6)='0' AND D( 5)='1' )then
          cVar2S3S28N044P048nsss(0) <='1';
          else
          cVar2S3S28N044P048nsss(0) <='0';
          end if;
        if(cVar1S4S28P024N006P068P034(0)='1' AND  A( 6)='1' )then
          cVar2S4S28P007nsss(0) <='1';
          else
          cVar2S4S28P007nsss(0) <='0';
          end if;
        if(cVar1S5S28P024N006P068P034(0)='1' AND  A( 6)='0' AND B( 7)='0' )then
          cVar2S5S28N007P025nsss(0) <='1';
          else
          cVar2S5S28N007P025nsss(0) <='0';
          end if;
        if(cVar1S6S28P024N006P068P034(0)='1' AND  A( 2)='1' )then
          cVar2S6S28P015nsss(0) <='1';
          else
          cVar2S6S28P015nsss(0) <='0';
          end if;
        if(cVar1S10S28N024P040N002N004(0)='1' AND  A( 7)='1' )then
          cVar2S10S28P005nsss(0) <='1';
          else
          cVar2S10S28P005nsss(0) <='0';
          end if;
        if(cVar1S11S28N024P040N002N004(0)='1' AND  A( 7)='0' AND A( 8)='1' AND A( 2)='0' )then
          cVar2S11S28N005P003P015nsss(0) <='1';
          else
          cVar2S11S28N005P003P015nsss(0) <='0';
          end if;
        if(cVar1S12S28N024N040P044P023(0)='1' AND  A( 7)='1' )then
          cVar2S12S28P005nsss(0) <='1';
          else
          cVar2S12S28P005nsss(0) <='0';
          end if;
        if(cVar1S13S28N024N040P044P023(0)='1' AND  A( 7)='0' AND A(17)='1' )then
          cVar2S13S28N005P004nsss(0) <='1';
          else
          cVar2S13S28N005P004nsss(0) <='0';
          end if;
        if(cVar1S14S28N024N040P044P023(0)='1' AND  A( 7)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S14S28N005N004P007nsss(0) <='1';
          else
          cVar2S14S28N005N004P007nsss(0) <='0';
          end if;
        if(cVar1S15S28N024N040P044N023(0)='1' AND  B( 7)='1' AND A(12)='0' )then
          cVar2S15S28P025P014nsss(0) <='1';
          else
          cVar2S15S28P025P014nsss(0) <='0';
          end if;
        if(cVar1S16S28N024N040P044N023(0)='1' AND  B( 7)='0' AND E( 4)='1' )then
          cVar2S16S28N025P054nsss(0) <='1';
          else
          cVar2S16S28N025P054nsss(0) <='0';
          end if;
        if(cVar1S17S28N024N040P044N023(0)='1' AND  B( 7)='0' AND E( 4)='0' AND B(18)='1' )then
          cVar2S17S28N025N054P022nsss(0) <='1';
          else
          cVar2S17S28N025N054P022nsss(0) <='0';
          end if;
        if(cVar1S18S28N024N040N044P042(0)='1' AND  B( 9)='0' )then
          cVar2S18S28P021nsss(0) <='1';
          else
          cVar2S18S28P021nsss(0) <='0';
          end if;
        if(cVar1S19S28N024N040N044P042(0)='1' AND  B( 9)='1' AND B( 0)='1' )then
          cVar2S19S28P021P039nsss(0) <='1';
          else
          cVar2S19S28P021P039nsss(0) <='0';
          end if;
        if(cVar1S20S28N024N040N044P042(0)='1' AND  B( 9)='1' AND B( 0)='0' AND E(12)='1' )then
          cVar2S20S28P021N039P055nsss(0) <='1';
          else
          cVar2S20S28P021N039P055nsss(0) <='0';
          end if;
        if(cVar1S21S28N024N040N044P042(0)='1' AND  E( 3)='1' )then
          cVar2S21S28P058nsss(0) <='1';
          else
          cVar2S21S28P058nsss(0) <='0';
          end if;
        if(cVar1S22S28N024N040N044P042(0)='1' AND  E( 3)='0' AND E(15)='1' )then
          cVar2S22S28N058P043nsss(0) <='1';
          else
          cVar2S22S28N058P043nsss(0) <='0';
          end if;
        if(cVar1S2S29P024P006N047N045(0)='1' AND  D( 6)='1' )then
          cVar2S2S29P044nsss(0) <='1';
          else
          cVar2S2S29P044nsss(0) <='0';
          end if;
        if(cVar1S3S29P024P006N047N045(0)='1' AND  D( 6)='0' AND D( 5)='1' )then
          cVar2S3S29N044P048nsss(0) <='1';
          else
          cVar2S3S29N044P048nsss(0) <='0';
          end if;
        if(cVar1S4S29P024N006P068P007(0)='1' AND  D(14)='1' )then
          cVar2S4S29P045nsss(0) <='1';
          else
          cVar2S4S29P045nsss(0) <='0';
          end if;
        if(cVar1S5S29P024N006P068P007(0)='1' AND  D(14)='0' AND D(13)='1' )then
          cVar2S5S29N045P049nsss(0) <='1';
          else
          cVar2S5S29N045P049nsss(0) <='0';
          end if;
        if(cVar1S6S29P024N006P068N007(0)='1' AND  B( 7)='0' AND D(11)='0' )then
          cVar2S6S29P025P057nsss(0) <='1';
          else
          cVar2S6S29P025P057nsss(0) <='0';
          end if;
        if(cVar1S8S29P024N006P068N012(0)='1' AND  A(15)='1' )then
          cVar2S8S29P008nsss(0) <='1';
          else
          cVar2S8S29P008nsss(0) <='0';
          end if;
        if(cVar1S10S29N024P040N002P034(0)='1' AND  B( 9)='1' AND A( 8)='1' )then
          cVar2S10S29P021P003nsss(0) <='1';
          else
          cVar2S10S29P021P003nsss(0) <='0';
          end if;
        if(cVar1S11S29N024P040N002P034(0)='1' AND  B( 9)='1' AND A( 8)='0' AND A( 7)='1' )then
          cVar2S11S29P021N003P005nsss(0) <='1';
          else
          cVar2S11S29P021N003P005nsss(0) <='0';
          end if;
        if(cVar1S12S29N024P040N002P034(0)='1' AND  B( 9)='0' AND E( 1)='0' )then
          cVar2S12S29N021P066nsss(0) <='1';
          else
          cVar2S12S29N021P066nsss(0) <='0';
          end if;
        if(cVar1S13S29N024P040N002P034(0)='1' AND  B( 9)='0' AND E( 1)='1' AND A( 1)='1' )then
          cVar2S13S29N021P066P017nsss(0) <='1';
          else
          cVar2S13S29N021P066P017nsss(0) <='0';
          end if;
        if(cVar1S14S29N024N040P044P023(0)='1' AND  A( 7)='1' )then
          cVar2S14S29P005nsss(0) <='1';
          else
          cVar2S14S29P005nsss(0) <='0';
          end if;
        if(cVar1S15S29N024N040P044P023(0)='1' AND  A( 7)='0' AND A(17)='1' )then
          cVar2S15S29N005P004nsss(0) <='1';
          else
          cVar2S15S29N005P004nsss(0) <='0';
          end if;
        if(cVar1S16S29N024N040P044P023(0)='1' AND  A( 7)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S16S29N005N004P007nsss(0) <='1';
          else
          cVar2S16S29N005N004P007nsss(0) <='0';
          end if;
        if(cVar1S17S29N024N040P044N023(0)='1' AND  B( 7)='1' AND A( 2)='0' )then
          cVar2S17S29P025P015nsss(0) <='1';
          else
          cVar2S17S29P025P015nsss(0) <='0';
          end if;
        if(cVar1S18S29N024N040P044N023(0)='1' AND  B( 7)='0' )then
          cVar2S18S29N025psss(0) <='1';
          else
          cVar2S18S29N025psss(0) <='0';
          end if;
        if(cVar1S19S29N024N040N044P041(0)='1' AND  B(19)='1' AND A( 8)='1' )then
          cVar2S19S29P020P003nsss(0) <='1';
          else
          cVar2S19S29P020P003nsss(0) <='0';
          end if;
        if(cVar1S20S29N024N040N044P041(0)='1' AND  B(19)='1' AND A( 8)='0' AND A(18)='1' )then
          cVar2S20S29P020N003P002nsss(0) <='1';
          else
          cVar2S20S29P020N003P002nsss(0) <='0';
          end if;
        if(cVar1S21S29N024N040N044P041(0)='1' AND  B(19)='0' AND A( 7)='1' )then
          cVar2S21S29N020P005nsss(0) <='1';
          else
          cVar2S21S29N020P005nsss(0) <='0';
          end if;
        if(cVar1S22S29N024N040N044P041(0)='1' AND  B(19)='0' AND A( 7)='0' AND A( 8)='1' )then
          cVar2S22S29N020N005P003nsss(0) <='1';
          else
          cVar2S22S29N020N005P003nsss(0) <='0';
          end if;
        if(cVar1S23S29N024N040N044N041(0)='1' AND  B( 0)='0' AND A( 7)='1' AND E(15)='1' )then
          cVar2S23S29P039P005P043nsss(0) <='1';
          else
          cVar2S23S29P039P005P043nsss(0) <='0';
          end if;
        if(cVar1S1S30P067P018P048N025(0)='1' AND  B( 6)='1' )then
          cVar2S1S30P027nsss(0) <='1';
          else
          cVar2S1S30P027nsss(0) <='0';
          end if;
        if(cVar1S2S30P067P018P048N025(0)='1' AND  B( 6)='0' AND B(17)='1' )then
          cVar2S2S30N027P024nsss(0) <='1';
          else
          cVar2S2S30N027P024nsss(0) <='0';
          end if;
        if(cVar1S3S30P067P018P048N025(0)='1' AND  B( 6)='0' AND B(17)='0' AND A( 3)='1' )then
          cVar2S3S30N027N024P013nsss(0) <='1';
          else
          cVar2S3S30N027N024P013nsss(0) <='0';
          end if;
        if(cVar1S4S30P067P018N048P014(0)='1' AND  B(12)='1' AND A( 2)='0' AND B( 2)='0' )then
          cVar2S4S30P034P015P035nsss(0) <='1';
          else
          cVar2S4S30P034P015P035nsss(0) <='0';
          end if;
        if(cVar1S5S30P067P018N048P014(0)='1' AND  B(12)='1' AND A( 2)='1' AND E(10)='1' )then
          cVar2S5S30P034P015P063nsss(0) <='1';
          else
          cVar2S5S30P034P015P063nsss(0) <='0';
          end if;
        if(cVar1S6S30P067P018N048P014(0)='1' AND  B(12)='0' AND B(13)='1' AND D( 9)='0' )then
          cVar2S6S30N034P032P065nsss(0) <='1';
          else
          cVar2S6S30N034P032P065nsss(0) <='0';
          end if;
        if(cVar1S7S30P067P018N048P014(0)='1' AND  B(12)='0' AND B(13)='0' )then
          cVar2S7S30N034N032psss(0) <='1';
          else
          cVar2S7S30N034N032psss(0) <='0';
          end if;
        if(cVar1S8S30P067P018N048N014(0)='1' AND  B(14)='1' AND B( 4)='0' )then
          cVar2S8S30P030P031nsss(0) <='1';
          else
          cVar2S8S30P030P031nsss(0) <='0';
          end if;
        if(cVar1S9S30P067P018N048N014(0)='1' AND  B(14)='0' )then
          cVar2S9S30N030psss(0) <='1';
          else
          cVar2S9S30N030psss(0) <='0';
          end if;
        if(cVar1S10S30P067P018P060P011(0)='1' AND  A( 8)='1' )then
          cVar2S10S30P003nsss(0) <='1';
          else
          cVar2S10S30P003nsss(0) <='0';
          end if;
        if(cVar1S11S30P067P018P060P011(0)='1' AND  A( 8)='0' AND B( 5)='1' )then
          cVar2S11S30N003P029nsss(0) <='1';
          else
          cVar2S11S30N003P029nsss(0) <='0';
          end if;
        if(cVar1S12S30P067P018P060P011(0)='1' AND  A( 8)='0' AND B( 5)='0' AND D( 8)='0' )then
          cVar2S12S30N003N029P069nsss(0) <='1';
          else
          cVar2S12S30N003N029P069nsss(0) <='0';
          end if;
        if(cVar1S13S30P067P018P060N011(0)='1' AND  E( 4)='0' AND B(17)='1' )then
          cVar2S13S30P054P024nsss(0) <='1';
          else
          cVar2S13S30P054P024nsss(0) <='0';
          end if;
        if(cVar1S14S30P067P018P060N011(0)='1' AND  E( 4)='0' AND B(17)='0' AND D( 7)='1' )then
          cVar2S14S30P054N024P040nsss(0) <='1';
          else
          cVar2S14S30P054N024P040nsss(0) <='0';
          end if;
        if(cVar1S15S30P067P018P060N011(0)='1' AND  E( 4)='1' AND A( 3)='1' AND B( 4)='1' )then
          cVar2S15S30P054P013P031nsss(0) <='1';
          else
          cVar2S15S30P054P013P031nsss(0) <='0';
          end if;
        if(cVar1S16S30P067P018P060P013(0)='1' AND  B( 3)='1' )then
          cVar2S16S30P033nsss(0) <='1';
          else
          cVar2S16S30P033nsss(0) <='0';
          end if;
        if(cVar1S17S30P067P018P060P013(0)='1' AND  B( 3)='0' AND E( 2)='0' AND A( 1)='0' )then
          cVar2S17S30N033P062P017nsss(0) <='1';
          else
          cVar2S17S30N033P062P017nsss(0) <='0';
          end if;
        if(cVar1S18S30P067P018P060N013(0)='1' AND  E( 5)='1' )then
          cVar2S18S30P050nsss(0) <='1';
          else
          cVar2S18S30P050nsss(0) <='0';
          end if;
        if(cVar1S19S30P067P018P060N013(0)='1' AND  E( 5)='0' AND B( 2)='1' AND E( 3)='0' )then
          cVar2S19S30N050P035P058nsss(0) <='1';
          else
          cVar2S19S30N050P035P058nsss(0) <='0';
          end if;
        if(cVar1S20S30P067P069P018P016(0)='1' AND  D( 2)='0' AND D( 4)='1' )then
          cVar2S20S30P060P052nsss(0) <='1';
          else
          cVar2S20S30P060P052nsss(0) <='0';
          end if;
        if(cVar1S21S30P067P069P018P016(0)='1' AND  D( 2)='0' AND D( 4)='0' AND A( 5)='0' )then
          cVar2S21S30P060N052P009nsss(0) <='1';
          else
          cVar2S21S30P060N052P009nsss(0) <='0';
          end if;
        if(cVar1S22S30P067P069P018P016(0)='1' AND  D( 2)='1' AND A( 1)='1' )then
          cVar2S22S30P060P017nsss(0) <='1';
          else
          cVar2S22S30P060P017nsss(0) <='0';
          end if;
        if(cVar1S23S30P067P069P018P016(0)='1' AND  B( 4)='0' AND D( 5)='0' AND D( 1)='0' )then
          cVar2S23S30P031P048P064nsss(0) <='1';
          else
          cVar2S23S30P031P048P064nsss(0) <='0';
          end if;
        if(cVar1S24S30P067P069N018P019(0)='1' AND  B(11)='0' )then
          cVar2S24S30P036nsss(0) <='1';
          else
          cVar2S24S30P036nsss(0) <='0';
          end if;
        if(cVar1S25S30P067P069N018P019(0)='1' AND  B(11)='1' AND E( 1)='0' AND A(13)='0' )then
          cVar2S25S30P036P066P012nsss(0) <='1';
          else
          cVar2S25S30P036P066P012nsss(0) <='0';
          end if;
        if(cVar1S26S30P067P069N018N019(0)='1' AND  A(11)='1' AND B(11)='1' AND B( 1)='0' )then
          cVar2S26S30P016P036P037nsss(0) <='1';
          else
          cVar2S26S30P016P036P037nsss(0) <='0';
          end if;
        if(cVar1S27S30P067P069N018N019(0)='1' AND  A(11)='1' AND B(11)='0' AND D( 0)='1' )then
          cVar2S27S30P016N036P068nsss(0) <='1';
          else
          cVar2S27S30P016N036P068nsss(0) <='0';
          end if;
        if(cVar1S28S30P067P069N018N019(0)='1' AND  A(11)='0' AND A( 1)='1' AND A( 2)='0' )then
          cVar2S28S30N016P017P015nsss(0) <='1';
          else
          cVar2S28S30N016P017P015nsss(0) <='0';
          end if;
        if(cVar1S30S30P067N069P065P063(0)='1' AND  B(12)='1' )then
          cVar2S30S30P034nsss(0) <='1';
          else
          cVar2S30S30P034nsss(0) <='0';
          end if;
        if(cVar1S32S30P067N069N065N052(0)='1' AND  E(10)='0' AND D(10)='1' )then
          cVar2S32S30P063P061nsss(0) <='1';
          else
          cVar2S32S30P063P061nsss(0) <='0';
          end if;
        if(cVar1S0S31P018P060P054P062(0)='1' AND  E(10)='0' AND A(11)='0' )then
          cVar2S0S31P063P016nsss(0) <='1';
          else
          cVar2S0S31P063P016nsss(0) <='0';
          end if;
        if(cVar1S1S31P018P060P054P062(0)='1' AND  E(10)='0' AND A(11)='1' AND D( 8)='0' )then
          cVar2S1S31P063P016P069nsss(0) <='1';
          else
          cVar2S1S31P063P016P069nsss(0) <='0';
          end if;
        if(cVar1S2S31P018P060P054P062(0)='1' AND  E(10)='1' AND B(12)='1' AND D( 0)='0' )then
          cVar2S2S31P063P034P068nsss(0) <='1';
          else
          cVar2S2S31P063P034P068nsss(0) <='0';
          end if;
        if(cVar1S3S31P018P060P054P062(0)='1' AND  D( 1)='1' AND E( 5)='1' )then
          cVar2S3S31P064P050nsss(0) <='1';
          else
          cVar2S3S31P064P050nsss(0) <='0';
          end if;
        if(cVar1S4S31P018P060P054P062(0)='1' AND  D( 1)='1' AND E( 5)='0' AND E(11)='0' )then
          cVar2S4S31P064N050P059nsss(0) <='1';
          else
          cVar2S4S31P064N050P059nsss(0) <='0';
          end if;
        if(cVar1S5S31P018P060P054P062(0)='1' AND  D( 1)='0' AND A( 2)='1' AND A( 1)='0' )then
          cVar2S5S31N064P015P017nsss(0) <='1';
          else
          cVar2S5S31N064P015P017nsss(0) <='0';
          end if;
        if(cVar1S6S31P018P060P054P011(0)='1' AND  A( 2)='0' )then
          cVar2S6S31P015nsss(0) <='1';
          else
          cVar2S6S31P015nsss(0) <='0';
          end if;
        if(cVar1S7S31P018P060P054N011(0)='1' AND  D( 9)='0' AND A( 3)='1' AND D( 3)='1' )then
          cVar2S7S31P065P013P056nsss(0) <='1';
          else
          cVar2S7S31P065P013P056nsss(0) <='0';
          end if;
        if(cVar1S9S31P018P060P029N050(0)='1' AND  B(14)='0' AND A(12)='1' AND B(13)='1' )then
          cVar2S9S31P030P014P032nsss(0) <='1';
          else
          cVar2S9S31P030P014P032nsss(0) <='0';
          end if;
        if(cVar1S10S31P018P060P029N050(0)='1' AND  B(14)='0' AND A(12)='0' AND A( 2)='1' )then
          cVar2S10S31P030N014P015nsss(0) <='1';
          else
          cVar2S10S31P030N014P015nsss(0) <='0';
          end if;
        if(cVar1S12S31N018P048P025N007(0)='1' AND  A(16)='1' )then
          cVar2S12S31P006nsss(0) <='1';
          else
          cVar2S12S31P006nsss(0) <='0';
          end if;
        if(cVar1S13S31N018P048P025N007(0)='1' AND  A(16)='0' AND A( 5)='1' )then
          cVar2S13S31N006P009nsss(0) <='1';
          else
          cVar2S13S31N006P009nsss(0) <='0';
          end if;
        if(cVar1S15S31N018N048P014P034(0)='1' AND  B( 3)='0' AND B( 2)='0' )then
          cVar2S15S31P033P035nsss(0) <='1';
          else
          cVar2S15S31P033P035nsss(0) <='0';
          end if;
        if(cVar1S16S31N018N048P014N034(0)='1' AND  B(13)='1' AND A(14)='0' )then
          cVar2S16S31P032P010nsss(0) <='1';
          else
          cVar2S16S31P032P010nsss(0) <='0';
          end if;
        if(cVar1S17S31N018N048P014N034(0)='1' AND  B(13)='0' AND A(15)='1' AND A(16)='0' )then
          cVar2S17S31N032P008P006nsss(0) <='1';
          else
          cVar2S17S31N032P008P006nsss(0) <='0';
          end if;
        if(cVar1S18S31N018N048P014N034(0)='1' AND  B(13)='0' AND A(15)='0' AND A(13)='1' )then
          cVar2S18S31N032N008P012nsss(0) <='1';
          else
          cVar2S18S31N032N008P012nsss(0) <='0';
          end if;
        if(cVar1S19S31N018N048N014P030(0)='1' AND  A(13)='1' AND A(11)='0' AND A( 4)='0' )then
          cVar2S19S31P012P016P011nsss(0) <='1';
          else
          cVar2S19S31P012P016P011nsss(0) <='0';
          end if;
        if(cVar1S20S31N018N048N014P030(0)='1' AND  A(13)='1' AND A(11)='1' AND A( 2)='1' )then
          cVar2S20S31P012P016P015nsss(0) <='1';
          else
          cVar2S20S31P012P016P015nsss(0) <='0';
          end if;
        if(cVar1S21S31N018N048N014P030(0)='1' AND  A(13)='0' AND A(14)='1' )then
          cVar2S21S31N012P010nsss(0) <='1';
          else
          cVar2S21S31N012P010nsss(0) <='0';
          end if;
        if(cVar1S22S31N018N048N014P030(0)='1' AND  A(13)='0' AND A(14)='0' AND A( 3)='1' )then
          cVar2S22S31N012N010P013nsss(0) <='1';
          else
          cVar2S22S31N012N010P013nsss(0) <='0';
          end if;
        if(cVar1S23S31N018N048N014N030(0)='1' AND  B( 8)='1' AND A( 7)='1' )then
          cVar2S23S31P023P005nsss(0) <='1';
          else
          cVar2S23S31P023P005nsss(0) <='0';
          end if;
        if(cVar1S24S31N018N048N014N030(0)='1' AND  B( 8)='1' AND A( 7)='0' AND E( 7)='1' )then
          cVar2S24S31P023N005P042nsss(0) <='1';
          else
          cVar2S24S31P023N005P042nsss(0) <='0';
          end if;
        if(cVar1S25S31N018N048N014N030(0)='1' AND  B( 8)='0' AND A( 7)='0' AND A( 2)='1' )then
          cVar2S25S31N023P005P015nsss(0) <='1';
          else
          cVar2S25S31N023P005P015nsss(0) <='0';
          end if;
        if(cVar1S26S31N018N048N014N030(0)='1' AND  B( 8)='0' AND A( 7)='1' AND B( 9)='1' )then
          cVar2S26S31N023P005P021nsss(0) <='1';
          else
          cVar2S26S31N023P005P021nsss(0) <='0';
          end if;
        if(cVar1S1S32P015P018P040N021(0)='1' AND  B(19)='1' )then
          cVar2S1S32P020nsss(0) <='1';
          else
          cVar2S1S32P020nsss(0) <='0';
          end if;
        if(cVar1S2S32P015P018P040N021(0)='1' AND  B(19)='0' AND B( 8)='1' )then
          cVar2S2S32N020P023nsss(0) <='1';
          else
          cVar2S2S32N020P023nsss(0) <='0';
          end if;
        if(cVar1S3S32P015P018P040N021(0)='1' AND  B(19)='0' AND B( 8)='0' AND B(18)='1' )then
          cVar2S3S32N020N023P022nsss(0) <='1';
          else
          cVar2S3S32N020N023P022nsss(0) <='0';
          end if;
        if(cVar1S4S32P015P018N040P063(0)='1' AND  A(11)='1' AND A(13)='0' AND A(14)='0' )then
          cVar2S4S32P016P012P010nsss(0) <='1';
          else
          cVar2S4S32P016P012P010nsss(0) <='0';
          end if;
        if(cVar1S5S32P015P018N040P063(0)='1' AND  A(11)='1' AND A(13)='1' AND B(12)='1' )then
          cVar2S5S32P016P012P034nsss(0) <='1';
          else
          cVar2S5S32P016P012P034nsss(0) <='0';
          end if;
        if(cVar1S6S32P015P018N040P063(0)='1' AND  A(11)='0' AND A( 1)='1' AND A( 0)='0' )then
          cVar2S6S32N016P017P019nsss(0) <='1';
          else
          cVar2S6S32N016P017P019nsss(0) <='0';
          end if;
        if(cVar1S7S32P015P018N040P063(0)='1' AND  A(11)='0' AND A( 1)='0' AND A(12)='1' )then
          cVar2S7S32N016N017P014nsss(0) <='1';
          else
          cVar2S7S32N016N017P014nsss(0) <='0';
          end if;
        if(cVar1S8S32P015P018N040N063(0)='1' AND  A(11)='0' AND B(11)='0' )then
          cVar2S8S32P016P036nsss(0) <='1';
          else
          cVar2S8S32P016P036nsss(0) <='0';
          end if;
        if(cVar1S9S32P015P018N040N063(0)='1' AND  A(11)='0' AND B(11)='1' AND A( 1)='1' )then
          cVar2S9S32P016P036P017nsss(0) <='1';
          else
          cVar2S9S32P016P036P017nsss(0) <='0';
          end if;
        if(cVar1S10S32P015P018N040N063(0)='1' AND  A(11)='1' AND E( 2)='1' AND A(13)='0' )then
          cVar2S10S32P016P062P012nsss(0) <='1';
          else
          cVar2S10S32P016P062P012nsss(0) <='0';
          end if;
        if(cVar1S11S32P015P018N040N063(0)='1' AND  A(11)='1' AND E( 2)='0' AND B(11)='1' )then
          cVar2S11S32P016N062P036nsss(0) <='1';
          else
          cVar2S11S32P016N062P036nsss(0) <='0';
          end if;
        if(cVar1S12S32P015P018P004P062(0)='1' AND  D(11)='0' AND A( 1)='1' )then
          cVar2S12S32P057P017nsss(0) <='1';
          else
          cVar2S12S32P057P017nsss(0) <='0';
          end if;
        if(cVar1S13S32P015P018P004P062(0)='1' AND  D(11)='0' AND A( 1)='0' AND D( 8)='1' )then
          cVar2S13S32P057N017P069nsss(0) <='1';
          else
          cVar2S13S32P057N017P069nsss(0) <='0';
          end if;
        if(cVar1S14S32P015P018P004P062(0)='1' AND  D(11)='1' AND A( 3)='1' AND B(14)='1' )then
          cVar2S14S32P057P013P030nsss(0) <='1';
          else
          cVar2S14S32P057P013P030nsss(0) <='0';
          end if;
        if(cVar1S15S32P015P018P004P062(0)='1' AND  D(11)='1' AND A( 3)='0' AND E(13)='1' )then
          cVar2S15S32P057N013P051nsss(0) <='1';
          else
          cVar2S15S32P057N013P051nsss(0) <='0';
          end if;
        if(cVar1S16S32P015P018P004P062(0)='1' AND  D( 9)='0' AND B(11)='1' AND B( 1)='0' )then
          cVar2S16S32P065P036P037nsss(0) <='1';
          else
          cVar2S16S32P065P036P037nsss(0) <='0';
          end if;
        if(cVar1S17S32P015P018P004P062(0)='1' AND  D( 9)='1' AND B( 1)='0' AND A( 0)='1' )then
          cVar2S17S32P065P037P019nsss(0) <='1';
          else
          cVar2S17S32P065P037P019nsss(0) <='0';
          end if;
        if(cVar1S19S32P015P018P004N041(0)='1' AND  A(16)='1' )then
          cVar2S19S32P006nsss(0) <='1';
          else
          cVar2S19S32P006nsss(0) <='0';
          end if;
        if(cVar1S20S32P015P018P004N041(0)='1' AND  A(16)='0' AND E( 7)='1' )then
          cVar2S20S32N006P042nsss(0) <='1';
          else
          cVar2S20S32N006P042nsss(0) <='0';
          end if;
        if(cVar1S21S32P015P018P004N041(0)='1' AND  A(16)='0' AND E( 7)='0' AND D(14)='1' )then
          cVar2S21S32N006N042P045nsss(0) <='1';
          else
          cVar2S21S32N006N042P045nsss(0) <='0';
          end if;
        if(cVar1S22S32P015P017P060P063(0)='1' AND  B( 3)='1' AND A(10)='0' AND A(11)='0' )then
          cVar2S22S32P033P018P016nsss(0) <='1';
          else
          cVar2S22S32P033P018P016nsss(0) <='0';
          end if;
        if(cVar1S23S32P015P017P060P063(0)='1' AND  B( 3)='1' AND A(10)='1' AND D(10)='1' )then
          cVar2S23S32P033P018P061nsss(0) <='1';
          else
          cVar2S23S32P033P018P061nsss(0) <='0';
          end if;
        if(cVar1S24S32P015P017P060P063(0)='1' AND  B( 3)='0' AND B( 2)='1' AND E( 3)='0' )then
          cVar2S24S32N033P035P058nsss(0) <='1';
          else
          cVar2S24S32N033P035P058nsss(0) <='0';
          end if;
        if(cVar1S25S32P015P017P060P063(0)='1' AND  B( 3)='0' AND B( 2)='0' AND B( 1)='1' )then
          cVar2S25S32N033N035P037nsss(0) <='1';
          else
          cVar2S25S32N033N035P037nsss(0) <='0';
          end if;
        if(cVar1S26S32P015P017N060P018(0)='1' AND  A(14)='0' )then
          cVar2S26S32P010nsss(0) <='1';
          else
          cVar2S26S32P010nsss(0) <='0';
          end if;
        if(cVar1S27S32P015P017N060P018(0)='1' AND  A(14)='1' AND E(12)='1' )then
          cVar2S27S32P010P055nsss(0) <='1';
          else
          cVar2S27S32P010P055nsss(0) <='0';
          end if;
        if(cVar1S28S32P015P017N060N018(0)='1' AND  D( 1)='1' AND B( 2)='1' AND A( 3)='0' )then
          cVar2S28S32P064P035P013nsss(0) <='1';
          else
          cVar2S28S32P064P035P013nsss(0) <='0';
          end if;
        if(cVar1S29S32P015P017N060N018(0)='1' AND  D( 1)='1' AND B( 2)='0' AND A(11)='1' )then
          cVar2S29S32P064N035P016nsss(0) <='1';
          else
          cVar2S29S32P064N035P016nsss(0) <='0';
          end if;
        if(cVar1S30S32P015P017N060N018(0)='1' AND  D( 1)='0' AND A( 6)='1' )then
          cVar2S30S32N064P007nsss(0) <='1';
          else
          cVar2S30S32N064P007nsss(0) <='0';
          end if;
        if(cVar1S31S32P015P017N060N018(0)='1' AND  D( 1)='0' AND A( 6)='0' AND A(13)='1' )then
          cVar2S31S32N064N007P012nsss(0) <='1';
          else
          cVar2S31S32N064N007P012nsss(0) <='0';
          end if;
        if(cVar1S33S32P015P017P008P066(0)='1' AND  A(13)='0' AND A(10)='1' )then
          cVar2S33S32P012P018nsss(0) <='1';
          else
          cVar2S33S32P012P018nsss(0) <='0';
          end if;
        if(cVar1S34S32P015P017N008P056(0)='1' AND  D(13)='1' AND A( 3)='0' )then
          cVar2S34S32P049P013nsss(0) <='1';
          else
          cVar2S34S32P049P013nsss(0) <='0';
          end if;
        if(cVar1S35S32P015P017N008P056(0)='1' AND  D(13)='0' AND A(12)='1' AND B(13)='1' )then
          cVar2S35S32N049P014P032nsss(0) <='1';
          else
          cVar2S35S32N049P014P032nsss(0) <='0';
          end if;
        if(cVar1S36S32P015P017N008P056(0)='1' AND  E( 1)='1' )then
          cVar2S36S32P066nsss(0) <='1';
          else
          cVar2S36S32P066nsss(0) <='0';
          end if;
        if(cVar1S0S33P016P063P056P059(0)='1' AND  B(12)='1' AND B( 2)='0' )then
          cVar2S0S33P034P035nsss(0) <='1';
          else
          cVar2S0S33P034P035nsss(0) <='0';
          end if;
        if(cVar1S1S33P016P063P056P059(0)='1' AND  B(12)='1' AND B( 2)='1' AND A(12)='0' )then
          cVar2S1S33P034P035P014nsss(0) <='1';
          else
          cVar2S1S33P034P035P014nsss(0) <='0';
          end if;
        if(cVar1S2S33P016P063P056P059(0)='1' AND  B(12)='0' AND B(11)='1' AND B( 1)='0' )then
          cVar2S2S33N034P036P037nsss(0) <='1';
          else
          cVar2S2S33N034P036P037nsss(0) <='0';
          end if;
        if(cVar1S3S33P016P063P056P059(0)='1' AND  B(12)='0' AND B(11)='0' AND B( 2)='1' )then
          cVar2S3S33N034N036P035nsss(0) <='1';
          else
          cVar2S3S33N034N036P035nsss(0) <='0';
          end if;
        if(cVar1S4S33P016P063P056P059(0)='1' AND  B(13)='0' AND D(11)='0' AND E( 9)='0' )then
          cVar2S4S33P032P057P067nsss(0) <='1';
          else
          cVar2S4S33P032P057P067nsss(0) <='0';
          end if;
        if(cVar1S5S33P016P063P056P062(0)='1' AND  E( 4)='0' )then
          cVar2S5S33P054nsss(0) <='1';
          else
          cVar2S5S33P054nsss(0) <='0';
          end if;
        if(cVar1S6S33P016N063P059P014(0)='1' AND  E( 2)='0' AND A(17)='1' )then
          cVar2S6S33P062P004nsss(0) <='1';
          else
          cVar2S6S33P062P004nsss(0) <='0';
          end if;
        if(cVar1S7S33P016N063P059P014(0)='1' AND  E( 2)='0' AND A(17)='0' AND A( 0)='0' )then
          cVar2S7S33P062N004P019nsss(0) <='1';
          else
          cVar2S7S33P062N004P019nsss(0) <='0';
          end if;
        if(cVar1S8S33P016N063P059P014(0)='1' AND  E( 2)='1' AND A(15)='0' AND B(12)='1' )then
          cVar2S8S33P062P008P034nsss(0) <='1';
          else
          cVar2S8S33P062P008P034nsss(0) <='0';
          end if;
        if(cVar1S9S33P016N063P059N014(0)='1' AND  D( 1)='1' AND A(14)='0' AND A( 1)='0' )then
          cVar2S9S33P064P010P017nsss(0) <='1';
          else
          cVar2S9S33P064P010P017nsss(0) <='0';
          end if;
        if(cVar1S10S33P016N063P059N014(0)='1' AND  D( 1)='0' AND E( 1)='1' AND A( 1)='0' )then
          cVar2S10S33N064P066P017nsss(0) <='1';
          else
          cVar2S10S33N064P066P017nsss(0) <='0';
          end if;
        if(cVar1S11S33P016N063P059N014(0)='1' AND  D( 1)='0' AND E( 1)='0' AND A(19)='1' )then
          cVar2S11S33N064N066P000nsss(0) <='1';
          else
          cVar2S11S33N064N066P000nsss(0) <='0';
          end if;
        if(cVar1S12S33P016N063P059P032(0)='1' AND  A(13)='1' AND A( 2)='0' )then
          cVar2S12S33P012P015nsss(0) <='1';
          else
          cVar2S12S33P012P015nsss(0) <='0';
          end if;
        if(cVar1S13S33P016N063P059P032(0)='1' AND  A(13)='0' AND A(12)='1' AND A( 0)='1' )then
          cVar2S13S33N012P014P019nsss(0) <='1';
          else
          cVar2S13S33N012P014P019nsss(0) <='0';
          end if;
        if(cVar1S14S33P016N063P059N032(0)='1' AND  D( 8)='1' AND D(10)='1' )then
          cVar2S14S33P069P061nsss(0) <='1';
          else
          cVar2S14S33P069P061nsss(0) <='0';
          end if;
        if(cVar1S15S33P016N063P059N032(0)='1' AND  D( 8)='0' AND A( 4)='1' AND A( 0)='0' )then
          cVar2S15S33N069P011P019nsss(0) <='1';
          else
          cVar2S15S33N069P011P019nsss(0) <='0';
          end if;
        if(cVar1S16S33N016P034P040P021(0)='1' AND  A(18)='1' )then
          cVar2S16S33P002nsss(0) <='1';
          else
          cVar2S16S33P002nsss(0) <='0';
          end if;
        if(cVar1S17S33N016P034P040P021(0)='1' AND  A(18)='0' AND A( 8)='1' )then
          cVar2S17S33N002P003nsss(0) <='1';
          else
          cVar2S17S33N002P003nsss(0) <='0';
          end if;
        if(cVar1S18S33N016P034P040P021(0)='1' AND  A(18)='0' AND A( 8)='0' AND A(17)='1' )then
          cVar2S18S33N002N003P004nsss(0) <='1';
          else
          cVar2S18S33N002N003P004nsss(0) <='0';
          end if;
        if(cVar1S19S33N016P034P040N021(0)='1' AND  A(17)='1' )then
          cVar2S19S33P004nsss(0) <='1';
          else
          cVar2S19S33P004nsss(0) <='0';
          end if;
        if(cVar1S20S33N016P034P040N021(0)='1' AND  A(17)='0' AND A( 5)='0' )then
          cVar2S20S33N004P009nsss(0) <='1';
          else
          cVar2S20S33N004P009nsss(0) <='0';
          end if;
        if(cVar1S21S33N016P034N040P044(0)='1' AND  B( 8)='1' )then
          cVar2S21S33P023nsss(0) <='1';
          else
          cVar2S21S33P023nsss(0) <='0';
          end if;
        if(cVar1S22S33N016P034N040P044(0)='1' AND  B( 8)='0' AND A(16)='1' )then
          cVar2S22S33N023P006nsss(0) <='1';
          else
          cVar2S22S33N023P006nsss(0) <='0';
          end if;
        if(cVar1S23S33N016P034N040P044(0)='1' AND  B( 8)='0' AND A(16)='0' AND E( 4)='1' )then
          cVar2S23S33N023N006P054nsss(0) <='1';
          else
          cVar2S23S33N023N006P054nsss(0) <='0';
          end if;
        if(cVar1S24S33N016P034N040N044(0)='1' AND  E( 5)='1' AND A(12)='0' )then
          cVar2S24S33P050P014nsss(0) <='1';
          else
          cVar2S24S33P050P014nsss(0) <='0';
          end if;
        if(cVar1S25S33N016P034N040N044(0)='1' AND  E( 5)='1' AND A(12)='1' AND D( 0)='1' )then
          cVar2S25S33P050P014P068nsss(0) <='1';
          else
          cVar2S25S33P050P014P068nsss(0) <='0';
          end if;
        if(cVar1S26S33N016P034N040N044(0)='1' AND  E( 5)='0' AND D( 9)='0' AND D(15)='1' )then
          cVar2S26S33N050P065P041nsss(0) <='1';
          else
          cVar2S26S33N050P065P041nsss(0) <='0';
          end if;
        if(cVar1S27S33N016P034N040N044(0)='1' AND  E( 5)='0' AND D( 9)='1' AND A( 1)='1' )then
          cVar2S27S33N050P065P017nsss(0) <='1';
          else
          cVar2S27S33N050P065P017nsss(0) <='0';
          end if;
        if(cVar1S28S33N016P034P014P053(0)='1' AND  E( 1)='0' AND D( 3)='0' AND A( 3)='0' )then
          cVar2S28S33P066P056P013nsss(0) <='1';
          else
          cVar2S28S33P066P056P013nsss(0) <='0';
          end if;
        if(cVar1S29S33N016P034P014P053(0)='1' AND  E( 1)='1' AND A(13)='1' )then
          cVar2S29S33P066P012nsss(0) <='1';
          else
          cVar2S29S33P066P012nsss(0) <='0';
          end if;
        if(cVar1S30S33N016P034P014P053(0)='1' AND  E( 1)='1' AND A(13)='0' AND D( 9)='1' )then
          cVar2S30S33P066N012P065nsss(0) <='1';
          else
          cVar2S30S33P066N012P065nsss(0) <='0';
          end if;
        if(cVar1S31S33N016P034N014P017(0)='1' AND  D( 1)='0' AND B( 2)='0' AND E( 1)='0' )then
          cVar2S31S33P064P035P066nsss(0) <='1';
          else
          cVar2S31S33P064P035P066nsss(0) <='0';
          end if;
        if(cVar1S0S34P067P062P008P049(0)='1' AND  B(16)='1' )then
          cVar2S0S34P026nsss(0) <='1';
          else
          cVar2S0S34P026nsss(0) <='0';
          end if;
        if(cVar1S1S34P067P062P008P049(0)='1' AND  B(16)='0' AND B(17)='1' )then
          cVar2S1S34N026P024nsss(0) <='1';
          else
          cVar2S1S34N026P024nsss(0) <='0';
          end if;
        if(cVar1S2S34P067P062P008N049(0)='1' AND  E(13)='1' AND A(11)='0' AND E( 1)='0' )then
          cVar2S2S34P051P016P066nsss(0) <='1';
          else
          cVar2S2S34P051P016P066nsss(0) <='0';
          end if;
        if(cVar1S3S34P067P062P008N049(0)='1' AND  E(13)='1' AND A(11)='1' AND B(16)='0' )then
          cVar2S3S34P051P016P026nsss(0) <='1';
          else
          cVar2S3S34P051P016P026nsss(0) <='0';
          end if;
        if(cVar1S4S34P067P062P008N049(0)='1' AND  E(13)='0' AND B( 6)='1' )then
          cVar2S4S34N051P027nsss(0) <='1';
          else
          cVar2S4S34N051P027nsss(0) <='0';
          end if;
        if(cVar1S5S34P067P062P008N049(0)='1' AND  E(13)='0' AND B( 6)='0' AND D( 9)='0' )then
          cVar2S5S34N051N027P065nsss(0) <='1';
          else
          cVar2S5S34N051N027P065nsss(0) <='0';
          end if;
        if(cVar1S6S34P067P062N008P035(0)='1' AND  E( 3)='1' AND B( 3)='1' AND B(12)='0' )then
          cVar2S6S34P058P033P034nsss(0) <='1';
          else
          cVar2S6S34P058P033P034nsss(0) <='0';
          end if;
        if(cVar1S7S34P067P062N008P035(0)='1' AND  E( 3)='1' AND B( 3)='0' AND A(13)='1' )then
          cVar2S7S34P058N033P012nsss(0) <='1';
          else
          cVar2S7S34P058N033P012nsss(0) <='0';
          end if;
        if(cVar1S8S34P067P062N008P035(0)='1' AND  E( 3)='0' AND D( 2)='0' )then
          cVar2S8S34N058P060nsss(0) <='1';
          else
          cVar2S8S34N058P060nsss(0) <='0';
          end if;
        if(cVar1S9S34P067P062N008P035(0)='1' AND  E( 3)='0' AND D( 2)='1' AND D(11)='1' )then
          cVar2S9S34N058P060P057nsss(0) <='1';
          else
          cVar2S9S34N058P060P057nsss(0) <='0';
          end if;
        if(cVar1S10S34P067P062N008P035(0)='1' AND  E(10)='1' AND A( 1)='1' AND B(12)='0' )then
          cVar2S10S34P063P017P034nsss(0) <='1';
          else
          cVar2S10S34P063P017P034nsss(0) <='0';
          end if;
        if(cVar1S11S34P067P062N008P035(0)='1' AND  E(10)='1' AND A( 1)='0' AND A(10)='1' )then
          cVar2S11S34P063N017P018nsss(0) <='1';
          else
          cVar2S11S34P063N017P018nsss(0) <='0';
          end if;
        if(cVar1S12S34P067P062N008P035(0)='1' AND  E(10)='0' AND B( 1)='1' AND A( 3)='1' )then
          cVar2S12S34N063P037P013nsss(0) <='1';
          else
          cVar2S12S34N063P037P013nsss(0) <='0';
          end if;
        if(cVar1S13S34P067P062N008P035(0)='1' AND  E(10)='0' AND B( 1)='0' AND A( 2)='1' )then
          cVar2S13S34N063N037P015nsss(0) <='1';
          else
          cVar2S13S34N063N037P015nsss(0) <='0';
          end if;
        if(cVar1S14S34P067P062P055P035(0)='1' AND  A(14)='0' AND A( 4)='0' AND B(12)='0' )then
          cVar2S14S34P010P011P034nsss(0) <='1';
          else
          cVar2S14S34P010P011P034nsss(0) <='0';
          end if;
        if(cVar1S15S34P067P062P055P035(0)='1' AND  A(14)='0' AND A( 4)='1' AND D( 2)='1' )then
          cVar2S15S34P010P011P060nsss(0) <='1';
          else
          cVar2S15S34P010P011P060nsss(0) <='0';
          end if;
        if(cVar1S16S34P067P062P055P035(0)='1' AND  A(14)='1' AND A( 1)='1' AND A( 2)='1' )then
          cVar2S16S34P010P017P015nsss(0) <='1';
          else
          cVar2S16S34P010P017P015nsss(0) <='0';
          end if;
        if(cVar1S17S34P067P062P055N035(0)='1' AND  A(11)='1' AND B(12)='1' )then
          cVar2S17S34P016P034nsss(0) <='1';
          else
          cVar2S17S34P016P034nsss(0) <='0';
          end if;
        if(cVar1S18S34P067P062P055N035(0)='1' AND  A(11)='1' AND B(12)='0' AND B(11)='1' )then
          cVar2S18S34P016N034P036nsss(0) <='1';
          else
          cVar2S18S34P016N034P036nsss(0) <='0';
          end if;
        if(cVar1S19S34P067P062P055N035(0)='1' AND  A(11)='0' AND D( 9)='0' AND D( 3)='1' )then
          cVar2S19S34N016P065P056nsss(0) <='1';
          else
          cVar2S19S34N016P065P056nsss(0) <='0';
          end if;
        if(cVar1S21S34P067P010P069P031(0)='1' AND  E( 4)='0' AND D( 4)='1' )then
          cVar2S21S34P054P052nsss(0) <='1';
          else
          cVar2S21S34P054P052nsss(0) <='0';
          end if;
        if(cVar1S22S34P067P010P069P031(0)='1' AND  E( 4)='0' AND D( 4)='0' AND B(15)='0' )then
          cVar2S22S34P054N052P028nsss(0) <='1';
          else
          cVar2S22S34P054N052P028nsss(0) <='0';
          end if;
        if(cVar1S23S34P067P010P069P031(0)='1' AND  E( 4)='1' AND A( 4)='1' )then
          cVar2S23S34P054P011nsss(0) <='1';
          else
          cVar2S23S34P054P011nsss(0) <='0';
          end if;
        if(cVar1S24S34P067P010P069P031(0)='1' AND  E( 3)='0' AND D(11)='1' )then
          cVar2S24S34P058P057nsss(0) <='1';
          else
          cVar2S24S34P058P057nsss(0) <='0';
          end if;
        if(cVar1S26S34P067P010P015P036(0)='1' AND  D( 8)='1' AND A( 1)='0' )then
          cVar2S26S34P069P017nsss(0) <='1';
          else
          cVar2S26S34P069P017nsss(0) <='0';
          end if;
        if(cVar1S27S34P067P010P015P036(0)='1' AND  A(11)='1' )then
          cVar2S27S34P016nsss(0) <='1';
          else
          cVar2S27S34P016nsss(0) <='0';
          end if;
        if(cVar1S29S34P067P010N015N050(0)='1' AND  A( 7)='0' AND D(12)='1' )then
          cVar2S29S34P005P053nsss(0) <='1';
          else
          cVar2S29S34P005P053nsss(0) <='0';
          end if;
        if(cVar1S0S35P058P035P013P066(0)='1' AND  B( 4)='1' )then
          cVar2S0S35P031nsss(0) <='1';
          else
          cVar2S0S35P031nsss(0) <='0';
          end if;
        if(cVar1S1S35P058P035P013P066(0)='1' AND  B( 4)='0' AND B( 3)='1' )then
          cVar2S1S35N031P033nsss(0) <='1';
          else
          cVar2S1S35N031P033nsss(0) <='0';
          end if;
        if(cVar1S2S35P058P035P013P066(0)='1' AND  B( 4)='0' AND B( 3)='0' AND B( 1)='1' )then
          cVar2S2S35N031N033P037nsss(0) <='1';
          else
          cVar2S2S35N031N033P037nsss(0) <='0';
          end if;
        if(cVar1S3S35P058P035P013P066(0)='1' AND  A(13)='0' AND D( 0)='1' )then
          cVar2S3S35P012P068nsss(0) <='1';
          else
          cVar2S3S35P012P068nsss(0) <='0';
          end if;
        if(cVar1S4S35P058P035N013P004(0)='1' AND  B( 4)='0' AND A(12)='1' AND D( 2)='1' )then
          cVar2S4S35P031P014P060nsss(0) <='1';
          else
          cVar2S4S35P031P014P060nsss(0) <='0';
          end if;
        if(cVar1S5S35P058P035N013P004(0)='1' AND  B( 4)='0' AND A(12)='0' AND A( 4)='0' )then
          cVar2S5S35P031N014P011nsss(0) <='1';
          else
          cVar2S5S35P031N014P011nsss(0) <='0';
          end if;
        if(cVar1S6S35P058P035N013P004(0)='1' AND  B( 4)='1' AND A(13)='1' )then
          cVar2S6S35P031P012nsss(0) <='1';
          else
          cVar2S6S35P031P012nsss(0) <='0';
          end if;
        if(cVar1S7S35P058P035P060P034(0)='1' AND  D( 8)='0' AND A( 5)='0' AND A(12)='1' )then
          cVar2S7S35P069P009P014nsss(0) <='1';
          else
          cVar2S7S35P069P009P014nsss(0) <='0';
          end if;
        if(cVar1S8S35N058P030P012P031(0)='1' AND  D( 3)='1' )then
          cVar2S8S35P056nsss(0) <='1';
          else
          cVar2S8S35P056nsss(0) <='0';
          end if;
        if(cVar1S9S35N058P030P012P031(0)='1' AND  D( 3)='0' AND D(11)='1' )then
          cVar2S9S35N056P057nsss(0) <='1';
          else
          cVar2S9S35N056P057nsss(0) <='0';
          end if;
        if(cVar1S10S35N058P030P012P031(0)='1' AND  D( 3)='0' AND D(11)='0' AND E(11)='1' )then
          cVar2S10S35N056N057P059nsss(0) <='1';
          else
          cVar2S10S35N056N057P059nsss(0) <='0';
          end if;
        if(cVar1S11S35N058P030N012P010(0)='1' AND  D(11)='1' )then
          cVar2S11S35P057nsss(0) <='1';
          else
          cVar2S11S35P057nsss(0) <='0';
          end if;
        if(cVar1S12S35N058P030N012P010(0)='1' AND  D(11)='0' AND E( 4)='1' )then
          cVar2S12S35N057P054nsss(0) <='1';
          else
          cVar2S12S35N057P054nsss(0) <='0';
          end if;
        if(cVar1S13S35N058P030N012N010(0)='1' AND  A( 3)='1' AND D(11)='1' )then
          cVar2S13S35P013P057nsss(0) <='1';
          else
          cVar2S13S35P013P057nsss(0) <='0';
          end if;
        if(cVar1S14S35N058N030P024P006(0)='1' AND  E(14)='1' )then
          cVar2S14S35P047nsss(0) <='1';
          else
          cVar2S14S35P047nsss(0) <='0';
          end if;
        if(cVar1S15S35N058N030P024P006(0)='1' AND  E(14)='0' AND E(15)='1' )then
          cVar2S15S35N047P043nsss(0) <='1';
          else
          cVar2S15S35N047P043nsss(0) <='0';
          end if;
        if(cVar1S16S35N058N030P024P006(0)='1' AND  E(14)='0' AND E(15)='0' AND D( 6)='1' )then
          cVar2S16S35N047N043P044nsss(0) <='1';
          else
          cVar2S16S35N047N043P044nsss(0) <='0';
          end if;
        if(cVar1S17S35N058N030P024N006(0)='1' AND  B( 7)='0' AND E(14)='1' AND E( 1)='0' )then
          cVar2S17S35P025P047P066nsss(0) <='1';
          else
          cVar2S17S35P025P047P066nsss(0) <='0';
          end if;
        if(cVar1S18S35N058N030P024N006(0)='1' AND  B( 7)='0' AND E(14)='0' AND D(14)='1' )then
          cVar2S18S35P025N047P045nsss(0) <='1';
          else
          cVar2S18S35P025N047P045nsss(0) <='0';
          end if;
        if(cVar1S19S35N058N030N024P037(0)='1' AND  D(11)='0' AND D( 4)='0' AND E( 4)='0' )then
          cVar2S19S35P057P052P054nsss(0) <='1';
          else
          cVar2S19S35P057P052P054nsss(0) <='0';
          end if;
        if(cVar1S20S35N058N030N024P037(0)='1' AND  D(11)='0' AND D( 4)='1' AND E( 9)='1' )then
          cVar2S20S35P057P052P067nsss(0) <='1';
          else
          cVar2S20S35P057P052P067nsss(0) <='0';
          end if;
        if(cVar1S21S35N058N030N024P037(0)='1' AND  D(11)='1' AND D( 0)='1' AND A(10)='1' )then
          cVar2S21S35P057P068P018nsss(0) <='1';
          else
          cVar2S21S35P057P068P018nsss(0) <='0';
          end if;
        if(cVar1S22S35N058N030N024N037(0)='1' AND  B( 4)='1' AND E( 4)='1' )then
          cVar2S22S35P031P054nsss(0) <='1';
          else
          cVar2S22S35P031P054nsss(0) <='0';
          end if;
        if(cVar1S23S35N058N030N024N037(0)='1' AND  B( 4)='1' AND E( 4)='0' AND A( 3)='1' )then
          cVar2S23S35P031N054P013nsss(0) <='1';
          else
          cVar2S23S35P031N054P013nsss(0) <='0';
          end if;
        if(cVar1S24S35N058N030N024N037(0)='1' AND  B( 4)='0' AND B(15)='1' AND A(14)='1' )then
          cVar2S24S35N031P028P010nsss(0) <='1';
          else
          cVar2S24S35N031P028P010nsss(0) <='0';
          end if;
        if(cVar1S25S35N058N030N024N037(0)='1' AND  B( 4)='0' AND B(15)='0' AND B( 5)='1' )then
          cVar2S25S35N031N028P029nsss(0) <='1';
          else
          cVar2S25S35N031N028P029nsss(0) <='0';
          end if;
        if(cVar1S1S36P037P048N025P009(0)='1' AND  B( 6)='1' )then
          cVar2S1S36P027nsss(0) <='1';
          else
          cVar2S1S36P027nsss(0) <='0';
          end if;
        if(cVar1S2S36P037P048N025P009(0)='1' AND  B( 6)='0' AND A( 3)='0' )then
          cVar2S2S36N027P013nsss(0) <='1';
          else
          cVar2S2S36N027P013nsss(0) <='0';
          end if;
        if(cVar1S3S36P037P048N025N009(0)='1' AND  B(17)='1' AND A(12)='0' )then
          cVar2S3S36P024P014nsss(0) <='1';
          else
          cVar2S3S36P024P014nsss(0) <='0';
          end if;
        if(cVar1S4S36P037P048N025N009(0)='1' AND  B(17)='0' AND D( 4)='0' AND B(14)='1' )then
          cVar2S4S36N024P052P030nsss(0) <='1';
          else
          cVar2S4S36N024P052P030nsss(0) <='0';
          end if;
        if(cVar1S5S36P037N048P046P009(0)='1' AND  B( 6)='0' AND E( 5)='0' )then
          cVar2S5S36P027P050nsss(0) <='1';
          else
          cVar2S5S36P027P050nsss(0) <='0';
          end if;
        if(cVar1S6S36P037N048P046P009(0)='1' AND  B( 6)='1' AND A( 6)='1' )then
          cVar2S6S36P027P007nsss(0) <='1';
          else
          cVar2S6S36P027P007nsss(0) <='0';
          end if;
        if(cVar1S7S36P037N048P046P009(0)='1' AND  B( 6)='1' AND A( 6)='0' AND E( 5)='1' )then
          cVar2S7S36P027N007P050nsss(0) <='1';
          else
          cVar2S7S36P027N007P050nsss(0) <='0';
          end if;
        if(cVar1S8S36P037N048P046P009(0)='1' AND  D(13)='1' AND A( 1)='0' )then
          cVar2S8S36P049P017nsss(0) <='1';
          else
          cVar2S8S36P049P017nsss(0) <='0';
          end if;
        if(cVar1S9S36P037N048P046P009(0)='1' AND  D(13)='0' AND D( 4)='1' AND A( 3)='0' )then
          cVar2S9S36N049P052P013nsss(0) <='1';
          else
          cVar2S9S36N049P052P013nsss(0) <='0';
          end if;
        if(cVar1S10S36P037N048P046P009(0)='1' AND  D(13)='0' AND D( 4)='0' AND A( 6)='1' )then
          cVar2S10S36N049N052P007nsss(0) <='1';
          else
          cVar2S10S36N049N052P007nsss(0) <='0';
          end if;
        if(cVar1S11S36P037N048P046P044(0)='1' AND  B( 7)='1' AND A( 6)='1' )then
          cVar2S11S36P025P007nsss(0) <='1';
          else
          cVar2S11S36P025P007nsss(0) <='0';
          end if;
        if(cVar1S12S36P037N048P046P044(0)='1' AND  B( 7)='1' AND A( 6)='0' AND A(16)='1' )then
          cVar2S12S36P025N007P006nsss(0) <='1';
          else
          cVar2S12S36P025N007P006nsss(0) <='0';
          end if;
        if(cVar1S13S36P037N048P046P044(0)='1' AND  B( 7)='0' AND A(17)='1' )then
          cVar2S13S36N025P004nsss(0) <='1';
          else
          cVar2S13S36N025P004nsss(0) <='0';
          end if;
        if(cVar1S14S36P037N048P046P044(0)='1' AND  B( 7)='0' AND A(17)='0' AND A(10)='1' )then
          cVar2S14S36N025N004P018nsss(0) <='1';
          else
          cVar2S14S36N025N004P018nsss(0) <='0';
          end if;
        if(cVar1S15S36P037N048P046N044(0)='1' AND  A( 0)='0' AND A( 1)='1' )then
          cVar2S15S36P019P017nsss(0) <='1';
          else
          cVar2S15S36P019P017nsss(0) <='0';
          end if;
        if(cVar1S16S36P037P059P005P035(0)='1' AND  A(12)='1' )then
          cVar2S16S36P014nsss(0) <='1';
          else
          cVar2S16S36P014nsss(0) <='0';
          end if;
        if(cVar1S17S36P037P059P005P035(0)='1' AND  A(12)='0' AND E( 9)='0' AND B(17)='1' )then
          cVar2S17S36N014P067P024nsss(0) <='1';
          else
          cVar2S17S36N014P067P024nsss(0) <='0';
          end if;
        if(cVar1S18S36P037P059P005N035(0)='1' AND  B(11)='0' AND B( 7)='1' AND E( 6)='1' )then
          cVar2S18S36P036P025P046nsss(0) <='1';
          else
          cVar2S18S36P036P025P046nsss(0) <='0';
          end if;
        if(cVar1S19S36P037P059P005N035(0)='1' AND  B(11)='1' AND A(12)='1' AND D( 8)='0' )then
          cVar2S19S36P036P014P069nsss(0) <='1';
          else
          cVar2S19S36P036P014P069nsss(0) <='0';
          end if;
        if(cVar1S20S36P037P059P005N035(0)='1' AND  B(11)='1' AND A(12)='0' AND A( 3)='1' )then
          cVar2S20S36P036N014P013nsss(0) <='1';
          else
          cVar2S20S36P036N014P013nsss(0) <='0';
          end if;
        if(cVar1S21S36P037P059P005P063(0)='1' AND  B( 3)='0' AND A( 8)='0' AND A(14)='1' )then
          cVar2S21S36P033P003P010nsss(0) <='1';
          else
          cVar2S21S36P033P003P010nsss(0) <='0';
          end if;
        if(cVar1S23S36P037P059N008P060(0)='1' AND  E( 2)='1' )then
          cVar2S23S36P062nsss(0) <='1';
          else
          cVar2S23S36P062nsss(0) <='0';
          end if;
        if(cVar1S24S36P037P059N008N060(0)='1' AND  A(12)='1' AND D( 0)='0' AND D( 1)='1' )then
          cVar2S24S36P014P068P064nsss(0) <='1';
          else
          cVar2S24S36P014P068P064nsss(0) <='0';
          end if;
        if(cVar1S2S37P048P025N007N004(0)='1' AND  A(16)='1' )then
          cVar2S2S37P006nsss(0) <='1';
          else
          cVar2S2S37P006nsss(0) <='0';
          end if;
        if(cVar1S3S37P048P025N007N004(0)='1' AND  A(16)='0' AND A( 5)='1' )then
          cVar2S3S37N006P009nsss(0) <='1';
          else
          cVar2S3S37N006P009nsss(0) <='0';
          end if;
        if(cVar1S4S37P048P025N007N004(0)='1' AND  A(16)='0' AND A( 5)='0' AND A( 7)='1' )then
          cVar2S4S37N006N009P005nsss(0) <='1';
          else
          cVar2S4S37N006N009P005nsss(0) <='0';
          end if;
        if(cVar1S6S37P048N025P037P017(0)='1' AND  D( 2)='1' )then
          cVar2S6S37P060nsss(0) <='1';
          else
          cVar2S6S37P060nsss(0) <='0';
          end if;
        if(cVar1S7S37P048N025P037P017(0)='1' AND  D( 2)='0' AND A( 6)='1' )then
          cVar2S7S37N060P007nsss(0) <='1';
          else
          cVar2S7S37N060P007nsss(0) <='0';
          end if;
        if(cVar1S8S37P048N025P037P017(0)='1' AND  D( 2)='0' AND A( 6)='0' AND A(15)='1' )then
          cVar2S8S37N060N007P008nsss(0) <='1';
          else
          cVar2S8S37N060N007P008nsss(0) <='0';
          end if;
        if(cVar1S10S37P048N025P037N006(0)='1' AND  B(11)='0' AND E( 2)='1' )then
          cVar2S10S37P036P062nsss(0) <='1';
          else
          cVar2S10S37P036P062nsss(0) <='0';
          end if;
        if(cVar1S12S37N048P044N004P005(0)='1' AND  B( 8)='1' )then
          cVar2S12S37P023nsss(0) <='1';
          else
          cVar2S12S37P023nsss(0) <='0';
          end if;
        if(cVar1S13S37N048P044N004P005(0)='1' AND  B( 8)='0' AND E( 6)='1' )then
          cVar2S13S37N023P046nsss(0) <='1';
          else
          cVar2S13S37N023P046nsss(0) <='0';
          end if;
        if(cVar1S14S37N048P044N004N005(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S14S37P006P024nsss(0) <='1';
          else
          cVar2S14S37P006P024nsss(0) <='0';
          end if;
        if(cVar1S15S37N048P044N004N005(0)='1' AND  A(16)='1' AND B(17)='0' AND B( 7)='1' )then
          cVar2S15S37P006N024P025nsss(0) <='1';
          else
          cVar2S15S37P006N024P025nsss(0) <='0';
          end if;
        if(cVar1S16S37N048P044N004N005(0)='1' AND  A(16)='0' AND B( 9)='1' )then
          cVar2S16S37N006P021nsss(0) <='1';
          else
          cVar2S16S37N006P021nsss(0) <='0';
          end if;
        if(cVar1S17S37N048P044N004N005(0)='1' AND  A(16)='0' AND B( 9)='0' AND A( 6)='1' )then
          cVar2S17S37N006N021P007nsss(0) <='1';
          else
          cVar2S17S37N006N021P007nsss(0) <='0';
          end if;
        if(cVar1S18S37N048N044P046P025(0)='1' AND  B(16)='1' AND D(13)='1' )then
          cVar2S18S37P026P049nsss(0) <='1';
          else
          cVar2S18S37P026P049nsss(0) <='0';
          end if;
        if(cVar1S19S37N048N044P046P025(0)='1' AND  B(16)='1' AND D(13)='0' AND E(12)='0' )then
          cVar2S19S37P026N049P055nsss(0) <='1';
          else
          cVar2S19S37P026N049P055nsss(0) <='0';
          end if;
        if(cVar1S20S37N048N044P046P025(0)='1' AND  B(16)='0' AND B(17)='1' AND E(14)='1' )then
          cVar2S20S37N026P024P047nsss(0) <='1';
          else
          cVar2S20S37N026P024P047nsss(0) <='0';
          end if;
        if(cVar1S21S37N048N044P046P025(0)='1' AND  A( 6)='1' AND E(14)='1' )then
          cVar2S21S37P007P047nsss(0) <='1';
          else
          cVar2S21S37P007P047nsss(0) <='0';
          end if;
        if(cVar1S22S37N048N044P046P025(0)='1' AND  A( 6)='1' AND E(14)='0' AND E(15)='1' )then
          cVar2S22S37P007N047P043nsss(0) <='1';
          else
          cVar2S22S37P007N047P043nsss(0) <='0';
          end if;
        if(cVar1S23S37N048N044P046P025(0)='1' AND  A( 6)='0' AND A( 5)='1' )then
          cVar2S23S37N007P009nsss(0) <='1';
          else
          cVar2S23S37N007P009nsss(0) <='0';
          end if;
        if(cVar1S24S37N048N044P046P027(0)='1' AND  E( 4)='1' )then
          cVar2S24S37P054nsss(0) <='1';
          else
          cVar2S24S37P054nsss(0) <='0';
          end if;
        if(cVar1S2S38P048P025N007N004(0)='1' AND  A( 5)='1' )then
          cVar2S2S38P009nsss(0) <='1';
          else
          cVar2S2S38P009nsss(0) <='0';
          end if;
        if(cVar1S3S38P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S3S38N009P006nsss(0) <='1';
          else
          cVar2S3S38N009P006nsss(0) <='0';
          end if;
        if(cVar1S4S38P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S4S38N009N006P005nsss(0) <='1';
          else
          cVar2S4S38N009N006P005nsss(0) <='0';
          end if;
        if(cVar1S5S38P048N025P052P027(0)='1' AND  A( 6)='1' )then
          cVar2S5S38P007nsss(0) <='1';
          else
          cVar2S5S38P007nsss(0) <='0';
          end if;
        if(cVar1S6S38P048N025P052P027(0)='1' AND  A( 6)='0' AND A(16)='1' )then
          cVar2S6S38N007P006nsss(0) <='1';
          else
          cVar2S6S38N007P006nsss(0) <='0';
          end if;
        if(cVar1S7S38P048N025P052P027(0)='1' AND  A( 6)='0' AND A(16)='0' AND A( 5)='1' )then
          cVar2S7S38N007N006P009nsss(0) <='1';
          else
          cVar2S7S38N007N006P009nsss(0) <='0';
          end if;
        if(cVar1S8S38P048N025P052N027(0)='1' AND  B( 1)='0' AND B(14)='1' )then
          cVar2S8S38P037P030nsss(0) <='1';
          else
          cVar2S8S38P037P030nsss(0) <='0';
          end if;
        if(cVar1S9S38P048N025P052N027(0)='1' AND  B( 1)='0' AND B(14)='0' AND A(19)='0' )then
          cVar2S9S38P037N030P000nsss(0) <='1';
          else
          cVar2S9S38P037N030P000nsss(0) <='0';
          end if;
        if(cVar1S10S38P048N025P052N027(0)='1' AND  B( 1)='1' AND A(16)='1' )then
          cVar2S10S38P037P006nsss(0) <='1';
          else
          cVar2S10S38P037P006nsss(0) <='0';
          end if;
        if(cVar1S12S38P048N025P052N046(0)='1' AND  A( 5)='1' )then
          cVar2S12S38P009nsss(0) <='1';
          else
          cVar2S12S38P009nsss(0) <='0';
          end if;
        if(cVar1S13S38N048P025P046P018(0)='1' AND  D(14)='0' AND E(15)='0' )then
          cVar2S13S38P045P043nsss(0) <='1';
          else
          cVar2S13S38P045P043nsss(0) <='0';
          end if;
        if(cVar1S14S38N048P025P046P018(0)='1' AND  D(14)='1' AND B(18)='1' )then
          cVar2S14S38P045P022nsss(0) <='1';
          else
          cVar2S14S38P045P022nsss(0) <='0';
          end if;
        if(cVar1S15S38N048P025P046P018(0)='1' AND  D(14)='1' AND B(18)='0' AND B(17)='1' )then
          cVar2S15S38P045N022P024nsss(0) <='1';
          else
          cVar2S15S38P045N022P024nsss(0) <='0';
          end if;
        if(cVar1S16S38N048P025P046N018(0)='1' AND  A(11)='1' AND D( 9)='1' AND E( 4)='0' )then
          cVar2S16S38P016P065P054nsss(0) <='1';
          else
          cVar2S16S38P016P065P054nsss(0) <='0';
          end if;
        if(cVar1S17S38N048P025P046N018(0)='1' AND  A(11)='1' AND D( 9)='0' AND B( 4)='0' )then
          cVar2S17S38P016N065P031nsss(0) <='1';
          else
          cVar2S17S38P016N065P031nsss(0) <='0';
          end if;
        if(cVar1S18S38N048P025P046N018(0)='1' AND  A(11)='0' AND B(11)='0' )then
          cVar2S18S38N016P036nsss(0) <='1';
          else
          cVar2S18S38N016P036nsss(0) <='0';
          end if;
        if(cVar1S19S38N048P025P046N018(0)='1' AND  A(11)='0' AND B(11)='1' AND A( 1)='1' )then
          cVar2S19S38N016P036P017nsss(0) <='1';
          else
          cVar2S19S38N016P036P017nsss(0) <='0';
          end if;
        if(cVar1S20S38N048P025P046P027(0)='1' AND  A(10)='1' AND A( 0)='0' )then
          cVar2S20S38P018P019nsss(0) <='1';
          else
          cVar2S20S38P018P019nsss(0) <='0';
          end if;
        if(cVar1S21S38N048P025P046P027(0)='1' AND  A(10)='0' AND D( 3)='1' )then
          cVar2S21S38N018P056nsss(0) <='1';
          else
          cVar2S21S38N018P056nsss(0) <='0';
          end if;
        if(cVar1S22S38N048P025P046P027(0)='1' AND  A(10)='0' AND D( 3)='0' AND A(17)='1' )then
          cVar2S22S38N018N056P004nsss(0) <='1';
          else
          cVar2S22S38N018N056P004nsss(0) <='0';
          end if;
        if(cVar1S23S38N048P025P007P009(0)='1' AND  D( 6)='1' )then
          cVar2S23S38P044nsss(0) <='1';
          else
          cVar2S23S38P044nsss(0) <='0';
          end if;
        if(cVar1S24S38N048P025P007P009(0)='1' AND  D( 6)='0' AND E(15)='1' )then
          cVar2S24S38N044P043nsss(0) <='1';
          else
          cVar2S24S38N044P043nsss(0) <='0';
          end if;
        if(cVar1S25S38N048P025P007P009(0)='1' AND  D( 6)='0' AND E(15)='0' AND D(13)='1' )then
          cVar2S25S38N044N043P049nsss(0) <='1';
          else
          cVar2S25S38N044N043P049nsss(0) <='0';
          end if;
        if(cVar1S26S38N048P025N007P044(0)='1' AND  A(16)='1' )then
          cVar2S26S38P006nsss(0) <='1';
          else
          cVar2S26S38P006nsss(0) <='0';
          end if;
        if(cVar1S27S38N048P025N007N044(0)='1' AND  A( 5)='1' )then
          cVar2S27S38P009nsss(0) <='1';
          else
          cVar2S27S38P009nsss(0) <='0';
          end if;
        if(cVar1S2S39P048P025N007N004(0)='1' AND  A( 5)='1' )then
          cVar2S2S39P009nsss(0) <='1';
          else
          cVar2S2S39P009nsss(0) <='0';
          end if;
        if(cVar1S3S39P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S3S39N009P006nsss(0) <='1';
          else
          cVar2S3S39N009P006nsss(0) <='0';
          end if;
        if(cVar1S4S39P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S4S39N009N006P005nsss(0) <='1';
          else
          cVar2S4S39N009N006P005nsss(0) <='0';
          end if;
        if(cVar1S6S39P048N025P027N007(0)='1' AND  A(16)='1' )then
          cVar2S6S39P006nsss(0) <='1';
          else
          cVar2S6S39P006nsss(0) <='0';
          end if;
        if(cVar1S7S39P048N025P027N007(0)='1' AND  A(16)='0' AND A( 5)='1' AND E( 5)='1' )then
          cVar2S7S39N006P009P050nsss(0) <='1';
          else
          cVar2S7S39N006P009P050nsss(0) <='0';
          end if;
        if(cVar1S8S39P048N025P027N007(0)='1' AND  A(16)='0' AND A( 5)='0' AND A(15)='1' )then
          cVar2S8S39N006N009P008nsss(0) <='1';
          else
          cVar2S8S39N006N009P008nsss(0) <='0';
          end if;
        if(cVar1S10S39P048N025N027N058(0)='1' AND  B(14)='1' )then
          cVar2S10S39P030nsss(0) <='1';
          else
          cVar2S10S39P030nsss(0) <='0';
          end if;
        if(cVar1S11S39P048N025N027N058(0)='1' AND  B(14)='0' AND B(17)='1' AND A( 3)='0' )then
          cVar2S11S39N030P024P013nsss(0) <='1';
          else
          cVar2S11S39N030P024P013nsss(0) <='0';
          end if;
        if(cVar1S12S39P048N025N027N058(0)='1' AND  B(14)='0' AND B(17)='0' AND D(14)='1' )then
          cVar2S12S39N030N024P045nsss(0) <='1';
          else
          cVar2S12S39N030N024P045nsss(0) <='0';
          end if;
        if(cVar1S14S39N048P044N004P005(0)='1' AND  B( 8)='1' )then
          cVar2S14S39P023nsss(0) <='1';
          else
          cVar2S14S39P023nsss(0) <='0';
          end if;
        if(cVar1S15S39N048P044N004P005(0)='1' AND  B( 8)='0' AND E( 6)='1' )then
          cVar2S15S39N023P046nsss(0) <='1';
          else
          cVar2S15S39N023P046nsss(0) <='0';
          end if;
        if(cVar1S16S39N048P044N004N005(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S16S39P006P024nsss(0) <='1';
          else
          cVar2S16S39P006P024nsss(0) <='0';
          end if;
        if(cVar1S17S39N048P044N004N005(0)='1' AND  A(16)='1' AND B(17)='0' AND B( 7)='1' )then
          cVar2S17S39P006N024P025nsss(0) <='1';
          else
          cVar2S17S39P006N024P025nsss(0) <='0';
          end if;
        if(cVar1S18S39N048P044N004N005(0)='1' AND  A(16)='0' AND B( 9)='1' )then
          cVar2S18S39N006P021nsss(0) <='1';
          else
          cVar2S18S39N006P021nsss(0) <='0';
          end if;
        if(cVar1S19S39N048P044N004N005(0)='1' AND  A(16)='0' AND B( 9)='0' AND E( 7)='0' )then
          cVar2S19S39N006N021P042nsss(0) <='1';
          else
          cVar2S19S39N006N021P042nsss(0) <='0';
          end if;
        if(cVar1S20S39N048N044P046P052(0)='1' AND  E( 9)='1' AND A( 2)='1' )then
          cVar2S20S39P067P015nsss(0) <='1';
          else
          cVar2S20S39P067P015nsss(0) <='0';
          end if;
        if(cVar1S21S39N048N044P046P052(0)='1' AND  E( 9)='1' AND A( 2)='0' AND B( 5)='0' )then
          cVar2S21S39P067N015P029nsss(0) <='1';
          else
          cVar2S21S39P067N015P029nsss(0) <='0';
          end if;
        if(cVar1S22S39N048N044P046P052(0)='1' AND  E( 9)='0' AND D( 9)='1' )then
          cVar2S22S39N067P065nsss(0) <='1';
          else
          cVar2S22S39N067P065nsss(0) <='0';
          end if;
        if(cVar1S23S39N048N044P046P052(0)='1' AND  E( 9)='0' AND D( 9)='0' AND B(12)='0' )then
          cVar2S23S39N067N065P034nsss(0) <='1';
          else
          cVar2S23S39N067N065P034nsss(0) <='0';
          end if;
        if(cVar1S24S39N048N044P046N052(0)='1' AND  A(10)='1' AND A(11)='0' AND B(12)='0' )then
          cVar2S24S39P018P016P034nsss(0) <='1';
          else
          cVar2S24S39P018P016P034nsss(0) <='0';
          end if;
        if(cVar1S25S39N048N044P046N052(0)='1' AND  A(10)='1' AND A(11)='1' AND E(10)='1' )then
          cVar2S25S39P018P016P063nsss(0) <='1';
          else
          cVar2S25S39P018P016P063nsss(0) <='0';
          end if;
        if(cVar1S26S39N048N044P046N052(0)='1' AND  A(10)='0' AND A(11)='1' AND D( 9)='1' )then
          cVar2S26S39N018P016P065nsss(0) <='1';
          else
          cVar2S26S39N018P016P065nsss(0) <='0';
          end if;
        if(cVar1S27S39N048N044P046P027(0)='1' AND  A( 0)='0' AND A(10)='1' )then
          cVar2S27S39P019P018nsss(0) <='1';
          else
          cVar2S27S39P019P018nsss(0) <='0';
          end if;
        if(cVar1S28S39N048N044P046P027(0)='1' AND  A( 0)='0' AND A(10)='0' AND A( 3)='1' )then
          cVar2S28S39P019N018P013nsss(0) <='1';
          else
          cVar2S28S39P019N018P013nsss(0) <='0';
          end if;
        if(cVar1S1S40P018P048N025P027(0)='1' AND  A( 5)='1' )then
          cVar2S1S40P009nsss(0) <='1';
          else
          cVar2S1S40P009nsss(0) <='0';
          end if;
        if(cVar1S2S40P018P048N025P027(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S2S40N009P006nsss(0) <='1';
          else
          cVar2S2S40N009P006nsss(0) <='0';
          end if;
        if(cVar1S3S40P018P048N025P027(0)='1' AND  A( 5)='0' AND A(16)='0' AND A( 6)='1' )then
          cVar2S3S40N009N006P007nsss(0) <='1';
          else
          cVar2S3S40N009N006P007nsss(0) <='0';
          end if;
        if(cVar1S4S40P018P048N025N027(0)='1' AND  E( 3)='1' )then
          cVar2S4S40P058nsss(0) <='1';
          else
          cVar2S4S40P058nsss(0) <='0';
          end if;
        if(cVar1S5S40P018P048N025N027(0)='1' AND  E( 3)='0' AND B(17)='1' AND E( 6)='1' )then
          cVar2S5S40N058P024P046nsss(0) <='1';
          else
          cVar2S5S40N058P024P046nsss(0) <='0';
          end if;
        if(cVar1S6S40P018N048P010P032(0)='1' AND  E(11)='1' AND A( 0)='0' AND E( 3)='0' )then
          cVar2S6S40P059P019P058nsss(0) <='1';
          else
          cVar2S6S40P059P019P058nsss(0) <='0';
          end if;
        if(cVar1S7S40P018N048P010P032(0)='1' AND  E(11)='1' AND A( 0)='1' AND E( 1)='0' )then
          cVar2S7S40P059P019P066nsss(0) <='1';
          else
          cVar2S7S40P059P019P066nsss(0) <='0';
          end if;
        if(cVar1S8S40P018N048P010P032(0)='1' AND  E(11)='0' AND D( 2)='1' )then
          cVar2S8S40N059P060nsss(0) <='1';
          else
          cVar2S8S40N059P060nsss(0) <='0';
          end if;
        if(cVar1S9S40P018N048P010P032(0)='1' AND  E(11)='0' AND D( 2)='0' AND A( 2)='1' )then
          cVar2S9S40N059N060P015nsss(0) <='1';
          else
          cVar2S9S40N059N060P015nsss(0) <='0';
          end if;
        if(cVar1S10S40P018N048P010N032(0)='1' AND  B( 2)='1' AND B(12)='0' AND D(11)='0' )then
          cVar2S10S40P035P034P057nsss(0) <='1';
          else
          cVar2S10S40P035P034P057nsss(0) <='0';
          end if;
        if(cVar1S11S40P018N048P010N032(0)='1' AND  B( 2)='1' AND B(12)='1' AND A( 5)='1' )then
          cVar2S11S40P035P034P009nsss(0) <='1';
          else
          cVar2S11S40P035P034P009nsss(0) <='0';
          end if;
        if(cVar1S12S40P018N048P010N032(0)='1' AND  B( 2)='0' AND A( 4)='1' )then
          cVar2S12S40N035P011nsss(0) <='1';
          else
          cVar2S12S40N035P011nsss(0) <='0';
          end if;
        if(cVar1S13S40P018N048P010N032(0)='1' AND  B( 2)='0' AND A( 4)='0' AND B( 5)='0' )then
          cVar2S13S40N035N011P029nsss(0) <='1';
          else
          cVar2S13S40N035N011P029nsss(0) <='0';
          end if;
        if(cVar1S14S40P018N048P010P028(0)='1' AND  E(12)='1' )then
          cVar2S14S40P055nsss(0) <='1';
          else
          cVar2S14S40P055nsss(0) <='0';
          end if;
        if(cVar1S15S40P018N048P010P028(0)='1' AND  E(12)='0' AND E( 4)='1' )then
          cVar2S15S40N055P054nsss(0) <='1';
          else
          cVar2S15S40N055P054nsss(0) <='0';
          end if;
        if(cVar1S16S40P018N048P010P028(0)='1' AND  E(12)='0' AND E( 4)='0' AND E(13)='1' )then
          cVar2S16S40N055N054P051nsss(0) <='1';
          else
          cVar2S16S40N055N054P051nsss(0) <='0';
          end if;
        if(cVar1S17S40P018N048P010N028(0)='1' AND  B(14)='1' AND D(11)='1' )then
          cVar2S17S40P030P057nsss(0) <='1';
          else
          cVar2S17S40P030P057nsss(0) <='0';
          end if;
        if(cVar1S18S40P018N048P010N028(0)='1' AND  B(14)='1' AND D(11)='0' AND D( 3)='1' )then
          cVar2S18S40P030N057P056nsss(0) <='1';
          else
          cVar2S18S40P030N057P056nsss(0) <='0';
          end if;
        if(cVar1S19S40P018N048P010N028(0)='1' AND  B(14)='0' AND B( 5)='1' AND B( 1)='0' )then
          cVar2S19S40N030P029P037nsss(0) <='1';
          else
          cVar2S19S40N030P029P037nsss(0) <='0';
          end if;
        if(cVar1S20S40P018P069P009P068(0)='1' AND  B(15)='0' AND D(11)='0' AND A(19)='0' )then
          cVar2S20S40P028P057P000nsss(0) <='1';
          else
          cVar2S20S40P028P057P000nsss(0) <='0';
          end if;
        if(cVar1S21S40P018P069P009P068(0)='1' AND  A( 6)='1' )then
          cVar2S21S40P007nsss(0) <='1';
          else
          cVar2S21S40P007nsss(0) <='0';
          end if;
        if(cVar1S22S40P018P069P009P068(0)='1' AND  A( 6)='0' AND A( 1)='0' AND B( 1)='0' )then
          cVar2S22S40N007P017P037nsss(0) <='1';
          else
          cVar2S22S40N007P017P037nsss(0) <='0';
          end if;
        if(cVar1S23S40P018P069N009P003(0)='1' AND  E( 1)='0' AND D( 1)='0' )then
          cVar2S23S40P066P064nsss(0) <='1';
          else
          cVar2S23S40P066P064nsss(0) <='0';
          end if;
        if(cVar1S24S40P018P069N009P003(0)='1' AND  E( 1)='1' AND A(11)='0' AND A( 1)='0' )then
          cVar2S24S40P066P016P017nsss(0) <='1';
          else
          cVar2S24S40P066P016P017nsss(0) <='0';
          end if;
        if(cVar1S25S40P018P069N009N003(0)='1' AND  A( 2)='0' AND A( 0)='0' AND E( 1)='1' )then
          cVar2S25S40P015P019P066nsss(0) <='1';
          else
          cVar2S25S40P015P019P066nsss(0) <='0';
          end if;
        if(cVar1S26S40P018P069N009N003(0)='1' AND  A( 2)='0' AND A( 0)='1' AND A( 6)='1' )then
          cVar2S26S40P015P019P007nsss(0) <='1';
          else
          cVar2S26S40P015P019P007nsss(0) <='0';
          end if;
        if(cVar1S27S40P018P069N009N003(0)='1' AND  A( 2)='1' AND A(13)='1' )then
          cVar2S27S40P015P012nsss(0) <='1';
          else
          cVar2S27S40P015P012nsss(0) <='0';
          end if;
        if(cVar1S28S40P018P069N009N003(0)='1' AND  A( 2)='1' AND A(13)='0' AND D( 1)='1' )then
          cVar2S28S40P015N012P064nsss(0) <='1';
          else
          cVar2S28S40P015N012P064nsss(0) <='0';
          end if;
        if(cVar1S2S41P048P025N007N004(0)='1' AND  A( 5)='1' )then
          cVar2S2S41P009nsss(0) <='1';
          else
          cVar2S2S41P009nsss(0) <='0';
          end if;
        if(cVar1S3S41P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S3S41N009P006nsss(0) <='1';
          else
          cVar2S3S41N009P006nsss(0) <='0';
          end if;
        if(cVar1S4S41P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S4S41N009N006P005nsss(0) <='1';
          else
          cVar2S4S41N009N006P005nsss(0) <='0';
          end if;
        if(cVar1S5S41P048N025P052P065(0)='1' AND  E( 5)='1' AND B( 6)='1' )then
          cVar2S5S41P050P027nsss(0) <='1';
          else
          cVar2S5S41P050P027nsss(0) <='0';
          end if;
        if(cVar1S6S41P048N025P052P065(0)='1' AND  E( 5)='1' AND B( 6)='0' AND A( 4)='0' )then
          cVar2S6S41P050N027P011nsss(0) <='1';
          else
          cVar2S6S41P050N027P011nsss(0) <='0';
          end if;
        if(cVar1S7S41P048N025P052P065(0)='1' AND  E( 5)='0' AND A( 7)='0' AND A( 1)='0' )then
          cVar2S7S41N050P005P017nsss(0) <='1';
          else
          cVar2S7S41N050P005P017nsss(0) <='0';
          end if;
        if(cVar1S8S41P048N025P052P065(0)='1' AND  E( 6)='1' )then
          cVar2S8S41P046nsss(0) <='1';
          else
          cVar2S8S41P046nsss(0) <='0';
          end if;
        if(cVar1S10S41P048N025P052N015(0)='1' AND  E( 4)='1' )then
          cVar2S10S41P054nsss(0) <='1';
          else
          cVar2S10S41P054nsss(0) <='0';
          end if;
        if(cVar1S11S41P048N025P052N015(0)='1' AND  E( 4)='0' AND E( 6)='1' )then
          cVar2S11S41N054P046nsss(0) <='1';
          else
          cVar2S11S41N054P046nsss(0) <='0';
          end if;
        if(cVar1S12S41N048P018P059P045(0)='1' AND  E(15)='0' AND B( 7)='0' AND B(18)='0' )then
          cVar2S12S41P043P025P022nsss(0) <='1';
          else
          cVar2S12S41P043P025P022nsss(0) <='0';
          end if;
        if(cVar1S13S41N048P018P059P045(0)='1' AND  E(15)='0' AND B( 7)='1' AND A( 1)='1' )then
          cVar2S13S41P043P025P017nsss(0) <='1';
          else
          cVar2S13S41P043P025P017nsss(0) <='0';
          end if;
        if(cVar1S14S41N048P018P059P045(0)='1' AND  E(15)='1' AND A( 0)='0' AND D(15)='1' )then
          cVar2S14S41P043P019P041nsss(0) <='1';
          else
          cVar2S14S41P043P019P041nsss(0) <='0';
          end if;
        if(cVar1S15S41N048P018P059P045(0)='1' AND  B(18)='1' )then
          cVar2S15S41P022nsss(0) <='1';
          else
          cVar2S15S41P022nsss(0) <='0';
          end if;
        if(cVar1S16S41N048P018P059P045(0)='1' AND  B(18)='0' AND A( 6)='1' )then
          cVar2S16S41N022P007nsss(0) <='1';
          else
          cVar2S16S41N022P007nsss(0) <='0';
          end if;
        if(cVar1S17S41N048P018P059P045(0)='1' AND  B(18)='0' AND A( 6)='0' AND A( 7)='1' )then
          cVar2S17S41N022N007P005nsss(0) <='1';
          else
          cVar2S17S41N022N007P005nsss(0) <='0';
          end if;
        if(cVar1S19S41N048P018P059N050(0)='1' AND  A(17)='0' AND D(10)='1' AND A( 5)='1' )then
          cVar2S19S41P004P061P009nsss(0) <='1';
          else
          cVar2S19S41P004P061P009nsss(0) <='0';
          end if;
        if(cVar1S20S41N048P018P059N050(0)='1' AND  A(17)='0' AND D(10)='0' AND D(11)='1' )then
          cVar2S20S41P004N061P057nsss(0) <='1';
          else
          cVar2S20S41P004N061P057nsss(0) <='0';
          end if;
        if(cVar1S21S41N048N018P032P028(0)='1' AND  D( 9)='0' AND A(12)='1' )then
          cVar2S21S41P065P014nsss(0) <='1';
          else
          cVar2S21S41P065P014nsss(0) <='0';
          end if;
        if(cVar1S22S41N048N018P032P028(0)='1' AND  D( 9)='0' AND A(12)='0' AND A(13)='1' )then
          cVar2S22S41P065N014P012nsss(0) <='1';
          else
          cVar2S22S41P065N014P012nsss(0) <='0';
          end if;
        if(cVar1S23S41N048N018P032P028(0)='1' AND  D( 9)='1' AND B( 1)='1' )then
          cVar2S23S41P065P037nsss(0) <='1';
          else
          cVar2S23S41P065P037nsss(0) <='0';
          end if;
        if(cVar1S24S41N048N018N032P056(0)='1' AND  A( 3)='1' AND B( 4)='1' )then
          cVar2S24S41P013P031nsss(0) <='1';
          else
          cVar2S24S41P013P031nsss(0) <='0';
          end if;
        if(cVar1S25S41N048N018N032P056(0)='1' AND  A( 3)='1' AND B( 4)='0' AND A(14)='1' )then
          cVar2S25S41P013N031P010nsss(0) <='1';
          else
          cVar2S25S41P013N031P010nsss(0) <='0';
          end if;
        if(cVar1S26S41N048N018N032P056(0)='1' AND  A( 3)='0' AND A( 4)='1' )then
          cVar2S26S41N013P011nsss(0) <='1';
          else
          cVar2S26S41N013P011nsss(0) <='0';
          end if;
        if(cVar1S27S41N048N018N032P056(0)='1' AND  A( 3)='0' AND A( 4)='0' AND A(14)='1' )then
          cVar2S27S41N013N011P010nsss(0) <='1';
          else
          cVar2S27S41N013N011P010nsss(0) <='0';
          end if;
        if(cVar1S28S41N048N018N032N056(0)='1' AND  B( 2)='1' AND A(13)='0' AND A( 1)='1' )then
          cVar2S28S41P035P012P017nsss(0) <='1';
          else
          cVar2S28S41P035P012P017nsss(0) <='0';
          end if;
        if(cVar1S29S41N048N018N032N056(0)='1' AND  B( 2)='1' AND A(13)='1' AND A(12)='1' )then
          cVar2S29S41P035P012P014nsss(0) <='1';
          else
          cVar2S29S41P035P012P014nsss(0) <='0';
          end if;
        if(cVar1S30S41N048N018N032N056(0)='1' AND  B( 2)='0' AND B(17)='1' AND A(16)='1' )then
          cVar2S30S41N035P024P006nsss(0) <='1';
          else
          cVar2S30S41N035P024P006nsss(0) <='0';
          end if;
        if(cVar1S1S42P018P048N025P027(0)='1' AND  A( 5)='1' )then
          cVar2S1S42P009nsss(0) <='1';
          else
          cVar2S1S42P009nsss(0) <='0';
          end if;
        if(cVar1S2S42P018P048N025P027(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S2S42N009P006nsss(0) <='1';
          else
          cVar2S2S42N009P006nsss(0) <='0';
          end if;
        if(cVar1S3S42P018P048N025P027(0)='1' AND  A( 5)='0' AND A(16)='0' AND A(15)='1' )then
          cVar2S3S42N009N006P008nsss(0) <='1';
          else
          cVar2S3S42N009N006P008nsss(0) <='0';
          end if;
        if(cVar1S4S42P018P048N025N027(0)='1' AND  E( 2)='1' AND E( 1)='0' )then
          cVar2S4S42P062P066nsss(0) <='1';
          else
          cVar2S4S42P062P066nsss(0) <='0';
          end if;
        if(cVar1S5S42P018P048N025N027(0)='1' AND  E( 2)='0' AND A(16)='1' )then
          cVar2S5S42N062P006nsss(0) <='1';
          else
          cVar2S5S42N062P006nsss(0) <='0';
          end if;
        if(cVar1S6S42P018P048N025N027(0)='1' AND  E( 2)='0' AND A(16)='0' AND D( 7)='1' )then
          cVar2S6S42N062N006P040nsss(0) <='1';
          else
          cVar2S6S42N062N006P040nsss(0) <='0';
          end if;
        if(cVar1S8S42P018N048P038N002(0)='1' AND  A( 2)='0' AND B( 9)='1' )then
          cVar2S8S42P015P021nsss(0) <='1';
          else
          cVar2S8S42P015P021nsss(0) <='0';
          end if;
        if(cVar1S9S42P018N048P038N002(0)='1' AND  A( 2)='0' AND B( 9)='0' AND A(17)='1' )then
          cVar2S9S42P015N021P004nsss(0) <='1';
          else
          cVar2S9S42P015N021P004nsss(0) <='0';
          end if;
        if(cVar1S10S42P018N048N038P000(0)='1' AND  B(18)='1' AND E(15)='1' AND A(14)='0' )then
          cVar2S10S42P022P043P010nsss(0) <='1';
          else
          cVar2S10S42P022P043P010nsss(0) <='0';
          end if;
        if(cVar1S11S42P018N048N038P000(0)='1' AND  B(18)='1' AND E(15)='0' AND A( 6)='1' )then
          cVar2S11S42P022N043P007nsss(0) <='1';
          else
          cVar2S11S42P022N043P007nsss(0) <='0';
          end if;
        if(cVar1S12S42P018N048N038P000(0)='1' AND  B(18)='0' AND E( 6)='0' AND A( 7)='0' )then
          cVar2S12S42N022P046P005nsss(0) <='1';
          else
          cVar2S12S42N022P046P005nsss(0) <='0';
          end if;
        if(cVar1S13S42P018N048N038P000(0)='1' AND  B(18)='0' AND E( 6)='1' AND B( 7)='1' )then
          cVar2S13S42N022P046P025nsss(0) <='1';
          else
          cVar2S13S42N022P046P025nsss(0) <='0';
          end if;
        if(cVar1S14S42P018N048N038P000(0)='1' AND  E(14)='0' AND E(10)='0' AND E( 2)='0' )then
          cVar2S14S42P047P063P062nsss(0) <='1';
          else
          cVar2S14S42P047P063P062nsss(0) <='0';
          end if;
        if(cVar1S15S42P018P048P011P008(0)='1' AND  A(12)='1' )then
          cVar2S15S42P014nsss(0) <='1';
          else
          cVar2S15S42P014nsss(0) <='0';
          end if;
        if(cVar1S16S42P018P048P011P008(0)='1' AND  A(12)='0' AND A( 1)='0' )then
          cVar2S16S42N014P017nsss(0) <='1';
          else
          cVar2S16S42N014P017nsss(0) <='0';
          end if;
        if(cVar1S17S42P018P048P011P008(0)='1' AND  A(12)='0' AND A( 1)='1' AND E( 6)='0' )then
          cVar2S17S42N014P017P046nsss(0) <='1';
          else
          cVar2S17S42N014P017P046nsss(0) <='0';
          end if;
        if(cVar1S18S42P018P048P011P008(0)='1' AND  A(11)='0' )then
          cVar2S18S42P016nsss(0) <='1';
          else
          cVar2S18S42P016nsss(0) <='0';
          end if;
        if(cVar1S19S42P018P048P011P013(0)='1' AND  A( 1)='1' )then
          cVar2S19S42P017nsss(0) <='1';
          else
          cVar2S19S42P017nsss(0) <='0';
          end if;
        if(cVar1S21S42P018N048P044N023(0)='1' AND  E( 6)='1' )then
          cVar2S21S42P046nsss(0) <='1';
          else
          cVar2S21S42P046nsss(0) <='0';
          end if;
        if(cVar1S22S42P018N048P044N023(0)='1' AND  E( 6)='0' AND A( 2)='0' )then
          cVar2S22S42N046P015nsss(0) <='1';
          else
          cVar2S22S42N046P015nsss(0) <='0';
          end if;
        if(cVar1S23S42P018N048N044P004(0)='1' AND  E( 7)='0' AND B( 8)='1' AND E( 9)='1' )then
          cVar2S23S42P042P023P067nsss(0) <='1';
          else
          cVar2S23S42P042P023P067nsss(0) <='0';
          end if;
        if(cVar1S24S42P018N048N044P004(0)='1' AND  E( 7)='1' AND E( 1)='0' AND A( 3)='1' )then
          cVar2S24S42P042P066P013nsss(0) <='1';
          else
          cVar2S24S42P042P066P013nsss(0) <='0';
          end if;
        if(cVar1S25S42P018N048N044P004(0)='1' AND  A( 1)='1' AND A( 0)='1' AND A(13)='0' )then
          cVar2S25S42P017P019P012nsss(0) <='1';
          else
          cVar2S25S42P017P019P012nsss(0) <='0';
          end if;
        if(cVar1S26S42P018N048N044P004(0)='1' AND  A( 1)='0' AND D(15)='1' )then
          cVar2S26S42N017P041nsss(0) <='1';
          else
          cVar2S26S42N017P041nsss(0) <='0';
          end if;
        if(cVar1S27S42P018N048N044P004(0)='1' AND  A( 1)='0' AND D(15)='0' AND A( 5)='1' )then
          cVar2S27S42N017N041P009nsss(0) <='1';
          else
          cVar2S27S42N017N041P009nsss(0) <='0';
          end if;
        if(cVar1S2S43P048P025N007N004(0)='1' AND  A( 5)='1' )then
          cVar2S2S43P009nsss(0) <='1';
          else
          cVar2S2S43P009nsss(0) <='0';
          end if;
        if(cVar1S3S43P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='1' )then
          cVar2S3S43N009P006nsss(0) <='1';
          else
          cVar2S3S43N009P006nsss(0) <='0';
          end if;
        if(cVar1S4S43P048P025N007N004(0)='1' AND  A( 5)='0' AND A(16)='0' AND A(15)='1' )then
          cVar2S4S43N009N006P008nsss(0) <='1';
          else
          cVar2S4S43N009N006P008nsss(0) <='0';
          end if;
        if(cVar1S6S43P048N025P062N058(0)='1' AND  B( 1)='0' )then
          cVar2S6S43P037nsss(0) <='1';
          else
          cVar2S6S43P037nsss(0) <='0';
          end if;
        if(cVar1S7S43P048N025N062P027(0)='1' AND  A( 6)='1' )then
          cVar2S7S43P007nsss(0) <='1';
          else
          cVar2S7S43P007nsss(0) <='0';
          end if;
        if(cVar1S8S43P048N025N062P027(0)='1' AND  A( 6)='0' AND A(16)='1' )then
          cVar2S8S43N007P006nsss(0) <='1';
          else
          cVar2S8S43N007P006nsss(0) <='0';
          end if;
        if(cVar1S9S43P048N025N062P027(0)='1' AND  A( 6)='0' AND A(16)='0' AND A( 5)='1' )then
          cVar2S9S43N007N006P009nsss(0) <='1';
          else
          cVar2S9S43N007N006P009nsss(0) <='0';
          end if;
        if(cVar1S10S43P048N025N062N027(0)='1' AND  D(14)='1' )then
          cVar2S10S43P045nsss(0) <='1';
          else
          cVar2S10S43P045nsss(0) <='0';
          end if;
        if(cVar1S11S43P048N025N062N027(0)='1' AND  D(14)='0' AND A(19)='0' )then
          cVar2S11S43N045P000nsss(0) <='1';
          else
          cVar2S11S43N045P000nsss(0) <='0';
          end if;
        if(cVar1S12S43N048P022P043P012(0)='1' AND  A(14)='0' )then
          cVar2S12S43P010nsss(0) <='1';
          else
          cVar2S12S43P010nsss(0) <='0';
          end if;
        if(cVar1S13S43N048P022N043P004(0)='1' AND  E( 7)='1' )then
          cVar2S13S43P042nsss(0) <='1';
          else
          cVar2S13S43P042nsss(0) <='0';
          end if;
        if(cVar1S14S43N048P022N043N004(0)='1' AND  D(13)='0' AND E( 9)='0' AND B(11)='1' )then
          cVar2S14S43P049P067P036nsss(0) <='1';
          else
          cVar2S14S43P049P067P036nsss(0) <='0';
          end if;
        if(cVar1S15S43N048N022P038P021(0)='1' AND  A(18)='1' )then
          cVar2S15S43P002nsss(0) <='1';
          else
          cVar2S15S43P002nsss(0) <='0';
          end if;
        if(cVar1S16S43N048N022P038P021(0)='1' AND  A(18)='0' AND A( 2)='0' )then
          cVar2S16S43N002P015nsss(0) <='1';
          else
          cVar2S16S43N002P015nsss(0) <='0';
          end if;
        if(cVar1S17S43N048N022P038N021(0)='1' AND  D(15)='1' )then
          cVar2S17S43P041nsss(0) <='1';
          else
          cVar2S17S43P041nsss(0) <='0';
          end if;
        if(cVar1S18S43N048N022P038N021(0)='1' AND  D(15)='0' AND E( 9)='0' AND A( 8)='0' )then
          cVar2S18S43N041P067P003nsss(0) <='1';
          else
          cVar2S18S43N041P067P003nsss(0) <='0';
          end if;
        if(cVar1S19S43N048N022N038P004(0)='1' AND  A(15)='1' AND D(13)='1' )then
          cVar2S19S43P008P049nsss(0) <='1';
          else
          cVar2S19S43P008P049nsss(0) <='0';
          end if;
        if(cVar1S20S43N048N022N038P004(0)='1' AND  A(15)='1' AND D(13)='0' AND E(13)='1' )then
          cVar2S20S43P008N049P051nsss(0) <='1';
          else
          cVar2S20S43P008N049P051nsss(0) <='0';
          end if;
        if(cVar1S21S43N048N022N038P004(0)='1' AND  A(15)='0' AND B(14)='1' AND A(13)='1' )then
          cVar2S21S43N008P030P012nsss(0) <='1';
          else
          cVar2S21S43N008P030P012nsss(0) <='0';
          end if;
        if(cVar1S22S43N048N022N038P004(0)='1' AND  E( 7)='1' )then
          cVar2S22S43P042nsss(0) <='1';
          else
          cVar2S22S43P042nsss(0) <='0';
          end if;
        if(cVar1S23S43N048N022N038P004(0)='1' AND  E( 7)='0' AND A( 1)='1' AND A(13)='0' )then
          cVar2S23S43N042P017P012nsss(0) <='1';
          else
          cVar2S23S43N042P017P012nsss(0) <='0';
          end if;
        if(cVar1S24S43N048N022N038P004(0)='1' AND  E( 7)='0' AND A( 1)='0' AND D(14)='1' )then
          cVar2S24S43N042N017P045nsss(0) <='1';
          else
          cVar2S24S43N042N017P045nsss(0) <='0';
          end if;
        if(cVar1S3S44P022N043N004P047(0)='1' AND  E( 9)='0' AND A( 1)='0' )then
          cVar2S3S44P067P017nsss(0) <='1';
          else
          cVar2S3S44P067P017nsss(0) <='0';
          end if;
        if(cVar1S4S44N022P004P043P045(0)='1' AND  A(15)='1' )then
          cVar2S4S44P008nsss(0) <='1';
          else
          cVar2S4S44P008nsss(0) <='0';
          end if;
        if(cVar1S5S44N022P004P043P045(0)='1' AND  A(15)='0' AND E(14)='0' AND A(16)='0' )then
          cVar2S5S44N008P047P006nsss(0) <='1';
          else
          cVar2S5S44N008P047P006nsss(0) <='0';
          end if;
        if(cVar1S6S44N022P004P043P045(0)='1' AND  A(15)='0' AND E(14)='1' AND A(16)='1' )then
          cVar2S6S44N008P047P006nsss(0) <='1';
          else
          cVar2S6S44N008P047P006nsss(0) <='0';
          end if;
        if(cVar1S7S44N022P004P043P045(0)='1' AND  E(14)='1' AND A(16)='1' )then
          cVar2S7S44P047P006nsss(0) <='1';
          else
          cVar2S7S44P047P006nsss(0) <='0';
          end if;
        if(cVar1S8S44N022P004P043P045(0)='1' AND  E(14)='1' AND A(16)='0' AND A( 1)='0' )then
          cVar2S8S44P047N006P017nsss(0) <='1';
          else
          cVar2S8S44P047N006P017nsss(0) <='0';
          end if;
        if(cVar1S9S44N022P004P043P045(0)='1' AND  E(14)='0' AND E(13)='1' )then
          cVar2S9S44N047P051nsss(0) <='1';
          else
          cVar2S9S44N047P051nsss(0) <='0';
          end if;
        if(cVar1S10S44N022P004P043P045(0)='1' AND  E(14)='0' AND E(13)='0' AND D( 6)='1' )then
          cVar2S10S44N047N051P044nsss(0) <='1';
          else
          cVar2S10S44N047N051P044nsss(0) <='0';
          end if;
        if(cVar1S11S44N022P004P043P023(0)='1' AND  A( 7)='1' )then
          cVar2S11S44P005nsss(0) <='1';
          else
          cVar2S11S44P005nsss(0) <='0';
          end if;
        if(cVar1S12S44N022P004P043P023(0)='1' AND  A( 7)='0' AND D( 6)='0' )then
          cVar2S12S44N005P044nsss(0) <='1';
          else
          cVar2S12S44N005P044nsss(0) <='0';
          end if;
        if(cVar1S13S44N022P004P043N023(0)='1' AND  A(16)='1' )then
          cVar2S13S44P006nsss(0) <='1';
          else
          cVar2S13S44P006nsss(0) <='0';
          end if;
        if(cVar1S14S44N022P004P043N023(0)='1' AND  A(16)='0' AND A( 6)='1' )then
          cVar2S14S44N006P007nsss(0) <='1';
          else
          cVar2S14S44N006P007nsss(0) <='0';
          end if;
        if(cVar1S15S44N022P004P043N023(0)='1' AND  A(16)='0' AND A( 6)='0' AND A( 8)='1' )then
          cVar2S15S44N006N007P003nsss(0) <='1';
          else
          cVar2S15S44N006N007P003nsss(0) <='0';
          end if;
        if(cVar1S17S44N022P004N040P017(0)='1' AND  A(13)='0' AND D( 5)='1' )then
          cVar2S17S44P012P048nsss(0) <='1';
          else
          cVar2S17S44P012P048nsss(0) <='0';
          end if;
        if(cVar1S18S44N022P004N040P017(0)='1' AND  A(13)='0' AND D( 5)='0' AND A(11)='1' )then
          cVar2S18S44P012N048P016nsss(0) <='1';
          else
          cVar2S18S44P012N048P016nsss(0) <='0';
          end if;
        if(cVar1S19S44N022P004N040N017(0)='1' AND  D( 6)='1' AND B( 8)='1' )then
          cVar2S19S44P044P023nsss(0) <='1';
          else
          cVar2S19S44P044P023nsss(0) <='0';
          end if;
        if(cVar1S20S44N022P004N040N017(0)='1' AND  D( 6)='0' AND A( 2)='1' AND A(18)='1' )then
          cVar2S20S44N044P015P002nsss(0) <='1';
          else
          cVar2S20S44N044P015P002nsss(0) <='0';
          end if;
        if(cVar1S21S44N022P004N040N017(0)='1' AND  D( 6)='0' AND A( 2)='0' AND D(14)='1' )then
          cVar2S21S44N044N015P045nsss(0) <='1';
          else
          cVar2S21S44N044N015P045nsss(0) <='0';
          end if;
        if(cVar1S1S45P022P043N019P012(0)='1' AND  A( 3)='0' )then
          cVar2S1S45P013nsss(0) <='1';
          else
          cVar2S1S45P013nsss(0) <='0';
          end if;
        if(cVar1S4S45P022N043N004N007(0)='1' AND  B( 3)='1' )then
          cVar2S4S45P033nsss(0) <='1';
          else
          cVar2S4S45P033nsss(0) <='0';
          end if;
        if(cVar1S5S45P022N043N004N007(0)='1' AND  B( 3)='0' AND A(18)='1' )then
          cVar2S5S45N033P002nsss(0) <='1';
          else
          cVar2S5S45N033P002nsss(0) <='0';
          end if;
        if(cVar1S6S45P022N043N004N007(0)='1' AND  B( 3)='0' AND A(18)='0' AND A(15)='1' )then
          cVar2S6S45N033N002P008nsss(0) <='1';
          else
          cVar2S6S45N033N002P008nsss(0) <='0';
          end if;
        if(cVar1S8S45N022P047N006P008(0)='1' AND  B(16)='1' AND A(10)='1' )then
          cVar2S8S45P026P018nsss(0) <='1';
          else
          cVar2S8S45P026P018nsss(0) <='0';
          end if;
        if(cVar1S9S45N022P047N006P008(0)='1' AND  B(16)='1' AND A(10)='0' AND E( 5)='0' )then
          cVar2S9S45P026N018P050nsss(0) <='1';
          else
          cVar2S9S45P026N018P050nsss(0) <='0';
          end if;
        if(cVar1S10S45N022P047N006P008(0)='1' AND  B(16)='0' AND B(17)='1' )then
          cVar2S10S45N026P024nsss(0) <='1';
          else
          cVar2S10S45N026P024nsss(0) <='0';
          end if;
        if(cVar1S11S45N022P047N006N008(0)='1' AND  A( 6)='1' AND A( 2)='0' )then
          cVar2S11S45P007P015nsss(0) <='1';
          else
          cVar2S11S45P007P015nsss(0) <='0';
          end if;
        if(cVar1S12S45N022P047N006N008(0)='1' AND  A( 6)='0' AND A( 5)='1' AND E(13)='0' )then
          cVar2S12S45N007P009P051nsss(0) <='1';
          else
          cVar2S12S45N007P009P051nsss(0) <='0';
          end if;
        if(cVar1S13S45N022P047N006N008(0)='1' AND  A( 6)='0' AND A( 5)='0' AND D( 8)='1' )then
          cVar2S13S45N007N009P069nsss(0) <='1';
          else
          cVar2S13S45N007N009P069nsss(0) <='0';
          end if;
        if(cVar1S14S45N022N047P051P008(0)='1' AND  B(15)='1' )then
          cVar2S14S45P028nsss(0) <='1';
          else
          cVar2S14S45P028nsss(0) <='0';
          end if;
        if(cVar1S15S45N022N047P051P008(0)='1' AND  B(15)='0' AND B(16)='1' AND E( 1)='0' )then
          cVar2S15S45N028P026P066nsss(0) <='1';
          else
          cVar2S15S45N028P026P066nsss(0) <='0';
          end if;
        if(cVar1S16S45N022N047P051P008(0)='1' AND  B(15)='0' AND B(16)='0' AND D(12)='1' )then
          cVar2S16S45N028N026P053nsss(0) <='1';
          else
          cVar2S16S45N028N026P053nsss(0) <='0';
          end if;
        if(cVar1S17S45N022N047P051N008(0)='1' AND  B( 6)='1' AND A( 5)='1' )then
          cVar2S17S45P027P009nsss(0) <='1';
          else
          cVar2S17S45P027P009nsss(0) <='0';
          end if;
        if(cVar1S18S45N022N047P051N008(0)='1' AND  B( 6)='1' AND A( 5)='0' AND A( 4)='1' )then
          cVar2S18S45P027N009P011nsss(0) <='1';
          else
          cVar2S18S45P027N009P011nsss(0) <='0';
          end if;
        if(cVar1S19S45N022N047P051N008(0)='1' AND  B( 6)='0' AND A( 4)='1' )then
          cVar2S19S45N027P011nsss(0) <='1';
          else
          cVar2S19S45N027P011nsss(0) <='0';
          end if;
        if(cVar1S20S45N022N047N051P049(0)='1' AND  B( 8)='1' AND A( 7)='1' AND D( 0)='0' )then
          cVar2S20S45P023P005P068nsss(0) <='1';
          else
          cVar2S20S45P023P005P068nsss(0) <='0';
          end if;
        if(cVar1S21S45N022N047N051P049(0)='1' AND  B( 8)='1' AND A( 7)='0' AND A(17)='1' )then
          cVar2S21S45P023N005P004nsss(0) <='1';
          else
          cVar2S21S45P023N005P004nsss(0) <='0';
          end if;
        if(cVar1S22S45N022N047N051P049(0)='1' AND  B( 8)='0' AND E(15)='1' AND B(17)='1' )then
          cVar2S22S45N023P043P024nsss(0) <='1';
          else
          cVar2S22S45N023P043P024nsss(0) <='0';
          end if;
        if(cVar1S23S45N022N047N051P049(0)='1' AND  B( 3)='1' )then
          cVar2S23S45P033nsss(0) <='1';
          else
          cVar2S23S45P033nsss(0) <='0';
          end if;
        if(cVar1S24S45N022N047N051P049(0)='1' AND  B( 3)='0' AND B(12)='1' )then
          cVar2S24S45N033P034nsss(0) <='1';
          else
          cVar2S24S45N033P034nsss(0) <='0';
          end if;
        if(cVar1S3S46P022N043N004P047(0)='1' AND  D(10)='1' )then
          cVar2S3S46P061nsss(0) <='1';
          else
          cVar2S3S46P061nsss(0) <='0';
          end if;
        if(cVar1S4S46P022N043N004P047(0)='1' AND  D(10)='0' AND D( 8)='0' AND A( 8)='0' )then
          cVar2S4S46N061P069P003nsss(0) <='1';
          else
          cVar2S4S46N061P069P003nsss(0) <='0';
          end if;
        if(cVar1S5S46N022P048P025P050(0)='1' AND  E( 9)='0' )then
          cVar2S5S46P067nsss(0) <='1';
          else
          cVar2S5S46P067nsss(0) <='0';
          end if;
        if(cVar1S6S46N022P048N025P043(0)='1' AND  D(14)='1' )then
          cVar2S6S46P045nsss(0) <='1';
          else
          cVar2S6S46P045nsss(0) <='0';
          end if;
        if(cVar1S7S46N022P048N025P043(0)='1' AND  D(14)='0' AND D( 4)='0' )then
          cVar2S7S46N045P052nsss(0) <='1';
          else
          cVar2S7S46N045P052nsss(0) <='0';
          end if;
        if(cVar1S8S46N022P048N025P043(0)='1' AND  D(14)='0' AND D( 4)='1' AND A( 2)='1' )then
          cVar2S8S46N045P052P015nsss(0) <='1';
          else
          cVar2S8S46N045P052P015nsss(0) <='0';
          end if;
        if(cVar1S9S46N022N048P037P065(0)='1' AND  B( 7)='0' AND E(11)='0' AND B( 6)='0' )then
          cVar2S9S46P025P059P027nsss(0) <='1';
          else
          cVar2S9S46P025P059P027nsss(0) <='0';
          end if;
        if(cVar1S10S46N022N048P037P065(0)='1' AND  B( 7)='0' AND E(11)='1' AND A( 8)='0' )then
          cVar2S10S46P025P059P003nsss(0) <='1';
          else
          cVar2S10S46P025P059P003nsss(0) <='0';
          end if;
        if(cVar1S11S46N022N048P037P065(0)='1' AND  B( 7)='1' AND A(12)='1' )then
          cVar2S11S46P025P014nsss(0) <='1';
          else
          cVar2S11S46P025P014nsss(0) <='0';
          end if;
        if(cVar1S12S46N022N048P037P065(0)='1' AND  E( 2)='0' AND D( 8)='1' AND E( 9)='1' )then
          cVar2S12S46P062P069P067nsss(0) <='1';
          else
          cVar2S12S46P062P069P067nsss(0) <='0';
          end if;
        if(cVar1S13S46N022N048P037P065(0)='1' AND  E( 2)='0' AND D( 8)='0' AND D( 0)='0' )then
          cVar2S13S46P062N069P068nsss(0) <='1';
          else
          cVar2S13S46P062N069P068nsss(0) <='0';
          end if;
        if(cVar1S14S46N022N048N037P023(0)='1' AND  A( 7)='1' AND B( 0)='0' )then
          cVar2S14S46P005P039nsss(0) <='1';
          else
          cVar2S14S46P005P039nsss(0) <='0';
          end if;
        if(cVar1S15S46N022N048N037P023(0)='1' AND  A( 7)='0' AND A(17)='1' )then
          cVar2S15S46N005P004nsss(0) <='1';
          else
          cVar2S15S46N005P004nsss(0) <='0';
          end if;
        if(cVar1S16S46N022N048N037P023(0)='1' AND  A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S16S46N005N004P006nsss(0) <='1';
          else
          cVar2S16S46N005N004P006nsss(0) <='0';
          end if;
        if(cVar1S17S46N022N048N037N023(0)='1' AND  E(15)='0' AND D(14)='0' )then
          cVar2S17S46P043P045nsss(0) <='1';
          else
          cVar2S17S46P043P045nsss(0) <='0';
          end if;
        if(cVar1S18S46N022N048N037N023(0)='1' AND  E(15)='0' AND D(14)='1' AND B(17)='1' )then
          cVar2S18S46P043P045P024nsss(0) <='1';
          else
          cVar2S18S46P043P045P024nsss(0) <='0';
          end if;
        if(cVar1S19S46N022N048N037N023(0)='1' AND  E(15)='1' AND A(16)='1' )then
          cVar2S19S46P043P006nsss(0) <='1';
          else
          cVar2S19S46P043P006nsss(0) <='0';
          end if;
        if(cVar1S20S46N022N048N037N023(0)='1' AND  E(15)='1' AND A(16)='0' AND A( 6)='1' )then
          cVar2S20S46P043N006P007nsss(0) <='1';
          else
          cVar2S20S46P043N006P007nsss(0) <='0';
          end if;
        if(cVar1S1S47P022P043N019P013(0)='1' AND  A(17)='1' )then
          cVar2S1S47P004nsss(0) <='1';
          else
          cVar2S1S47P004nsss(0) <='0';
          end if;
        if(cVar1S2S47P022P043N019P013(0)='1' AND  A(17)='0' AND A( 7)='1' )then
          cVar2S2S47N004P005nsss(0) <='1';
          else
          cVar2S2S47N004P005nsss(0) <='0';
          end if;
        if(cVar1S3S47P022P043N019P013(0)='1' AND  A(17)='0' AND A( 7)='0' AND A( 6)='1' )then
          cVar2S3S47N004N005P007nsss(0) <='1';
          else
          cVar2S3S47N004N005P007nsss(0) <='0';
          end if;
        if(cVar1S5S47P022N043N004P047(0)='1' AND  D(10)='1' )then
          cVar2S5S47P061nsss(0) <='1';
          else
          cVar2S5S47P061nsss(0) <='0';
          end if;
        if(cVar1S6S47P022N043N004P047(0)='1' AND  D(10)='0' AND E( 9)='0' AND B(11)='1' )then
          cVar2S6S47N061P067P036nsss(0) <='1';
          else
          cVar2S6S47N061P067P036nsss(0) <='0';
          end if;
        if(cVar1S7S47N022P023P005P068(0)='1' AND  E(15)='1' )then
          cVar2S7S47P043nsss(0) <='1';
          else
          cVar2S7S47P043nsss(0) <='0';
          end if;
        if(cVar1S8S47N022P023P005P068(0)='1' AND  E(15)='0' AND E( 7)='1' )then
          cVar2S8S47N043P042nsss(0) <='1';
          else
          cVar2S8S47N043P042nsss(0) <='0';
          end if;
        if(cVar1S9S47N022P023N005P034(0)='1' AND  A( 6)='1' )then
          cVar2S9S47P007nsss(0) <='1';
          else
          cVar2S9S47P007nsss(0) <='0';
          end if;
        if(cVar1S10S47N022P023N005P034(0)='1' AND  A( 6)='0' AND A(17)='1' )then
          cVar2S10S47N007P004nsss(0) <='1';
          else
          cVar2S10S47N007P004nsss(0) <='0';
          end if;
        if(cVar1S11S47N022P023N005P034(0)='1' AND  A( 6)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S11S47N007N004P006nsss(0) <='1';
          else
          cVar2S11S47N007N004P006nsss(0) <='0';
          end if;
        if(cVar1S12S47N022N023P043P048(0)='1' AND  B( 7)='1' AND E( 5)='0' AND E( 9)='0' )then
          cVar2S12S47P025P050P067nsss(0) <='1';
          else
          cVar2S12S47P025P050P067nsss(0) <='0';
          end if;
        if(cVar1S13S47N022N023P043P048(0)='1' AND  B( 7)='0' AND D(14)='1' )then
          cVar2S13S47N025P045nsss(0) <='1';
          else
          cVar2S13S47N025P045nsss(0) <='0';
          end if;
        if(cVar1S14S47N022N023P043P048(0)='1' AND  B( 7)='0' AND D(14)='0' AND B(11)='0' )then
          cVar2S14S47N025N045P036nsss(0) <='1';
          else
          cVar2S14S47N025N045P036nsss(0) <='0';
          end if;
        if(cVar1S15S47N022N023P043N048(0)='1' AND  D(14)='0' AND B( 1)='1' AND B( 7)='0' )then
          cVar2S15S47P045P037P025nsss(0) <='1';
          else
          cVar2S15S47P045P037P025nsss(0) <='0';
          end if;
        if(cVar1S16S47N022N023P043N048(0)='1' AND  D(14)='0' AND B( 1)='0' AND A(11)='1' )then
          cVar2S16S47P045N037P016nsss(0) <='1';
          else
          cVar2S16S47P045N037P016nsss(0) <='0';
          end if;
        if(cVar1S17S47N022N023P043N048(0)='1' AND  D(14)='1' AND E(14)='1' )then
          cVar2S17S47P045P047nsss(0) <='1';
          else
          cVar2S17S47P045P047nsss(0) <='0';
          end if;
        if(cVar1S18S47N022N023P043N048(0)='1' AND  D(14)='1' AND E(14)='0' AND D( 2)='1' )then
          cVar2S18S47P045N047P060nsss(0) <='1';
          else
          cVar2S18S47P045N047P060nsss(0) <='0';
          end if;
        if(cVar1S20S47N022N023P043N006(0)='1' AND  A( 6)='1' AND B( 7)='1' )then
          cVar2S20S47P007P025nsss(0) <='1';
          else
          cVar2S20S47P007P025nsss(0) <='0';
          end if;
        if(cVar1S21S47N022N023P043N006(0)='1' AND  A( 6)='1' AND B( 7)='0' AND B(17)='1' )then
          cVar2S21S47P007N025P024nsss(0) <='1';
          else
          cVar2S21S47P007N025P024nsss(0) <='0';
          end if;
        if(cVar1S22S47N022N023P043N006(0)='1' AND  A( 6)='0' AND E(11)='1' )then
          cVar2S22S47N007P059nsss(0) <='1';
          else
          cVar2S22S47N007P059nsss(0) <='0';
          end if;
        if(cVar1S23S47N022N023P043N006(0)='1' AND  A( 6)='0' AND E(11)='0' AND B(19)='1' )then
          cVar2S23S47N007N059P020nsss(0) <='1';
          else
          cVar2S23S47N007N059P020nsss(0) <='0';
          end if;
        if(cVar1S0S48P016P065P034P059(0)='1' AND  E(12)='0' AND D( 3)='0' AND D( 2)='0' )then
          cVar2S0S48P055P056P060nsss(0) <='1';
          else
          cVar2S0S48P055P056P060nsss(0) <='0';
          end if;
        if(cVar1S1S48P016P065P034P059(0)='1' AND  E(12)='1' AND A( 1)='1' )then
          cVar2S1S48P055P017nsss(0) <='1';
          else
          cVar2S1S48P055P017nsss(0) <='0';
          end if;
        if(cVar1S2S48P016P065P034N059(0)='1' AND  B( 8)='1' AND A( 7)='1' )then
          cVar2S2S48P023P005nsss(0) <='1';
          else
          cVar2S2S48P023P005nsss(0) <='0';
          end if;
        if(cVar1S3S48P016P065P034N059(0)='1' AND  B( 8)='1' AND A( 7)='0' AND E( 7)='1' )then
          cVar2S3S48P023N005P042nsss(0) <='1';
          else
          cVar2S3S48P023N005P042nsss(0) <='0';
          end if;
        if(cVar1S4S48P016P065P034N059(0)='1' AND  B( 8)='0' AND B(15)='1' AND A(14)='1' )then
          cVar2S4S48N023P028P010nsss(0) <='1';
          else
          cVar2S4S48N023P028P010nsss(0) <='0';
          end if;
        if(cVar1S5S48P016P065P034N059(0)='1' AND  B( 8)='0' AND B(15)='0' )then
          cVar2S5S48N023N028psss(0) <='1';
          else
          cVar2S5S48N023N028psss(0) <='0';
          end if;
        if(cVar1S6S48P016P065P034P014(0)='1' AND  E( 2)='1' )then
          cVar2S6S48P062nsss(0) <='1';
          else
          cVar2S6S48P062nsss(0) <='0';
          end if;
        if(cVar1S7S48P016P065P034P014(0)='1' AND  E( 2)='0' AND E(11)='1' AND B(13)='0' )then
          cVar2S7S48N062P059P032nsss(0) <='1';
          else
          cVar2S7S48N062P059P032nsss(0) <='0';
          end if;
        if(cVar1S8S48P016P065P034P014(0)='1' AND  E( 2)='0' AND E(11)='0' AND B( 1)='1' )then
          cVar2S8S48N062N059P037nsss(0) <='1';
          else
          cVar2S8S48N062N059P037nsss(0) <='0';
          end if;
        if(cVar1S9S48P016P065P034N014(0)='1' AND  D( 1)='0' AND A(18)='1' )then
          cVar2S9S48P064P002nsss(0) <='1';
          else
          cVar2S9S48P064P002nsss(0) <='0';
          end if;
        if(cVar1S11S48P016P065P067P063(0)='1' AND  B( 2)='1' AND A(10)='1' )then
          cVar2S11S48P035P018nsss(0) <='1';
          else
          cVar2S11S48P035P018nsss(0) <='0';
          end if;
        if(cVar1S12S48P016P065P067P063(0)='1' AND  B( 2)='0' AND E( 2)='0' AND B(12)='1' )then
          cVar2S12S48N035P062P034nsss(0) <='1';
          else
          cVar2S12S48N035P062P034nsss(0) <='0';
          end if;
        if(cVar1S13S48P016P065N067P066(0)='1' AND  B(12)='1' AND A(12)='1' AND A( 2)='0' )then
          cVar2S13S48P034P014P015nsss(0) <='1';
          else
          cVar2S13S48P034P014P015nsss(0) <='0';
          end if;
        if(cVar1S14S48P016P065N067P066(0)='1' AND  B(12)='1' AND A(12)='0' AND A( 1)='1' )then
          cVar2S14S48P034N014P017nsss(0) <='1';
          else
          cVar2S14S48P034N014P017nsss(0) <='0';
          end if;
        if(cVar1S15S48P016P065N067P066(0)='1' AND  B(12)='0' AND B( 2)='1' AND E(10)='1' )then
          cVar2S15S48N034P035P063nsss(0) <='1';
          else
          cVar2S15S48N034P035P063nsss(0) <='0';
          end if;
        if(cVar1S16S48P016P065N067P066(0)='1' AND  A( 2)='1' AND A(10)='1' )then
          cVar2S16S48P015P018nsss(0) <='1';
          else
          cVar2S16S48P015P018nsss(0) <='0';
          end if;
        if(cVar1S17S48P016P065N067P066(0)='1' AND  A( 2)='0' AND A(13)='0' AND A(12)='1' )then
          cVar2S17S48N015P012P014nsss(0) <='1';
          else
          cVar2S17S48N015P012P014nsss(0) <='0';
          end if;
        if(cVar1S18S48P016P063P015P057(0)='1' AND  E( 1)='0' AND B(13)='0' )then
          cVar2S18S48P066P032nsss(0) <='1';
          else
          cVar2S18S48P066P032nsss(0) <='0';
          end if;
        if(cVar1S19S48P016P063P015P057(0)='1' AND  E( 1)='1' AND A(10)='1' AND B(11)='1' )then
          cVar2S19S48P066P018P036nsss(0) <='1';
          else
          cVar2S19S48P066P018P036nsss(0) <='0';
          end if;
        if(cVar1S20S48P016P063P015P057(0)='1' AND  E( 1)='1' AND A(10)='0' AND E( 9)='1' )then
          cVar2S20S48P066N018P067nsss(0) <='1';
          else
          cVar2S20S48P066N018P067nsss(0) <='0';
          end if;
        if(cVar1S21S48P016P063P015P056(0)='1' AND  A(10)='0' AND E( 2)='1' )then
          cVar2S21S48P018P062nsss(0) <='1';
          else
          cVar2S21S48P018P062nsss(0) <='0';
          end if;
        if(cVar1S22S48P016P063P015P056(0)='1' AND  A(10)='0' AND E( 2)='0' AND E( 1)='1' )then
          cVar2S22S48P018N062P066nsss(0) <='1';
          else
          cVar2S22S48P018N062P066nsss(0) <='0';
          end if;
        if(cVar1S23S48P016P063P015P056(0)='1' AND  A(10)='1' AND A( 3)='1' AND A( 0)='0' )then
          cVar2S23S48P018P013P019nsss(0) <='1';
          else
          cVar2S23S48P018P013P019nsss(0) <='0';
          end if;
        if(cVar1S24S48P016N063P052P061(0)='1' AND  A(17)='1' AND B(18)='1' )then
          cVar2S24S48P004P022nsss(0) <='1';
          else
          cVar2S24S48P004P022nsss(0) <='0';
          end if;
        if(cVar1S25S48P016N063P052P061(0)='1' AND  A(17)='1' AND B(18)='0' AND A( 0)='1' )then
          cVar2S25S48P004N022P019nsss(0) <='1';
          else
          cVar2S25S48P004N022P019nsss(0) <='0';
          end if;
        if(cVar1S26S48P016N063P052P061(0)='1' AND  A(17)='0' AND E( 2)='1' AND E(12)='0' )then
          cVar2S26S48N004P062P055nsss(0) <='1';
          else
          cVar2S26S48N004P062P055nsss(0) <='0';
          end if;
        if(cVar1S27S48P016N063P052P061(0)='1' AND  A(10)='1' AND A( 2)='1' AND A(12)='0' )then
          cVar2S27S48P018P015P014nsss(0) <='1';
          else
          cVar2S27S48P018P015P014nsss(0) <='0';
          end if;
        if(cVar1S28S48P016N063P052P061(0)='1' AND  A(10)='1' AND A( 2)='0' AND A(12)='1' )then
          cVar2S28S48P018N015P014nsss(0) <='1';
          else
          cVar2S28S48P018N015P014nsss(0) <='0';
          end if;
        if(cVar1S29S48P016N063P052P061(0)='1' AND  A(10)='0' AND B(13)='1' AND A( 2)='0' )then
          cVar2S29S48N018P032P015nsss(0) <='1';
          else
          cVar2S29S48N018P032P015nsss(0) <='0';
          end if;
        if(cVar1S30S48P016N063P052P060(0)='1' AND  B( 5)='1' AND A( 1)='1' )then
          cVar2S30S48P029P017nsss(0) <='1';
          else
          cVar2S30S48P029P017nsss(0) <='0';
          end if;
        if(cVar1S31S48P016N063P052P060(0)='1' AND  B( 5)='1' AND A( 1)='0' AND A( 5)='1' )then
          cVar2S31S48P029N017P009nsss(0) <='1';
          else
          cVar2S31S48P029N017P009nsss(0) <='0';
          end if;
        if(cVar1S2S49P023N005P034P007(0)='1' AND  E(15)='1' )then
          cVar2S2S49P043nsss(0) <='1';
          else
          cVar2S2S49P043nsss(0) <='0';
          end if;
        if(cVar1S3S49P023N005P034P007(0)='1' AND  E(15)='0' AND D( 6)='1' )then
          cVar2S3S49N043P044nsss(0) <='1';
          else
          cVar2S3S49N043P044nsss(0) <='0';
          end if;
        if(cVar1S4S49P023N005P034N007(0)='1' AND  E( 4)='1' )then
          cVar2S4S49P054nsss(0) <='1';
          else
          cVar2S4S49P054nsss(0) <='0';
          end if;
        if(cVar1S5S49P023N005P034N007(0)='1' AND  E( 4)='0' AND A(17)='1' AND D( 6)='1' )then
          cVar2S5S49N054P004P044nsss(0) <='1';
          else
          cVar2S5S49N054P004P044nsss(0) <='0';
          end if;
        if(cVar1S6S49P023N005P034N007(0)='1' AND  E( 4)='0' AND A(17)='0' AND A( 8)='1' )then
          cVar2S6S49N054N004P003nsss(0) <='1';
          else
          cVar2S6S49N054N004P003nsss(0) <='0';
          end if;
        if(cVar1S8S49N023P022P043N005(0)='1' AND  A( 0)='1' )then
          cVar2S8S49P019nsss(0) <='1';
          else
          cVar2S8S49P019nsss(0) <='0';
          end if;
        if(cVar1S9S49N023P022P043N005(0)='1' AND  A( 0)='0' AND A(17)='1' AND A(10)='0' )then
          cVar2S9S49N019P004P018nsss(0) <='1';
          else
          cVar2S9S49N019P004P018nsss(0) <='0';
          end if;
        if(cVar1S10S49N023P022P043N005(0)='1' AND  A( 0)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S10S49N019N004P007nsss(0) <='1';
          else
          cVar2S10S49N019N004P007nsss(0) <='0';
          end if;
        if(cVar1S12S49N023P022N043N004(0)='1' AND  A( 6)='1' )then
          cVar2S12S49P007nsss(0) <='1';
          else
          cVar2S12S49P007nsss(0) <='0';
          end if;
        if(cVar1S13S49N023P022N043N004(0)='1' AND  A( 6)='0' AND A(18)='1' )then
          cVar2S13S49N007P002nsss(0) <='1';
          else
          cVar2S13S49N007P002nsss(0) <='0';
          end if;
        if(cVar1S14S49N023P022N043N004(0)='1' AND  A( 6)='0' AND A(18)='0' AND A(10)='1' )then
          cVar2S14S49N007N002P018nsss(0) <='1';
          else
          cVar2S14S49N007N002P018nsss(0) <='0';
          end if;
        if(cVar1S15S49N023N022P016P035(0)='1' AND  B(12)='1' AND E(10)='1' AND B(11)='0' )then
          cVar2S15S49P034P063P036nsss(0) <='1';
          else
          cVar2S15S49P034P063P036nsss(0) <='0';
          end if;
        if(cVar1S16S49N023N022P016P035(0)='1' AND  B(12)='1' AND E(10)='0' AND E( 2)='1' )then
          cVar2S16S49P034N063P062nsss(0) <='1';
          else
          cVar2S16S49P034N063P062nsss(0) <='0';
          end if;
        if(cVar1S17S49N023N022P016P035(0)='1' AND  B(12)='0' AND B(11)='1' AND B( 1)='0' )then
          cVar2S17S49N034P036P037nsss(0) <='1';
          else
          cVar2S17S49N034P036P037nsss(0) <='0';
          end if;
        if(cVar1S18S49N023N022P016P035(0)='1' AND  E(13)='1' )then
          cVar2S18S49P051nsss(0) <='1';
          else
          cVar2S18S49P051nsss(0) <='0';
          end if;
        if(cVar1S19S49N023N022N016P028(0)='1' AND  A(14)='1' AND E(12)='1' AND A(13)='0' )then
          cVar2S19S49P010P055P012nsss(0) <='1';
          else
          cVar2S19S49P010P055P012nsss(0) <='0';
          end if;
        if(cVar1S20S49N023N022N016P028(0)='1' AND  A(14)='1' AND E(12)='0' AND E(13)='1' )then
          cVar2S20S49P010N055P051nsss(0) <='1';
          else
          cVar2S20S49P010N055P051nsss(0) <='0';
          end if;
        if(cVar1S21S49N023N022N016P028(0)='1' AND  A(14)='0' AND B( 5)='0' AND A(15)='1' )then
          cVar2S21S49N010P029P008nsss(0) <='1';
          else
          cVar2S21S49N010P029P008nsss(0) <='0';
          end if;
        if(cVar1S22S49N023N022N016N028(0)='1' AND  E(11)='1' AND B(13)='1' AND B( 2)='0' )then
          cVar2S22S49P059P032P035nsss(0) <='1';
          else
          cVar2S22S49P059P032P035nsss(0) <='0';
          end if;
        if(cVar1S23S49N023N022N016N028(0)='1' AND  E(11)='1' AND B(13)='0' AND A( 3)='1' )then
          cVar2S23S49P059N032P013nsss(0) <='1';
          else
          cVar2S23S49P059N032P013nsss(0) <='0';
          end if;
        if(cVar1S24S49N023N022N016N028(0)='1' AND  E(11)='0' AND E(14)='1' AND A(16)='1' )then
          cVar2S24S49N059P047P006nsss(0) <='1';
          else
          cVar2S24S49N059P047P006nsss(0) <='0';
          end if;
        if(cVar1S2S50P023N005P034P007(0)='1' AND  E(15)='1' )then
          cVar2S2S50P043nsss(0) <='1';
          else
          cVar2S2S50P043nsss(0) <='0';
          end if;
        if(cVar1S3S50P023N005P034P007(0)='1' AND  E(15)='0' AND A(10)='0' )then
          cVar2S3S50N043P018nsss(0) <='1';
          else
          cVar2S3S50N043P018nsss(0) <='0';
          end if;
        if(cVar1S4S50P023N005P034N007(0)='1' AND  D( 1)='1' )then
          cVar2S4S50P064nsss(0) <='1';
          else
          cVar2S4S50P064nsss(0) <='0';
          end if;
        if(cVar1S5S50P023N005P034N007(0)='1' AND  D( 1)='0' AND A(16)='1' )then
          cVar2S5S50N064P006nsss(0) <='1';
          else
          cVar2S5S50N064P006nsss(0) <='0';
          end if;
        if(cVar1S6S50N023P028P029P010(0)='1' AND  B( 4)='0' )then
          cVar2S6S50P031nsss(0) <='1';
          else
          cVar2S6S50P031nsss(0) <='0';
          end if;
        if(cVar1S7S50N023P028P029N010(0)='1' AND  A(15)='1' AND A(12)='0' )then
          cVar2S7S50P008P014nsss(0) <='1';
          else
          cVar2S7S50P008P014nsss(0) <='0';
          end if;
        if(cVar1S8S50N023P028P029N010(0)='1' AND  A(15)='0' AND E(10)='0' AND A( 4)='1' )then
          cVar2S8S50N008P063P011nsss(0) <='1';
          else
          cVar2S8S50N008P063P011nsss(0) <='0';
          end if;
        if(cVar1S9S50N023N028P053P025(0)='1' AND  A( 6)='1' )then
          cVar2S9S50P007nsss(0) <='1';
          else
          cVar2S9S50P007nsss(0) <='0';
          end if;
        if(cVar1S10S50N023N028P053P025(0)='1' AND  A( 6)='0' AND E( 6)='1' )then
          cVar2S10S50N007P046nsss(0) <='1';
          else
          cVar2S10S50N007P046nsss(0) <='0';
          end if;
        if(cVar1S11S50N023N028P053N025(0)='1' AND  B(17)='1' AND A(16)='1' AND A( 4)='0' )then
          cVar2S11S50P024P006P011nsss(0) <='1';
          else
          cVar2S11S50P024P006P011nsss(0) <='0';
          end if;
        if(cVar1S12S50N023N028P053N025(0)='1' AND  B(17)='1' AND A(16)='0' AND A(14)='0' )then
          cVar2S12S50P024N006P010nsss(0) <='1';
          else
          cVar2S12S50P024N006P010nsss(0) <='0';
          end if;
        if(cVar1S13S50N023N028P053N025(0)='1' AND  B(17)='0' AND D(14)='0' AND E(15)='0' )then
          cVar2S13S50N024P045P043nsss(0) <='1';
          else
          cVar2S13S50N024P045P043nsss(0) <='0';
          end if;
        if(cVar1S14S50N023N028P053N025(0)='1' AND  B(17)='0' AND D(14)='1' AND B(18)='1' )then
          cVar2S14S50N024P045P022nsss(0) <='1';
          else
          cVar2S14S50N024P045P022nsss(0) <='0';
          end if;
        if(cVar1S15S50N023N028P053P029(0)='1' AND  A( 4)='1' )then
          cVar2S15S50P011nsss(0) <='1';
          else
          cVar2S15S50P011nsss(0) <='0';
          end if;
        if(cVar1S16S50N023N028P053P029(0)='1' AND  A( 4)='0' AND A( 5)='1' )then
          cVar2S16S50N011P009nsss(0) <='1';
          else
          cVar2S16S50N011P009nsss(0) <='0';
          end if;
        if(cVar1S17S50N023N028P053N029(0)='1' AND  B(16)='1' AND B(11)='0' AND A( 4)='0' )then
          cVar2S17S50P026P036P011nsss(0) <='1';
          else
          cVar2S17S50P026P036P011nsss(0) <='0';
          end if;
        if(cVar1S18S50N023N028P053N029(0)='1' AND  B(16)='0' AND B( 6)='1' )then
          cVar2S18S50N026P027nsss(0) <='1';
          else
          cVar2S18S50N026P027nsss(0) <='0';
          end if;
        if(cVar1S19S50N023N028P053N029(0)='1' AND  B(16)='0' AND B( 6)='0' AND B( 2)='1' )then
          cVar2S19S50N026N027P035nsss(0) <='1';
          else
          cVar2S19S50N026N027P035nsss(0) <='0';
          end if;
        if(cVar1S0S51P028P029P010P031(0)='1' AND  D(12)='1' )then
          cVar2S0S51P053nsss(0) <='1';
          else
          cVar2S0S51P053nsss(0) <='0';
          end if;
        if(cVar1S1S51P028P029P010P031(0)='1' AND  D(12)='0' AND E(12)='1' AND A(13)='0' )then
          cVar2S1S51N053P055P012nsss(0) <='1';
          else
          cVar2S1S51N053P055P012nsss(0) <='0';
          end if;
        if(cVar1S2S51P028P029P010P031(0)='1' AND  D(12)='0' AND E(12)='0' AND E( 4)='1' )then
          cVar2S2S51N053N055P054nsss(0) <='1';
          else
          cVar2S2S51N053N055P054nsss(0) <='0';
          end if;
        if(cVar1S4S51P028P029N010N008(0)='1' AND  E(10)='0' AND D( 0)='0' AND A(12)='0' )then
          cVar2S4S51P063P068P014nsss(0) <='1';
          else
          cVar2S4S51P063P068P014nsss(0) <='0';
          end if;
        if(cVar1S6S51N028P023P005N042(0)='1' AND  E(15)='1' )then
          cVar2S6S51P043nsss(0) <='1';
          else
          cVar2S6S51P043nsss(0) <='0';
          end if;
        if(cVar1S7S51N028P023N005P049(0)='1' AND  B(16)='0' AND A( 6)='1' AND A( 2)='0' )then
          cVar2S7S51P026P007P015nsss(0) <='1';
          else
          cVar2S7S51P026P007P015nsss(0) <='0';
          end if;
        if(cVar1S8S51N028P023N005P049(0)='1' AND  B(16)='0' AND A( 6)='0' )then
          cVar2S8S51P026N007psss(0) <='1';
          else
          cVar2S8S51P026N007psss(0) <='0';
          end if;
        if(cVar1S10S51N028N023P025N007(0)='1' AND  E( 6)='1' )then
          cVar2S10S51P046nsss(0) <='1';
          else
          cVar2S10S51P046nsss(0) <='0';
          end if;
        if(cVar1S11S51N028N023P025N007(0)='1' AND  E( 6)='0' AND A( 8)='0' AND D(11)='1' )then
          cVar2S11S51N046P003P057nsss(0) <='1';
          else
          cVar2S11S51N046P003P057nsss(0) <='0';
          end if;
        if(cVar1S12S51N028N023N025P024(0)='1' AND  A(16)='1' AND E(14)='1' )then
          cVar2S12S51P006P047nsss(0) <='1';
          else
          cVar2S12S51P006P047nsss(0) <='0';
          end if;
        if(cVar1S13S51N028N023N025P024(0)='1' AND  A(16)='1' AND E(14)='0' AND E(15)='1' )then
          cVar2S13S51P006N047P043nsss(0) <='1';
          else
          cVar2S13S51P006N047P043nsss(0) <='0';
          end if;
        if(cVar1S14S51N028N023N025P024(0)='1' AND  A(16)='0' AND E(14)='1' )then
          cVar2S14S51N006P047nsss(0) <='1';
          else
          cVar2S14S51N006P047nsss(0) <='0';
          end if;
        if(cVar1S15S51N028N023N025N024(0)='1' AND  D(15)='1' AND B(19)='1' )then
          cVar2S15S51P041P020nsss(0) <='1';
          else
          cVar2S15S51P041P020nsss(0) <='0';
          end if;
        if(cVar1S16S51N028N023N025N024(0)='1' AND  D(15)='1' AND B(19)='0' AND A( 9)='1' )then
          cVar2S16S51P041N020P001nsss(0) <='1';
          else
          cVar2S16S51P041N020P001nsss(0) <='0';
          end if;
        if(cVar1S17S51N028N023N025N024(0)='1' AND  D(15)='0' AND B( 0)='1' AND D( 1)='1' )then
          cVar2S17S51N041P039P064nsss(0) <='1';
          else
          cVar2S17S51N041P039P064nsss(0) <='0';
          end if;
        if(cVar1S2S52P045P043N005N004(0)='1' AND  A(16)='1' )then
          cVar2S2S52P006nsss(0) <='1';
          else
          cVar2S2S52P006nsss(0) <='0';
          end if;
        if(cVar1S3S52P045P043N005N004(0)='1' AND  A(16)='0' AND A( 6)='1' AND A( 2)='0' )then
          cVar2S3S52N006P007P015nsss(0) <='1';
          else
          cVar2S3S52N006P007P015nsss(0) <='0';
          end if;
        if(cVar1S4S52P045P043N005N004(0)='1' AND  A(16)='0' AND A( 6)='0' AND A( 8)='1' )then
          cVar2S4S52N006N007P003nsss(0) <='1';
          else
          cVar2S4S52N006N007P003nsss(0) <='0';
          end if;
        if(cVar1S6S52P045N043P047N006(0)='1' AND  B(17)='1' )then
          cVar2S6S52P024nsss(0) <='1';
          else
          cVar2S6S52P024nsss(0) <='0';
          end if;
        if(cVar1S7S52P045N043P047N006(0)='1' AND  B(17)='0' AND A(11)='0' )then
          cVar2S7S52N024P016nsss(0) <='1';
          else
          cVar2S7S52N024P016nsss(0) <='0';
          end if;
        if(cVar1S9S52P045N043N047N048(0)='1' AND  D( 2)='1' )then
          cVar2S9S52P060nsss(0) <='1';
          else
          cVar2S9S52P060nsss(0) <='0';
          end if;
        if(cVar1S10S52P045N043N047N048(0)='1' AND  D( 2)='0' AND D( 6)='1' )then
          cVar2S10S52N060P044nsss(0) <='1';
          else
          cVar2S10S52N060P044nsss(0) <='0';
          end if;
        if(cVar1S11S52P045N043N047N048(0)='1' AND  D( 2)='0' AND D( 6)='0' AND E(10)='1' )then
          cVar2S11S52N060N044P063nsss(0) <='1';
          else
          cVar2S11S52N060N044P063nsss(0) <='0';
          end if;
        if(cVar1S12S52N045P028P010P055(0)='1' AND  A(13)='0' )then
          cVar2S12S52P012nsss(0) <='1';
          else
          cVar2S12S52P012nsss(0) <='0';
          end if;
        if(cVar1S13S52N045P028P010N055(0)='1' AND  B(12)='0' AND E( 4)='1' )then
          cVar2S13S52P034P054nsss(0) <='1';
          else
          cVar2S13S52P034P054nsss(0) <='0';
          end if;
        if(cVar1S14S52N045P028P010N055(0)='1' AND  B(12)='0' AND E( 4)='0' AND D(12)='1' )then
          cVar2S14S52P034N054P053nsss(0) <='1';
          else
          cVar2S14S52P034N054P053nsss(0) <='0';
          end if;
        if(cVar1S15S52N045P028N010P011(0)='1' AND  D(12)='1' )then
          cVar2S15S52P053nsss(0) <='1';
          else
          cVar2S15S52P053nsss(0) <='0';
          end if;
        if(cVar1S16S52N045P028N010P011(0)='1' AND  D(12)='0' AND D(11)='1' )then
          cVar2S16S52N053P057nsss(0) <='1';
          else
          cVar2S16S52N053P057nsss(0) <='0';
          end if;
        if(cVar1S17S52N045P028N010P011(0)='1' AND  D(12)='0' AND D(11)='0' AND A(11)='1' )then
          cVar2S17S52N053N057P016nsss(0) <='1';
          else
          cVar2S17S52N053N057P016nsss(0) <='0';
          end if;
        if(cVar1S18S52N045P028N010N011(0)='1' AND  B( 5)='0' AND A(15)='1' )then
          cVar2S18S52P029P008nsss(0) <='1';
          else
          cVar2S18S52P029P008nsss(0) <='0';
          end if;
        if(cVar1S19S52N045P028N010N011(0)='1' AND  B( 5)='0' AND A(15)='0' AND A(13)='1' )then
          cVar2S19S52P029N008P012nsss(0) <='1';
          else
          cVar2S19S52P029N008P012nsss(0) <='0';
          end if;
        if(cVar1S20S52N045N028P040P021(0)='1' AND  A(18)='1' )then
          cVar2S20S52P002nsss(0) <='1';
          else
          cVar2S20S52P002nsss(0) <='0';
          end if;
        if(cVar1S21S52N045N028P040P021(0)='1' AND  A(18)='0' AND A(11)='0' AND A( 1)='0' )then
          cVar2S21S52N002P016P017nsss(0) <='1';
          else
          cVar2S21S52N002P016P017nsss(0) <='0';
          end if;
        if(cVar1S22S52N045N028P040N021(0)='1' AND  B(19)='1' )then
          cVar2S22S52P020nsss(0) <='1';
          else
          cVar2S22S52P020nsss(0) <='0';
          end if;
        if(cVar1S23S52N045N028P040N021(0)='1' AND  B(19)='0' AND E( 1)='0' AND E( 5)='1' )then
          cVar2S23S52N020P066P050nsss(0) <='1';
          else
          cVar2S23S52N020P066P050nsss(0) <='0';
          end if;
        if(cVar1S24S52N045N028N040P025(0)='1' AND  E( 6)='1' AND E( 1)='0' )then
          cVar2S24S52P046P066nsss(0) <='1';
          else
          cVar2S24S52P046P066nsss(0) <='0';
          end if;
        if(cVar1S25S52N045N028N040P025(0)='1' AND  E( 6)='1' AND E( 1)='1' AND A(10)='0' )then
          cVar2S25S52P046P066P018nsss(0) <='1';
          else
          cVar2S25S52P046P066P018nsss(0) <='0';
          end if;
        if(cVar1S26S52N045N028N040P025(0)='1' AND  E( 6)='0' AND A( 6)='1' AND E(14)='1' )then
          cVar2S26S52N046P007P047nsss(0) <='1';
          else
          cVar2S26S52N046P007P047nsss(0) <='0';
          end if;
        if(cVar1S27S52N045N028N040N025(0)='1' AND  A( 2)='1' AND D( 3)='0' )then
          cVar2S27S52P015P056nsss(0) <='1';
          else
          cVar2S27S52P015P056nsss(0) <='0';
          end if;
        if(cVar1S28S52N045N028N040N025(0)='1' AND  A( 2)='1' AND D( 3)='1' AND D( 0)='1' )then
          cVar2S28S52P015P056P068nsss(0) <='1';
          else
          cVar2S28S52P015P056P068nsss(0) <='0';
          end if;
        if(cVar1S29S52N045N028N040N025(0)='1' AND  A( 2)='0' AND A( 7)='0' )then
          cVar2S29S52N015P005nsss(0) <='1';
          else
          cVar2S29S52N015P005nsss(0) <='0';
          end if;
        if(cVar1S30S52N045N028N040N025(0)='1' AND  A( 2)='0' AND A( 7)='1' AND B( 8)='1' )then
          cVar2S30S52N015P005P023nsss(0) <='1';
          else
          cVar2S30S52N015P005P023nsss(0) <='0';
          end if;
        if(cVar1S3S53P025N007P046N004(0)='1' AND  A(16)='1' )then
          cVar2S3S53P006nsss(0) <='1';
          else
          cVar2S3S53P006nsss(0) <='0';
          end if;
        if(cVar1S4S53P025N007P046N004(0)='1' AND  A(16)='0' AND D( 5)='1' )then
          cVar2S4S53N006P048nsss(0) <='1';
          else
          cVar2S4S53N006P048nsss(0) <='0';
          end if;
        if(cVar1S5S53P025N007N046P003(0)='1' AND  D(11)='1' )then
          cVar2S5S53P057nsss(0) <='1';
          else
          cVar2S5S53P057nsss(0) <='0';
          end if;
        if(cVar1S6S53P025N007N046P003(0)='1' AND  D(11)='0' AND B( 1)='0' AND B(12)='0' )then
          cVar2S6S53N057P037P034nsss(0) <='1';
          else
          cVar2S6S53N057P037P034nsss(0) <='0';
          end if;
        if(cVar1S8S53N025P028P010N055(0)='1' AND  A( 7)='0' AND A( 1)='1' )then
          cVar2S8S53P005P017nsss(0) <='1';
          else
          cVar2S8S53P005P017nsss(0) <='0';
          end if;
        if(cVar1S9S53N025P028P010N055(0)='1' AND  A( 7)='0' AND A( 1)='0' AND B(16)='0' )then
          cVar2S9S53P005N017P026nsss(0) <='1';
          else
          cVar2S9S53P005N017P026nsss(0) <='0';
          end if;
        if(cVar1S10S53N025P028N010P029(0)='1' AND  E(10)='0' AND D(12)='1' AND A(12)='0' )then
          cVar2S10S53P063P053P014nsss(0) <='1';
          else
          cVar2S10S53P063P053P014nsss(0) <='0';
          end if;
        if(cVar1S11S53N025P028N010P029(0)='1' AND  E(10)='0' AND D(12)='0' AND A(13)='1' )then
          cVar2S11S53P063N053P012nsss(0) <='1';
          else
          cVar2S11S53P063N053P012nsss(0) <='0';
          end if;
        if(cVar1S12S53N025P028N010P029(0)='1' AND  A( 4)='1' )then
          cVar2S12S53P011nsss(0) <='1';
          else
          cVar2S12S53P011nsss(0) <='0';
          end if;
        if(cVar1S13S53N025N028P040P021(0)='1' AND  A(18)='1' )then
          cVar2S13S53P002nsss(0) <='1';
          else
          cVar2S13S53P002nsss(0) <='0';
          end if;
        if(cVar1S14S53N025N028P040P021(0)='1' AND  A(18)='0' AND A( 2)='0' )then
          cVar2S14S53N002P015nsss(0) <='1';
          else
          cVar2S14S53N002P015nsss(0) <='0';
          end if;
        if(cVar1S15S53N025N028P040N021(0)='1' AND  E( 1)='0' AND B(19)='1' )then
          cVar2S15S53P066P020nsss(0) <='1';
          else
          cVar2S15S53P066P020nsss(0) <='0';
          end if;
        if(cVar1S16S53N025N028P040N021(0)='1' AND  E( 1)='0' AND B(19)='0' AND E(14)='1' )then
          cVar2S16S53P066N020P047nsss(0) <='1';
          else
          cVar2S16S53P066N020P047nsss(0) <='0';
          end if;
        if(cVar1S17S53N025N028N040P045(0)='1' AND  B(18)='1' )then
          cVar2S17S53P022nsss(0) <='1';
          else
          cVar2S17S53P022nsss(0) <='0';
          end if;
        if(cVar1S18S53N025N028N040P045(0)='1' AND  B(18)='0' AND B(17)='1' )then
          cVar2S18S53N022P024nsss(0) <='1';
          else
          cVar2S18S53N022P024nsss(0) <='0';
          end if;
        if(cVar1S19S53N025N028N040P045(0)='1' AND  B(18)='0' AND B(17)='0' AND B( 8)='1' )then
          cVar2S19S53N022N024P023nsss(0) <='1';
          else
          cVar2S19S53N022N024P023nsss(0) <='0';
          end if;
        if(cVar1S20S53N025N028N040N045(0)='1' AND  A( 2)='1' AND E(14)='0' AND D( 2)='1' )then
          cVar2S20S53P015P047P060nsss(0) <='1';
          else
          cVar2S20S53P015P047P060nsss(0) <='0';
          end if;
        if(cVar1S21S53N025N028N040N045(0)='1' AND  A( 2)='1' AND E(14)='1' AND B(16)='1' )then
          cVar2S21S53P015P047P026nsss(0) <='1';
          else
          cVar2S21S53P015P047P026nsss(0) <='0';
          end if;
        if(cVar1S22S53N025N028N040N045(0)='1' AND  A( 2)='0' AND A(10)='1' AND A(17)='0' )then
          cVar2S22S53N015P018P004nsss(0) <='1';
          else
          cVar2S22S53N015P018P004nsss(0) <='0';
          end if;
        if(cVar1S23S53N025N028N040N045(0)='1' AND  A( 2)='0' AND A(10)='0' AND A(11)='1' )then
          cVar2S23S53N015N018P016nsss(0) <='1';
          else
          cVar2S23S53N015N018P016nsss(0) <='0';
          end if;
        if(cVar1S2S54P018P040N002N004(0)='1' AND  A( 8)='1' AND A(12)='0' )then
          cVar2S2S54P003P014nsss(0) <='1';
          else
          cVar2S2S54P003P014nsss(0) <='0';
          end if;
        if(cVar1S3S54P018P040N002N004(0)='1' AND  A( 8)='0' AND A( 7)='1' )then
          cVar2S3S54N003P005nsss(0) <='1';
          else
          cVar2S3S54N003P005nsss(0) <='0';
          end if;
        if(cVar1S4S54P018P040N002N004(0)='1' AND  A( 8)='0' AND A( 7)='0' AND E( 5)='1' )then
          cVar2S4S54N003N005P050nsss(0) <='1';
          else
          cVar2S4S54N003N005P050nsss(0) <='0';
          end if;
        if(cVar1S6S54P018N040P045N004(0)='1' AND  B( 8)='1' )then
          cVar2S6S54P023nsss(0) <='1';
          else
          cVar2S6S54P023nsss(0) <='0';
          end if;
        if(cVar1S7S54P018N040P045N004(0)='1' AND  B( 8)='0' AND A(16)='1' )then
          cVar2S7S54N023P006nsss(0) <='1';
          else
          cVar2S7S54N023P006nsss(0) <='0';
          end if;
        if(cVar1S8S54P018N040P045N004(0)='1' AND  B( 8)='0' AND A(16)='0' AND A( 6)='1' )then
          cVar2S8S54N023N006P007nsss(0) <='1';
          else
          cVar2S8S54N023N006P007nsss(0) <='0';
          end if;
        if(cVar1S9S54P018N040N045P015(0)='1' AND  B(11)='0' AND E(14)='0' )then
          cVar2S9S54P036P047nsss(0) <='1';
          else
          cVar2S9S54P036P047nsss(0) <='0';
          end if;
        if(cVar1S10S54P018N040N045P015(0)='1' AND  B(11)='1' AND A( 5)='1' AND A( 0)='0' )then
          cVar2S10S54P036P009P019nsss(0) <='1';
          else
          cVar2S10S54P036P009P019nsss(0) <='0';
          end if;
        if(cVar1S11S54P018N040N045N015(0)='1' AND  B(15)='1' AND B( 5)='0' )then
          cVar2S11S54P028P029nsss(0) <='1';
          else
          cVar2S11S54P028P029nsss(0) <='0';
          end if;
        if(cVar1S12S54P018N040N045N015(0)='1' AND  B(15)='0' AND B( 7)='1' )then
          cVar2S12S54N028P025nsss(0) <='1';
          else
          cVar2S12S54N028P025nsss(0) <='0';
          end if;
        if(cVar1S13S54P018N040N045N015(0)='1' AND  B(15)='0' AND B( 7)='0' AND A(11)='0' )then
          cVar2S13S54N028N025P016nsss(0) <='1';
          else
          cVar2S13S54N028N025P016nsss(0) <='0';
          end if;
        if(cVar1S14S54P018P015P019P056(0)='1' AND  B( 6)='1' )then
          cVar2S14S54P027nsss(0) <='1';
          else
          cVar2S14S54P027nsss(0) <='0';
          end if;
        if(cVar1S15S54P018P015P019P056(0)='1' AND  B( 6)='0' AND D(14)='1' )then
          cVar2S15S54N027P045nsss(0) <='1';
          else
          cVar2S15S54N027P045nsss(0) <='0';
          end if;
        if(cVar1S16S54P018P015P019P056(0)='1' AND  B( 6)='0' AND D(14)='0' AND B( 8)='0' )then
          cVar2S16S54N027N045P023nsss(0) <='1';
          else
          cVar2S16S54N027N045P023nsss(0) <='0';
          end if;
        if(cVar1S17S54P018P015P019P056(0)='1' AND  A(13)='1' )then
          cVar2S17S54P012nsss(0) <='1';
          else
          cVar2S17S54P012nsss(0) <='0';
          end if;
        if(cVar1S19S54P018N015P019P007(0)='1' AND  A(16)='1' AND E( 1)='0' AND D( 8)='0' )then
          cVar2S19S54P006P066P069nsss(0) <='1';
          else
          cVar2S19S54P006P066P069nsss(0) <='0';
          end if;
        if(cVar1S20S54P018N015P019P007(0)='1' AND  A(16)='0' AND B( 3)='1' AND E( 9)='0' )then
          cVar2S20S54N006P033P067nsss(0) <='1';
          else
          cVar2S20S54N006P033P067nsss(0) <='0';
          end if;
        if(cVar1S21S54P018N015P019P007(0)='1' AND  B( 7)='1' )then
          cVar2S21S54P025nsss(0) <='1';
          else
          cVar2S21S54P025nsss(0) <='0';
          end if;
        if(cVar1S22S54P018N015P019P007(0)='1' AND  B( 7)='0' AND B(12)='0' AND A(13)='1' )then
          cVar2S22S54N025P034P012nsss(0) <='1';
          else
          cVar2S22S54N025P034P012nsss(0) <='0';
          end if;
        if(cVar1S23S54P018N015P019P059(0)='1' AND  A( 3)='1' )then
          cVar2S23S54P013nsss(0) <='1';
          else
          cVar2S23S54P013nsss(0) <='0';
          end if;
        if(cVar1S24S54P018N015P019P059(0)='1' AND  A( 3)='0' AND A(12)='1' )then
          cVar2S24S54N013P014nsss(0) <='1';
          else
          cVar2S24S54N013P014nsss(0) <='0';
          end if;
        if(cVar1S25S54P018N015P019N059(0)='1' AND  A( 6)='1' AND A( 4)='0' AND E( 1)='0' )then
          cVar2S25S54P007P011P066nsss(0) <='1';
          else
          cVar2S25S54P007P011P066nsss(0) <='0';
          end if;
        if(cVar1S26S54P018N015P019N059(0)='1' AND  A( 6)='0' AND B( 9)='1' )then
          cVar2S26S54N007P021nsss(0) <='1';
          else
          cVar2S26S54N007P021nsss(0) <='0';
          end if;
        if(cVar1S1S55P040N002P015P021(0)='1' AND  A( 8)='1' )then
          cVar2S1S55P003nsss(0) <='1';
          else
          cVar2S1S55P003nsss(0) <='0';
          end if;
        if(cVar1S2S55P040N002P015P021(0)='1' AND  A( 8)='0' AND A( 7)='1' AND B(10)='1' )then
          cVar2S2S55N003P005P038nsss(0) <='1';
          else
          cVar2S2S55N003P005P038nsss(0) <='0';
          end if;
        if(cVar1S3S55P040N002P015N021(0)='1' AND  A(17)='1' )then
          cVar2S3S55P004nsss(0) <='1';
          else
          cVar2S3S55P004nsss(0) <='0';
          end if;
        if(cVar1S4S55P040N002P015N021(0)='1' AND  A(17)='0' AND E( 5)='1' )then
          cVar2S4S55N004P050nsss(0) <='1';
          else
          cVar2S4S55N004P050nsss(0) <='0';
          end if;
        if(cVar1S5S55P040N002P015N021(0)='1' AND  A(17)='0' AND E( 5)='0' AND D( 0)='0' )then
          cVar2S5S55N004N050P068nsss(0) <='1';
          else
          cVar2S5S55N004N050P068nsss(0) <='0';
          end if;
        if(cVar1S7S55P040N002P015N013(0)='1' AND  A( 0)='1' )then
          cVar2S7S55P019nsss(0) <='1';
          else
          cVar2S7S55P019nsss(0) <='0';
          end if;
        if(cVar1S8S55N040P045P005P068(0)='1' AND  A(13)='0' )then
          cVar2S8S55P012nsss(0) <='1';
          else
          cVar2S8S55P012nsss(0) <='0';
          end if;
        if(cVar1S9S55N040P045N005P004(0)='1' AND  A( 3)='0' AND B(18)='1' )then
          cVar2S9S55P013P022nsss(0) <='1';
          else
          cVar2S9S55P013P022nsss(0) <='0';
          end if;
        if(cVar1S10S55N040P045N005P004(0)='1' AND  A( 3)='0' AND B(18)='0' AND E(15)='1' )then
          cVar2S10S55P013N022P043nsss(0) <='1';
          else
          cVar2S10S55P013N022P043nsss(0) <='0';
          end if;
        if(cVar1S11S55N040P045N005N004(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S11S55P006P024nsss(0) <='1';
          else
          cVar2S11S55P006P024nsss(0) <='0';
          end if;
        if(cVar1S12S55N040P045N005N004(0)='1' AND  A(16)='1' AND B(17)='0' AND B(18)='1' )then
          cVar2S12S55P006N024P022nsss(0) <='1';
          else
          cVar2S12S55P006N024P022nsss(0) <='0';
          end if;
        if(cVar1S13S55N040P045N005N004(0)='1' AND  A(16)='0' AND A( 6)='1' AND D( 0)='0' )then
          cVar2S13S55N006P007P068nsss(0) <='1';
          else
          cVar2S13S55N006P007P068nsss(0) <='0';
          end if;
        if(cVar1S14S55N040P045N005N004(0)='1' AND  A(16)='0' AND A( 6)='0' AND E(13)='1' )then
          cVar2S14S55N006N007P051nsss(0) <='1';
          else
          cVar2S14S55N006N007P051nsss(0) <='0';
          end if;
        if(cVar1S15S55N040N045P015P047(0)='1' AND  E( 7)='0' AND B(13)='1' AND B( 3)='0' )then
          cVar2S15S55P042P032P033nsss(0) <='1';
          else
          cVar2S15S55P042P032P033nsss(0) <='0';
          end if;
        if(cVar1S16S55N040N045P015P047(0)='1' AND  E( 7)='0' AND B(13)='0' )then
          cVar2S16S55P042N032psss(0) <='1';
          else
          cVar2S16S55P042N032psss(0) <='0';
          end if;
        if(cVar1S17S55N040N045P015P047(0)='1' AND  E( 7)='1' AND A(11)='1' AND D( 6)='1' )then
          cVar2S17S55P042P016P044nsss(0) <='1';
          else
          cVar2S17S55P042P016P044nsss(0) <='0';
          end if;
        if(cVar1S18S55N040N045P015P047(0)='1' AND  E( 7)='1' AND A(11)='0' AND B( 8)='1' )then
          cVar2S18S55P042N016P023nsss(0) <='1';
          else
          cVar2S18S55P042N016P023nsss(0) <='0';
          end if;
        if(cVar1S19S55N040N045P015P047(0)='1' AND  B( 3)='0' AND D(13)='1' AND B( 1)='1' )then
          cVar2S19S55P033P049P037nsss(0) <='1';
          else
          cVar2S19S55P033P049P037nsss(0) <='0';
          end if;
        if(cVar1S20S55N040N045N015P028(0)='1' AND  B( 5)='0' AND B( 4)='0' )then
          cVar2S20S55P029P031nsss(0) <='1';
          else
          cVar2S20S55P029P031nsss(0) <='0';
          end if;
        if(cVar1S21S55N040N045N015P028(0)='1' AND  B( 5)='1' AND A( 4)='1' )then
          cVar2S21S55P029P011nsss(0) <='1';
          else
          cVar2S21S55P029P011nsss(0) <='0';
          end if;
        if(cVar1S22S55N040N045N015N028(0)='1' AND  B( 7)='1' AND E( 6)='1' AND E( 1)='0' )then
          cVar2S22S55P025P046P066nsss(0) <='1';
          else
          cVar2S22S55P025P046P066nsss(0) <='0';
          end if;
        if(cVar1S23S55N040N045N015N028(0)='1' AND  B( 7)='1' AND E( 6)='0' AND A( 6)='1' )then
          cVar2S23S55P025N046P007nsss(0) <='1';
          else
          cVar2S23S55P025N046P007nsss(0) <='0';
          end if;
        if(cVar1S24S55N040N045N015N028(0)='1' AND  B( 7)='0' AND A(10)='1' AND A( 0)='0' )then
          cVar2S24S55N025P018P019nsss(0) <='1';
          else
          cVar2S24S55N025P018P019nsss(0) <='0';
          end if;
        if(cVar1S25S55N040N045N015N028(0)='1' AND  B( 7)='0' AND A(10)='0' AND A( 4)='1' )then
          cVar2S25S55N025N018P011nsss(0) <='1';
          else
          cVar2S25S55N025N018P011nsss(0) <='0';
          end if;
        if(cVar1S2S56P045N005N004P006(0)='1' AND  B(17)='1' )then
          cVar2S2S56P024nsss(0) <='1';
          else
          cVar2S2S56P024nsss(0) <='0';
          end if;
        if(cVar1S3S56P045N005N004P006(0)='1' AND  B(17)='0' AND B(18)='1' )then
          cVar2S3S56N024P022nsss(0) <='1';
          else
          cVar2S3S56N024P022nsss(0) <='0';
          end if;
        if(cVar1S4S56P045N005N004N006(0)='1' AND  A( 6)='1' AND D( 0)='0' )then
          cVar2S4S56P007P068nsss(0) <='1';
          else
          cVar2S4S56P007P068nsss(0) <='0';
          end if;
        if(cVar1S5S56P045N005N004N006(0)='1' AND  A( 6)='0' AND A( 8)='1' AND E(15)='1' )then
          cVar2S5S56N007P003P043nsss(0) <='1';
          else
          cVar2S5S56N007P003P043nsss(0) <='0';
          end if;
        if(cVar1S6S56P045N005N004N006(0)='1' AND  A( 6)='0' AND A( 8)='0' AND D( 5)='1' )then
          cVar2S6S56N007N003P048nsss(0) <='1';
          else
          cVar2S6S56N007N003P048nsss(0) <='0';
          end if;
        if(cVar1S8S56N045P040P021N002(0)='1' AND  A( 2)='0' AND A(11)='0' )then
          cVar2S8S56P015P016nsss(0) <='1';
          else
          cVar2S8S56P015P016nsss(0) <='0';
          end if;
        if(cVar1S9S56N045P040N021P066(0)='1' AND  B(19)='1' )then
          cVar2S9S56P020nsss(0) <='1';
          else
          cVar2S9S56P020nsss(0) <='0';
          end if;
        if(cVar1S10S56N045P040N021P066(0)='1' AND  B(19)='0' AND A(15)='0' )then
          cVar2S10S56N020P008nsss(0) <='1';
          else
          cVar2S10S56N020P008nsss(0) <='0';
          end if;
        if(cVar1S11S56N045N040P018P043(0)='1' AND  A( 2)='0' AND A( 8)='0' )then
          cVar2S11S56P015P003nsss(0) <='1';
          else
          cVar2S11S56P015P003nsss(0) <='0';
          end if;
        if(cVar1S12S56N045N040P018P043(0)='1' AND  A( 2)='0' AND A( 8)='1' AND B( 0)='1' )then
          cVar2S12S56P015P003P039nsss(0) <='1';
          else
          cVar2S12S56P015P003P039nsss(0) <='0';
          end if;
        if(cVar1S13S56N045N040P018P043(0)='1' AND  A( 2)='1' AND A(11)='0' AND B( 2)='1' )then
          cVar2S13S56P015P016P035nsss(0) <='1';
          else
          cVar2S13S56P015P016P035nsss(0) <='0';
          end if;
        if(cVar1S14S56N045N040P018P043(0)='1' AND  D(15)='1' )then
          cVar2S14S56P041nsss(0) <='1';
          else
          cVar2S14S56P041nsss(0) <='0';
          end if;
        if(cVar1S15S56N045N040P018P043(0)='1' AND  D(15)='0' AND A( 4)='1' )then
          cVar2S15S56N041P011nsss(0) <='1';
          else
          cVar2S15S56N041P011nsss(0) <='0';
          end if;
        if(cVar1S16S56N045N040P018P043(0)='1' AND  D(15)='0' AND A( 4)='0' AND D(13)='1' )then
          cVar2S16S56N041N011P049nsss(0) <='1';
          else
          cVar2S16S56N041N011P049nsss(0) <='0';
          end if;
        if(cVar1S17S56N045N040P018P060(0)='1' AND  A( 4)='0' AND B( 5)='1' AND A( 3)='1' )then
          cVar2S17S56P011P029P013nsss(0) <='1';
          else
          cVar2S17S56P011P029P013nsss(0) <='0';
          end if;
        if(cVar1S18S56N045N040P018P060(0)='1' AND  A( 4)='1' AND B( 5)='1' AND D( 4)='0' )then
          cVar2S18S56P011P029P052nsss(0) <='1';
          else
          cVar2S18S56P011P029P052nsss(0) <='0';
          end if;
        if(cVar1S19S56N045N040P018P060(0)='1' AND  A( 4)='1' AND B( 5)='0' AND A( 8)='1' )then
          cVar2S19S56P011N029P003nsss(0) <='1';
          else
          cVar2S19S56P011N029P003nsss(0) <='0';
          end if;
        if(cVar1S20S56N045N040P018P060(0)='1' AND  B(16)='0' AND B( 2)='1' AND E( 3)='0' )then
          cVar2S20S56P026P035P058nsss(0) <='1';
          else
          cVar2S20S56P026P035P058nsss(0) <='0';
          end if;
        if(cVar1S21S56N045N040P018P060(0)='1' AND  B(16)='0' AND B( 2)='0' AND A( 3)='1' )then
          cVar2S21S56P026N035P013nsss(0) <='1';
          else
          cVar2S21S56P026N035P013nsss(0) <='0';
          end if;
        if(cVar1S2S57P045N005N004P006(0)='1' AND  B(17)='1' )then
          cVar2S2S57P024nsss(0) <='1';
          else
          cVar2S2S57P024nsss(0) <='0';
          end if;
        if(cVar1S3S57P045N005N004P006(0)='1' AND  B(17)='0' AND B(18)='1' )then
          cVar2S3S57N024P022nsss(0) <='1';
          else
          cVar2S3S57N024P022nsss(0) <='0';
          end if;
        if(cVar1S4S57P045N005N004N006(0)='1' AND  A( 6)='1' AND D( 0)='0' )then
          cVar2S4S57P007P068nsss(0) <='1';
          else
          cVar2S4S57P007P068nsss(0) <='0';
          end if;
        if(cVar1S5S57P045N005N004N006(0)='1' AND  A( 6)='0' AND A(12)='1' AND E(15)='0' )then
          cVar2S5S57N007P014P043nsss(0) <='1';
          else
          cVar2S5S57N007P014P043nsss(0) <='0';
          end if;
        if(cVar1S6S57P045N005N004N006(0)='1' AND  A( 6)='0' AND A(12)='0' AND E(13)='1' )then
          cVar2S6S57N007N014P051nsss(0) <='1';
          else
          cVar2S6S57N007N014P051nsss(0) <='0';
          end if;
        if(cVar1S8S57N045P040P021N002(0)='1' AND  A( 8)='1' )then
          cVar2S8S57P003nsss(0) <='1';
          else
          cVar2S8S57P003nsss(0) <='0';
          end if;
        if(cVar1S9S57N045P040P021N002(0)='1' AND  A( 8)='0' AND A(17)='1' )then
          cVar2S9S57N003P004nsss(0) <='1';
          else
          cVar2S9S57N003P004nsss(0) <='0';
          end if;
        if(cVar1S10S57N045P040P021N002(0)='1' AND  A( 8)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S10S57N003N004P005nsss(0) <='1';
          else
          cVar2S10S57N003N004P005nsss(0) <='0';
          end if;
        if(cVar1S11S57N045P040N021P020(0)='1' AND  A(18)='1' )then
          cVar2S11S57P002nsss(0) <='1';
          else
          cVar2S11S57P002nsss(0) <='0';
          end if;
        if(cVar1S12S57N045P040N021N020(0)='1' AND  A(15)='0' AND D( 2)='1' )then
          cVar2S12S57P008P060nsss(0) <='1';
          else
          cVar2S12S57P008P060nsss(0) <='0';
          end if;
        if(cVar1S13S57N045P040N021N020(0)='1' AND  A(15)='0' AND D( 2)='0' AND B( 8)='1' )then
          cVar2S13S57P008N060P023nsss(0) <='1';
          else
          cVar2S13S57P008N060P023nsss(0) <='0';
          end if;
        if(cVar1S14S57N045N040P018P060(0)='1' AND  A( 4)='0' AND B( 5)='0' AND E( 7)='0' )then
          cVar2S14S57P011P029P042nsss(0) <='1';
          else
          cVar2S14S57P011P029P042nsss(0) <='0';
          end if;
        if(cVar1S15S57N045N040P018P060(0)='1' AND  A( 4)='0' AND B( 5)='1' AND A( 3)='1' )then
          cVar2S15S57P011P029P013nsss(0) <='1';
          else
          cVar2S15S57P011P029P013nsss(0) <='0';
          end if;
        if(cVar1S16S57N045N040P018P060(0)='1' AND  A( 4)='1' AND D(12)='1' )then
          cVar2S16S57P011P053nsss(0) <='1';
          else
          cVar2S16S57P011P053nsss(0) <='0';
          end if;
        if(cVar1S17S57N045N040P018P060(0)='1' AND  A( 4)='1' AND D(12)='0' AND E( 4)='1' )then
          cVar2S17S57P011N053P054nsss(0) <='1';
          else
          cVar2S17S57P011N053P054nsss(0) <='0';
          end if;
        if(cVar1S18S57N045N040P018P060(0)='1' AND  A( 9)='0' AND A( 1)='1' AND A( 8)='1' )then
          cVar2S18S57P001P017P003nsss(0) <='1';
          else
          cVar2S18S57P001P017P003nsss(0) <='0';
          end if;
        if(cVar1S19S57N045N040P018P060(0)='1' AND  A( 9)='0' AND A( 1)='0' AND A(11)='1' )then
          cVar2S19S57P001N017P016nsss(0) <='1';
          else
          cVar2S19S57P001N017P016nsss(0) <='0';
          end if;
        if(cVar1S20S57N045N040N018P043(0)='1' AND  A(15)='1' AND D(13)='1' )then
          cVar2S20S57P008P049nsss(0) <='1';
          else
          cVar2S20S57P008P049nsss(0) <='0';
          end if;
        if(cVar1S21S57N045N040N018P043(0)='1' AND  A(15)='1' AND D(13)='0' AND D( 1)='0' )then
          cVar2S21S57P008N049P064nsss(0) <='1';
          else
          cVar2S21S57P008N049P064nsss(0) <='0';
          end if;
        if(cVar1S22S57N045N040N018P043(0)='1' AND  A(15)='0' AND B( 9)='1' AND A( 8)='1' )then
          cVar2S22S57N008P021P003nsss(0) <='1';
          else
          cVar2S22S57N008P021P003nsss(0) <='0';
          end if;
        if(cVar1S23S57N045N040N018P043(0)='1' AND  D(15)='1' )then
          cVar2S23S57P041nsss(0) <='1';
          else
          cVar2S23S57P041nsss(0) <='0';
          end if;
        if(cVar1S24S57N045N040N018P043(0)='1' AND  D(15)='0' AND D(13)='1' )then
          cVar2S24S57N041P049nsss(0) <='1';
          else
          cVar2S24S57N041P049nsss(0) <='0';
          end if;
        if(cVar1S1S58P045N005P021P006(0)='1' AND  A(15)='0' )then
          cVar2S1S58P008nsss(0) <='1';
          else
          cVar2S1S58P008nsss(0) <='0';
          end if;
        if(cVar1S2S58P045N005P021N006(0)='1' AND  A(17)='1' AND A(10)='0' )then
          cVar2S2S58P004P018nsss(0) <='1';
          else
          cVar2S2S58P004P018nsss(0) <='0';
          end if;
        if(cVar1S3S58P045N005P021N006(0)='1' AND  A(17)='0' AND A( 6)='1' AND D( 0)='0' )then
          cVar2S3S58N004P007P068nsss(0) <='1';
          else
          cVar2S3S58N004P007P068nsss(0) <='0';
          end if;
        if(cVar1S4S58P045N005P021N006(0)='1' AND  A(17)='0' AND A( 6)='0' AND D( 5)='1' )then
          cVar2S4S58N004N007P048nsss(0) <='1';
          else
          cVar2S4S58N004N007P048nsss(0) <='0';
          end if;
        if(cVar1S6S58N045P018P040N002(0)='1' AND  B(10)='1' AND A( 2)='0' )then
          cVar2S6S58P038P015nsss(0) <='1';
          else
          cVar2S6S58P038P015nsss(0) <='0';
          end if;
        if(cVar1S7S58N045P018P040N002(0)='1' AND  B(10)='0' AND E( 2)='1' )then
          cVar2S7S58N038P062nsss(0) <='1';
          else
          cVar2S7S58N038P062nsss(0) <='0';
          end if;
        if(cVar1S8S58N045P018P040N002(0)='1' AND  B(10)='0' AND E( 2)='0' AND B( 8)='1' )then
          cVar2S8S58N038N062P023nsss(0) <='1';
          else
          cVar2S8S58N038N062P023nsss(0) <='0';
          end if;
        if(cVar1S9S58N045P018N040P043(0)='1' AND  B( 9)='0' AND B(10)='0' AND A(13)='0' )then
          cVar2S9S58P021P038P012nsss(0) <='1';
          else
          cVar2S9S58P021P038P012nsss(0) <='0';
          end if;
        if(cVar1S10S58N045P018N040P043(0)='1' AND  B( 9)='0' AND B(10)='1' AND B( 1)='1' )then
          cVar2S10S58P021P038P037nsss(0) <='1';
          else
          cVar2S10S58P021P038P037nsss(0) <='0';
          end if;
        if(cVar1S11S58N045P018N040P043(0)='1' AND  B( 9)='1' AND A( 8)='1' )then
          cVar2S11S58P021P003nsss(0) <='1';
          else
          cVar2S11S58P021P003nsss(0) <='0';
          end if;
        if(cVar1S12S58N045P018N040P043(0)='1' AND  B( 9)='1' AND A( 8)='0' AND A(16)='1' )then
          cVar2S12S58P021N003P006nsss(0) <='1';
          else
          cVar2S12S58P021N003P006nsss(0) <='0';
          end if;
        if(cVar1S13S58N045P018N040P043(0)='1' AND  D(15)='1' AND A( 7)='1' )then
          cVar2S13S58P041P005nsss(0) <='1';
          else
          cVar2S13S58P041P005nsss(0) <='0';
          end if;
        if(cVar1S14S58N045P018N040P043(0)='1' AND  D(15)='1' AND A( 7)='0' AND B(19)='1' )then
          cVar2S14S58P041N005P020nsss(0) <='1';
          else
          cVar2S14S58P041N005P020nsss(0) <='0';
          end if;
        if(cVar1S15S58N045P018N040P043(0)='1' AND  D(15)='0' AND A( 4)='1' )then
          cVar2S15S58N041P011nsss(0) <='1';
          else
          cVar2S15S58N041P011nsss(0) <='0';
          end if;
        if(cVar1S16S58N045P018N040P043(0)='1' AND  D(15)='0' AND A( 4)='0' AND A(11)='1' )then
          cVar2S16S58N041N011P016nsss(0) <='1';
          else
          cVar2S16S58N041N011P016nsss(0) <='0';
          end if;
        if(cVar1S17S58N045P018P019P056(0)='1' AND  B( 2)='1' AND D( 9)='1' )then
          cVar2S17S58P035P065nsss(0) <='1';
          else
          cVar2S17S58P035P065nsss(0) <='0';
          end if;
        if(cVar1S18S58N045P018P019P056(0)='1' AND  B( 2)='1' AND D( 9)='0' AND D( 0)='0' )then
          cVar2S18S58P035N065P068nsss(0) <='1';
          else
          cVar2S18S58P035N065P068nsss(0) <='0';
          end if;
        if(cVar1S19S58N045P018P019P056(0)='1' AND  B( 2)='0' AND B( 0)='1' )then
          cVar2S19S58N035P039nsss(0) <='1';
          else
          cVar2S19S58N035P039nsss(0) <='0';
          end if;
        if(cVar1S20S58N045P018P019P056(0)='1' AND  B( 2)='0' AND B( 0)='0' AND B( 9)='1' )then
          cVar2S20S58N035N039P021nsss(0) <='1';
          else
          cVar2S20S58N035N039P021nsss(0) <='0';
          end if;
        if(cVar1S21S58N045P018P019P056(0)='1' AND  D( 1)='1' )then
          cVar2S21S58P064nsss(0) <='1';
          else
          cVar2S21S58P064nsss(0) <='0';
          end if;
        if(cVar1S22S58N045P018P019P056(0)='1' AND  D( 1)='0' AND E(12)='1' )then
          cVar2S22S58N064P055nsss(0) <='1';
          else
          cVar2S22S58N064P055nsss(0) <='0';
          end if;
        if(cVar1S23S58N045P018N019P024(0)='1' AND  B(15)='1' AND A( 5)='0' )then
          cVar2S23S58P028P009nsss(0) <='1';
          else
          cVar2S23S58P028P009nsss(0) <='0';
          end if;
        if(cVar1S24S58N045P018N019P024(0)='1' AND  B(15)='0' AND E(12)='1' AND A( 3)='1' )then
          cVar2S24S58N028P055P013nsss(0) <='1';
          else
          cVar2S24S58N028P055P013nsss(0) <='0';
          end if;
        if(cVar1S25S58N045P018N019P024(0)='1' AND  B(11)='0' AND A(13)='1' )then
          cVar2S25S58P036P012nsss(0) <='1';
          else
          cVar2S25S58P036P012nsss(0) <='0';
          end if;
        if(cVar1S26S58N045P018N019P024(0)='1' AND  B(11)='0' AND A(13)='0' AND D(13)='1' )then
          cVar2S26S58P036N012P049nsss(0) <='1';
          else
          cVar2S26S58P036N012P049nsss(0) <='0';
          end if;
        if(cVar1S3S59P045N022N023P006(0)='1' AND  B(17)='1' )then
          cVar2S3S59P024nsss(0) <='1';
          else
          cVar2S3S59P024nsss(0) <='0';
          end if;
        if(cVar1S4S59P045N022N023N006(0)='1' AND  D( 6)='1' )then
          cVar2S4S59P044nsss(0) <='1';
          else
          cVar2S4S59P044nsss(0) <='0';
          end if;
        if(cVar1S5S59P045N022N023N006(0)='1' AND  D( 6)='0' AND E( 9)='1' )then
          cVar2S5S59N044P067nsss(0) <='1';
          else
          cVar2S5S59N044P067nsss(0) <='0';
          end if;
        if(cVar1S6S59P045N022N023N006(0)='1' AND  D( 6)='0' AND E( 9)='0' AND A(17)='1' )then
          cVar2S6S59N044N067P004nsss(0) <='1';
          else
          cVar2S6S59N044N067P004nsss(0) <='0';
          end if;
        if(cVar1S8S59N045P040P021N002(0)='1' AND  A( 8)='1' )then
          cVar2S8S59P003nsss(0) <='1';
          else
          cVar2S8S59P003nsss(0) <='0';
          end if;
        if(cVar1S9S59N045P040P021N002(0)='1' AND  A( 8)='0' AND A(17)='1' )then
          cVar2S9S59N003P004nsss(0) <='1';
          else
          cVar2S9S59N003P004nsss(0) <='0';
          end if;
        if(cVar1S10S59N045P040P021N002(0)='1' AND  A( 8)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S10S59N003N004P005nsss(0) <='1';
          else
          cVar2S10S59N003N004P005nsss(0) <='0';
          end if;
        if(cVar1S12S59N045P040N021P066(0)='1' AND  A(10)='0' AND B( 1)='0' )then
          cVar2S12S59P018P037nsss(0) <='1';
          else
          cVar2S12S59P018P037nsss(0) <='0';
          end if;
        if(cVar1S13S59N045N040P025P007(0)='1' AND  E( 1)='0' )then
          cVar2S13S59P066nsss(0) <='1';
          else
          cVar2S13S59P066nsss(0) <='0';
          end if;
        if(cVar1S14S59N045N040P025N007(0)='1' AND  E( 6)='1' AND A(17)='1' )then
          cVar2S14S59P046P004nsss(0) <='1';
          else
          cVar2S14S59P046P004nsss(0) <='0';
          end if;
        if(cVar1S15S59N045N040P025N007(0)='1' AND  E( 6)='1' AND A(17)='0' AND A(16)='1' )then
          cVar2S15S59P046N004P006nsss(0) <='1';
          else
          cVar2S15S59P046N004P006nsss(0) <='0';
          end if;
        if(cVar1S16S59N045N040P025N007(0)='1' AND  E( 6)='0' AND A( 8)='0' AND E( 3)='1' )then
          cVar2S16S59N046P003P058nsss(0) <='1';
          else
          cVar2S16S59N046P003P058nsss(0) <='0';
          end if;
        if(cVar1S17S59N045N040N025P018(0)='1' AND  B(18)='0' AND D(11)='0' AND B(13)='0' )then
          cVar2S17S59P022P057P032nsss(0) <='1';
          else
          cVar2S17S59P022P057P032nsss(0) <='0';
          end if;
        if(cVar1S18S59N045N040N025P018(0)='1' AND  B(18)='0' AND D(11)='1' AND D( 0)='1' )then
          cVar2S18S59P022P057P068nsss(0) <='1';
          else
          cVar2S18S59P022P057P068nsss(0) <='0';
          end if;
        if(cVar1S19S59N045N040N025N018(0)='1' AND  B(14)='1' AND B( 4)='0' AND A(13)='1' )then
          cVar2S19S59P030P031P012nsss(0) <='1';
          else
          cVar2S19S59P030P031P012nsss(0) <='0';
          end if;
        if(cVar1S20S59N045N040N025N018(0)='1' AND  B(14)='0' AND D(11)='0' AND E(10)='1' )then
          cVar2S20S59N030P057P063nsss(0) <='1';
          else
          cVar2S20S59N030P057P063nsss(0) <='0';
          end if;
        if(cVar1S21S59N045N040N025N018(0)='1' AND  B(14)='0' AND D(11)='1' AND B( 4)='1' )then
          cVar2S21S59N030P057P031nsss(0) <='1';
          else
          cVar2S21S59N030P057P031nsss(0) <='0';
          end if;
        if(cVar1S1S60P045N005P021P024(0)='1' AND  A(16)='1' )then
          cVar2S1S60P006nsss(0) <='1';
          else
          cVar2S1S60P006nsss(0) <='0';
          end if;
        if(cVar1S2S60P045N005P021P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S2S60N006P004nsss(0) <='1';
          else
          cVar2S2S60N006P004nsss(0) <='0';
          end if;
        if(cVar1S3S60P045N005P021P024(0)='1' AND  A(16)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S3S60N006N004P007nsss(0) <='1';
          else
          cVar2S3S60N006N004P007nsss(0) <='0';
          end if;
        if(cVar1S5S60N045P018P040P002(0)='1' AND  B( 9)='1' )then
          cVar2S5S60P021nsss(0) <='1';
          else
          cVar2S5S60P021nsss(0) <='0';
          end if;
        if(cVar1S6S60N045P018P040P002(0)='1' AND  B( 9)='0' AND B( 0)='1' )then
          cVar2S6S60N021P039nsss(0) <='1';
          else
          cVar2S6S60N021P039nsss(0) <='0';
          end if;
        if(cVar1S7S60N045P018P040P002(0)='1' AND  B( 9)='0' AND B( 0)='0' AND B(10)='1' )then
          cVar2S7S60N021N039P038nsss(0) <='1';
          else
          cVar2S7S60N021N039P038nsss(0) <='0';
          end if;
        if(cVar1S8S60N045P018P040N002(0)='1' AND  D(13)='1' )then
          cVar2S8S60P049nsss(0) <='1';
          else
          cVar2S8S60P049nsss(0) <='0';
          end if;
        if(cVar1S9S60N045P018P040N002(0)='1' AND  D(13)='0' AND B( 9)='1' )then
          cVar2S9S60N049P021nsss(0) <='1';
          else
          cVar2S9S60N049P021nsss(0) <='0';
          end if;
        if(cVar1S10S60N045P018P040N002(0)='1' AND  D(13)='0' AND B( 9)='0' AND E( 2)='1' )then
          cVar2S10S60N049N021P062nsss(0) <='1';
          else
          cVar2S10S60N049N021P062nsss(0) <='0';
          end if;
        if(cVar1S11S60N045P018N040P043(0)='1' AND  D( 9)='0' AND B(14)='1' AND B( 4)='0' )then
          cVar2S11S60P065P030P031nsss(0) <='1';
          else
          cVar2S11S60P065P030P031nsss(0) <='0';
          end if;
        if(cVar1S12S60N045P018N040P043(0)='1' AND  D( 9)='0' AND B(14)='0' )then
          cVar2S12S60P065N030psss(0) <='1';
          else
          cVar2S12S60P065N030psss(0) <='0';
          end if;
        if(cVar1S13S60N045P018N040P043(0)='1' AND  D( 9)='1' AND E( 1)='0' AND E( 3)='0' )then
          cVar2S13S60P065P066P058nsss(0) <='1';
          else
          cVar2S13S60P065P066P058nsss(0) <='0';
          end if;
        if(cVar1S14S60N045P018N040P043(0)='1' AND  D( 9)='1' AND E( 1)='1' AND D( 8)='1' )then
          cVar2S14S60P065P066P069nsss(0) <='1';
          else
          cVar2S14S60P065P066P069nsss(0) <='0';
          end if;
        if(cVar1S15S60N045P018N040P043(0)='1' AND  D(15)='1' AND B(18)='1' )then
          cVar2S15S60P041P022nsss(0) <='1';
          else
          cVar2S15S60P041P022nsss(0) <='0';
          end if;
        if(cVar1S16S60N045P018N040P043(0)='1' AND  D(15)='1' AND B(18)='0' AND B(19)='1' )then
          cVar2S16S60P041N022P020nsss(0) <='1';
          else
          cVar2S16S60P041N022P020nsss(0) <='0';
          end if;
        if(cVar1S17S60N045P018N040P043(0)='1' AND  D(15)='0' AND D(13)='1' )then
          cVar2S17S60N041P049nsss(0) <='1';
          else
          cVar2S17S60N041P049nsss(0) <='0';
          end if;
        if(cVar1S19S60N045P018P025N035(0)='1' AND  E( 1)='0' AND E( 6)='1' )then
          cVar2S19S60P066P046nsss(0) <='1';
          else
          cVar2S19S60P066P046nsss(0) <='0';
          end if;
        if(cVar1S20S60N045P018P025N035(0)='1' AND  E( 1)='0' AND E( 6)='0' AND A(12)='0' )then
          cVar2S20S60P066N046P014nsss(0) <='1';
          else
          cVar2S20S60P066N046P014nsss(0) <='0';
          end if;
        if(cVar1S21S60N045P018N025P037(0)='1' AND  E( 1)='1' AND B(11)='1' )then
          cVar2S21S60P066P036nsss(0) <='1';
          else
          cVar2S21S60P066P036nsss(0) <='0';
          end if;
        if(cVar1S22S60N045P018N025P037(0)='1' AND  E( 1)='0' AND D( 7)='1' )then
          cVar2S22S60N066P040nsss(0) <='1';
          else
          cVar2S22S60N066P040nsss(0) <='0';
          end if;
        if(cVar1S23S60N045P018N025P037(0)='1' AND  E( 1)='0' AND A(16)='1' AND A(11)='0' )then
          cVar2S23S60P066P006P016nsss(0) <='1';
          else
          cVar2S23S60P066P006P016nsss(0) <='0';
          end if;
        if(cVar1S24S60N045P018N025P037(0)='1' AND  E( 1)='0' AND A(16)='0' AND E( 3)='1' )then
          cVar2S24S60P066N006P058nsss(0) <='1';
          else
          cVar2S24S60P066N006P058nsss(0) <='0';
          end if;
        if(cVar1S25S60N045P018N025P037(0)='1' AND  E( 1)='1' AND D(12)='1' )then
          cVar2S25S60P066P053nsss(0) <='1';
          else
          cVar2S25S60P066P053nsss(0) <='0';
          end if;
        if(cVar1S1S61P045N005P021P024(0)='1' AND  A( 3)='1' )then
          cVar2S1S61P013nsss(0) <='1';
          else
          cVar2S1S61P013nsss(0) <='0';
          end if;
        if(cVar1S2S61P045N005P021P024(0)='1' AND  A( 3)='0' AND D( 0)='0' )then
          cVar2S2S61N013P068nsss(0) <='1';
          else
          cVar2S2S61N013P068nsss(0) <='0';
          end if;
        if(cVar1S3S61P045N005P021N024(0)='1' AND  B(18)='1' )then
          cVar2S3S61P022nsss(0) <='1';
          else
          cVar2S3S61P022nsss(0) <='0';
          end if;
        if(cVar1S4S61P045N005P021N024(0)='1' AND  B(18)='0' AND D( 6)='1' )then
          cVar2S4S61N022P044nsss(0) <='1';
          else
          cVar2S4S61N022P044nsss(0) <='0';
          end if;
        if(cVar1S5S61P045N005P021N024(0)='1' AND  B(18)='0' AND D( 6)='0' AND B( 7)='1' )then
          cVar2S5S61N022N044P025nsss(0) <='1';
          else
          cVar2S5S61N022N044P025nsss(0) <='0';
          end if;
        if(cVar1S6S61N045P018P037P061(0)='1' AND  A( 1)='1' AND B(11)='0' )then
          cVar2S6S61P017P036nsss(0) <='1';
          else
          cVar2S6S61P017P036nsss(0) <='0';
          end if;
        if(cVar1S7S61N045P018P037P061(0)='1' AND  A( 1)='0' AND A( 5)='1' )then
          cVar2S7S61N017P009nsss(0) <='1';
          else
          cVar2S7S61N017P009nsss(0) <='0';
          end if;
        if(cVar1S8S61N045P018P037P061(0)='1' AND  A( 1)='0' AND A( 5)='0' AND B(11)='1' )then
          cVar2S8S61N017N009P036nsss(0) <='1';
          else
          cVar2S8S61N017N009P036nsss(0) <='0';
          end if;
        if(cVar1S9S61N045P018P037N061(0)='1' AND  E(11)='0' AND D( 0)='1' AND A(12)='0' )then
          cVar2S9S61P059P068P014nsss(0) <='1';
          else
          cVar2S9S61P059P068P014nsss(0) <='0';
          end if;
        if(cVar1S10S61N045P018P037N061(0)='1' AND  E(11)='0' AND D( 0)='0' )then
          cVar2S10S61P059N068psss(0) <='1';
          else
          cVar2S10S61P059N068psss(0) <='0';
          end if;
        if(cVar1S11S61N045P018P037N061(0)='1' AND  E(11)='1' AND E(12)='1' )then
          cVar2S11S61P059P055nsss(0) <='1';
          else
          cVar2S11S61P059P055nsss(0) <='0';
          end if;
        if(cVar1S12S61N045P018P037P066(0)='1' AND  A(16)='1' AND A(11)='0' )then
          cVar2S12S61P006P016nsss(0) <='1';
          else
          cVar2S12S61P006P016nsss(0) <='0';
          end if;
        if(cVar1S13S61N045P018P037P066(0)='1' AND  A(16)='0' AND D( 0)='0' AND E( 4)='0' )then
          cVar2S13S61N006P068P054nsss(0) <='1';
          else
          cVar2S13S61N006P068P054nsss(0) <='0';
          end if;
        if(cVar1S14S61N045P018P037P066(0)='1' AND  A(11)='1' AND A( 8)='0' )then
          cVar2S14S61P016P003nsss(0) <='1';
          else
          cVar2S14S61P016P003nsss(0) <='0';
          end if;
        if(cVar1S15S61N045P018P037P066(0)='1' AND  A(11)='0' AND B(17)='0' AND B( 4)='1' )then
          cVar2S15S61N016P024P031nsss(0) <='1';
          else
          cVar2S15S61N016P024P031nsss(0) <='0';
          end if;
        if(cVar1S17S61N045N018P040N002(0)='1' AND  D(13)='1' )then
          cVar2S17S61P049nsss(0) <='1';
          else
          cVar2S17S61P049nsss(0) <='0';
          end if;
        if(cVar1S18S61N045N018P040N002(0)='1' AND  D(13)='0' AND B(12)='0' )then
          cVar2S18S61N049P034nsss(0) <='1';
          else
          cVar2S18S61N049P034nsss(0) <='0';
          end if;
        if(cVar1S19S61N045N018N040P000(0)='1' AND  B(15)='1' AND A(14)='1' )then
          cVar2S19S61P028P010nsss(0) <='1';
          else
          cVar2S19S61P028P010nsss(0) <='0';
          end if;
        if(cVar1S20S61N045N018N040P000(0)='1' AND  B(15)='1' AND A(14)='0' AND A( 4)='1' )then
          cVar2S20S61P028N010P011nsss(0) <='1';
          else
          cVar2S20S61P028N010P011nsss(0) <='0';
          end if;
        if(cVar1S21S61N045N018N040P000(0)='1' AND  B(15)='0' AND B( 5)='1' AND A( 4)='1' )then
          cVar2S21S61N028P029P011nsss(0) <='1';
          else
          cVar2S21S61N028P029P011nsss(0) <='0';
          end if;
        if(cVar1S22S61N045N018N040P000(0)='1' AND  E(10)='0' AND D( 2)='0' AND B(11)='0' )then
          cVar2S22S61P063P060P036nsss(0) <='1';
          else
          cVar2S22S61P063P060P036nsss(0) <='0';
          end if;
        if(cVar1S1S62P045N005P027P024(0)='1' AND  A(16)='1' )then
          cVar2S1S62P006nsss(0) <='1';
          else
          cVar2S1S62P006nsss(0) <='0';
          end if;
        if(cVar1S2S62P045N005P027P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S2S62N006P004nsss(0) <='1';
          else
          cVar2S2S62N006P004nsss(0) <='0';
          end if;
        if(cVar1S3S62P045N005P027P024(0)='1' AND  A(16)='0' AND A(17)='0' AND E(14)='1' )then
          cVar2S3S62N006N004P047nsss(0) <='1';
          else
          cVar2S3S62N006N004P047nsss(0) <='0';
          end if;
        if(cVar1S4S62P045N005P027N024(0)='1' AND  A(12)='1' AND B(18)='1' )then
          cVar2S4S62P014P022nsss(0) <='1';
          else
          cVar2S4S62P014P022nsss(0) <='0';
          end if;
        if(cVar1S5S62P045N005P027N024(0)='1' AND  A(12)='1' AND B(18)='0' AND A( 3)='0' )then
          cVar2S5S62P014N022P013nsss(0) <='1';
          else
          cVar2S5S62P014N022P013nsss(0) <='0';
          end if;
        if(cVar1S6S62P045N005P027N024(0)='1' AND  A(12)='0' AND D(10)='1' )then
          cVar2S6S62N014P061nsss(0) <='1';
          else
          cVar2S6S62N014P061nsss(0) <='0';
          end if;
        if(cVar1S7S62P045N005P027N024(0)='1' AND  A(12)='0' AND D(10)='0' AND A( 8)='1' )then
          cVar2S7S62N014N061P003nsss(0) <='1';
          else
          cVar2S7S62N014N061P003nsss(0) <='0';
          end if;
        if(cVar1S8S62N045P018P000P030(0)='1' AND  B( 4)='0' AND A(13)='1' )then
          cVar2S8S62P031P012nsss(0) <='1';
          else
          cVar2S8S62P031P012nsss(0) <='0';
          end if;
        if(cVar1S9S62N045P018P000P030(0)='1' AND  B( 4)='0' AND A(13)='0' AND A(14)='1' )then
          cVar2S9S62P031N012P010nsss(0) <='1';
          else
          cVar2S9S62P031N012P010nsss(0) <='0';
          end if;
        if(cVar1S10S62N045P018P000N030(0)='1' AND  B( 4)='1' AND A( 3)='1' )then
          cVar2S10S62P031P013nsss(0) <='1';
          else
          cVar2S10S62P031P013nsss(0) <='0';
          end if;
        if(cVar1S11S62N045P018P000N030(0)='1' AND  B( 4)='1' AND A( 3)='0' AND A( 4)='1' )then
          cVar2S11S62P031N013P011nsss(0) <='1';
          else
          cVar2S11S62P031N013P011nsss(0) <='0';
          end if;
        if(cVar1S12S62N045P018P000N030(0)='1' AND  B( 4)='0' AND E( 4)='0' AND A( 4)='0' )then
          cVar2S12S62N031P054P011nsss(0) <='1';
          else
          cVar2S12S62N031P054P011nsss(0) <='0';
          end if;
        if(cVar1S13S62N045P018P000N030(0)='1' AND  B( 4)='0' AND E( 4)='1' AND B( 5)='1' )then
          cVar2S13S62N031P054P029nsss(0) <='1';
          else
          cVar2S13S62N031P054P029nsss(0) <='0';
          end if;
        if(cVar1S15S62N045P018P000N040(0)='1' AND  B( 2)='0' AND A( 3)='1' AND A( 0)='1' )then
          cVar2S15S62P035P013P019nsss(0) <='1';
          else
          cVar2S15S62P035P013P019nsss(0) <='0';
          end if;
        if(cVar1S16S62N045P018P000N040(0)='1' AND  B( 2)='0' AND A( 3)='0' AND A( 8)='1' )then
          cVar2S16S62P035N013P003nsss(0) <='1';
          else
          cVar2S16S62P035N013P003nsss(0) <='0';
          end if;
        if(cVar1S18S62N045P018P061N035(0)='1' AND  A(12)='1' AND B(12)='1' )then
          cVar2S18S62P014P034nsss(0) <='1';
          else
          cVar2S18S62P014P034nsss(0) <='0';
          end if;
        if(cVar1S19S62N045P018P061N035(0)='1' AND  A(12)='1' AND B(12)='0' AND B( 1)='0' )then
          cVar2S19S62P014N034P037nsss(0) <='1';
          else
          cVar2S19S62P014N034P037nsss(0) <='0';
          end if;
        if(cVar1S20S62N045P018P061N035(0)='1' AND  A(12)='0' AND A( 2)='1' )then
          cVar2S20S62N014P015nsss(0) <='1';
          else
          cVar2S20S62N014P015nsss(0) <='0';
          end if;
        if(cVar1S21S62N045P018N061P025(0)='1' AND  B( 2)='1' )then
          cVar2S21S62P035nsss(0) <='1';
          else
          cVar2S21S62P035nsss(0) <='0';
          end if;
        if(cVar1S22S62N045P018N061P025(0)='1' AND  B( 2)='0' AND A( 4)='0' )then
          cVar2S22S62N035P011nsss(0) <='1';
          else
          cVar2S22S62N035P011nsss(0) <='0';
          end if;
        if(cVar1S23S62N045P018N061N025(0)='1' AND  E(10)='0' AND D( 9)='1' AND E( 9)='1' )then
          cVar2S23S62P063P065P067nsss(0) <='1';
          else
          cVar2S23S62P063P065P067nsss(0) <='0';
          end if;
        if(cVar1S24S62N045P018N061N025(0)='1' AND  E(10)='0' AND D( 9)='0' AND A(16)='1' )then
          cVar2S24S62P063N065P006nsss(0) <='1';
          else
          cVar2S24S62P063N065P006nsss(0) <='0';
          end if;
        if(cVar1S1S63P045N005P021P007(0)='1' AND  D( 0)='0' )then
          cVar2S1S63P068nsss(0) <='1';
          else
          cVar2S1S63P068nsss(0) <='0';
          end if;
        if(cVar1S2S63P045N005P021N007(0)='1' AND  A(16)='1' AND A(17)='0' )then
          cVar2S2S63P006P004nsss(0) <='1';
          else
          cVar2S2S63P006P004nsss(0) <='0';
          end if;
        if(cVar1S3S63P045N005P021N007(0)='1' AND  A(16)='0' AND A(17)='1' AND A(10)='0' )then
          cVar2S3S63N006P004P018nsss(0) <='1';
          else
          cVar2S3S63N006P004P018nsss(0) <='0';
          end if;
        if(cVar1S4S63P045N005P021N007(0)='1' AND  A(16)='0' AND A(17)='0' )then
          cVar2S4S63N006N004psss(0) <='1';
          else
          cVar2S4S63N006N004psss(0) <='0';
          end if;
        if(cVar1S5S63N045P018P019P056(0)='1' AND  B( 3)='0' AND B( 6)='1' AND E( 1)='0' )then
          cVar2S5S63P033P027P066nsss(0) <='1';
          else
          cVar2S5S63P033P027P066nsss(0) <='0';
          end if;
        if(cVar1S6S63N045P018P019P056(0)='1' AND  B( 3)='0' AND B( 6)='0' )then
          cVar2S6S63P033N027psss(0) <='1';
          else
          cVar2S6S63P033N027psss(0) <='0';
          end if;
        if(cVar1S7S63N045P018P019P056(0)='1' AND  B( 3)='1' AND E(11)='1' )then
          cVar2S7S63P033P059nsss(0) <='1';
          else
          cVar2S7S63P033P059nsss(0) <='0';
          end if;
        if(cVar1S8S63N045P018P019P056(0)='1' AND  B( 3)='1' AND E(11)='0' AND B(11)='1' )then
          cVar2S8S63P033N059P036nsss(0) <='1';
          else
          cVar2S8S63P033N059P036nsss(0) <='0';
          end if;
        if(cVar1S9S63N045P018P019P056(0)='1' AND  D( 1)='1' )then
          cVar2S9S63P064nsss(0) <='1';
          else
          cVar2S9S63P064nsss(0) <='0';
          end if;
        if(cVar1S10S63N045P018P019P056(0)='1' AND  D( 1)='0' AND A( 3)='1' AND B( 4)='1' )then
          cVar2S10S63N064P013P031nsss(0) <='1';
          else
          cVar2S10S63N064P013P031nsss(0) <='0';
          end if;
        if(cVar1S11S63N045P018P019P056(0)='1' AND  D( 1)='0' AND A( 3)='0' AND B(14)='1' )then
          cVar2S11S63N064N013P030nsss(0) <='1';
          else
          cVar2S11S63N064N013P030nsss(0) <='0';
          end if;
        if(cVar1S12S63N045P018N019P024(0)='1' AND  A( 6)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar2S12S63P007P031P013nsss(0) <='1';
          else
          cVar2S12S63P007P031P013nsss(0) <='0';
          end if;
        if(cVar1S13S63N045P018N019P024(0)='1' AND  A( 6)='0' AND B( 4)='0' AND A(17)='0' )then
          cVar2S13S63P007N031P004nsss(0) <='1';
          else
          cVar2S13S63P007N031P004nsss(0) <='0';
          end if;
        if(cVar1S14S63N045P018N019P024(0)='1' AND  A( 6)='1' AND D(13)='1' )then
          cVar2S14S63P007P049nsss(0) <='1';
          else
          cVar2S14S63P007P049nsss(0) <='0';
          end if;
        if(cVar1S15S63N045P018N019P024(0)='1' AND  A( 6)='1' AND D(13)='0' AND B( 7)='1' )then
          cVar2S15S63P007N049P025nsss(0) <='1';
          else
          cVar2S15S63P007N049P025nsss(0) <='0';
          end if;
        if(cVar1S16S63N045P018N019P024(0)='1' AND  B(11)='0' AND A(12)='1' )then
          cVar2S16S63P036P014nsss(0) <='1';
          else
          cVar2S16S63P036P014nsss(0) <='0';
          end if;
        if(cVar1S17S63N045N018P030P031(0)='1' AND  B( 2)='0' AND E(10)='0' )then
          cVar2S17S63P035P063nsss(0) <='1';
          else
          cVar2S17S63P035P063nsss(0) <='0';
          end if;
        if(cVar1S18S63N045N018P030P031(0)='1' AND  B( 2)='1' AND A( 4)='0' AND A( 0)='1' )then
          cVar2S18S63P035P011P019nsss(0) <='1';
          else
          cVar2S18S63P035P011P019nsss(0) <='0';
          end if;
        if(cVar1S19S63N045N018N030P031(0)='1' AND  A( 3)='1' )then
          cVar2S19S63P013nsss(0) <='1';
          else
          cVar2S19S63P013nsss(0) <='0';
          end if;
        if(cVar1S20S63N045N018N030P031(0)='1' AND  A( 3)='0' AND A( 4)='1' AND A(11)='0' )then
          cVar2S20S63N013P011P016nsss(0) <='1';
          else
          cVar2S20S63N013P011P016nsss(0) <='0';
          end if;
        if(cVar1S21S63N045N018N030P031(0)='1' AND  A( 3)='0' AND A( 4)='0' AND A(13)='1' )then
          cVar2S21S63N013N011P012nsss(0) <='1';
          else
          cVar2S21S63N013N011P012nsss(0) <='0';
          end if;
        if(cVar1S22S63N045N018N030N031(0)='1' AND  D(11)='0' AND A(12)='1' AND D( 2)='1' )then
          cVar2S22S63P057P014P060nsss(0) <='1';
          else
          cVar2S22S63P057P014P060nsss(0) <='0';
          end if;
        if(cVar1S23S63N045N018N030N031(0)='1' AND  D(11)='0' AND A(12)='0' AND D( 8)='1' )then
          cVar2S23S63P057N014P069nsss(0) <='1';
          else
          cVar2S23S63P057N014P069nsss(0) <='0';
          end if;
        if(cVar1S24S63N045N018N030N031(0)='1' AND  D(11)='1' AND B(15)='1' AND A(14)='1' )then
          cVar2S24S63P057P028P010nsss(0) <='1';
          else
          cVar2S24S63P057P028P010nsss(0) <='0';
          end if;
        if(cVar1S25S63N045N018N030N031(0)='1' AND  D(11)='1' AND B(15)='0' AND D( 2)='1' )then
          cVar2S25S63P057N028P060nsss(0) <='1';
          else
          cVar2S25S63P057N028P060nsss(0) <='0';
          end if;
        if(cVar1S0S64P018P069P011P029(0)='1' AND  D(12)='1' )then
          cVar2S0S64P053nsss(0) <='1';
          else
          cVar2S0S64P053nsss(0) <='0';
          end if;
        if(cVar1S1S64P018P069P011P029(0)='1' AND  D(12)='0' AND E( 4)='1' AND D(11)='0' )then
          cVar2S1S64N053P054P057nsss(0) <='1';
          else
          cVar2S1S64N053P054P057nsss(0) <='0';
          end if;
        if(cVar1S2S64P018P069P011P029(0)='1' AND  D(12)='0' AND E( 4)='0' AND D( 4)='1' )then
          cVar2S2S64N053N054P052nsss(0) <='1';
          else
          cVar2S2S64N053N054P052nsss(0) <='0';
          end if;
        if(cVar1S3S64P018P069P011N029(0)='1' AND  B(19)='1' )then
          cVar2S3S64P020nsss(0) <='1';
          else
          cVar2S3S64P020nsss(0) <='0';
          end if;
        if(cVar1S4S64P018P069P011N029(0)='1' AND  B(19)='0' AND A(12)='1' AND D( 3)='0' )then
          cVar2S4S64N020P014P056nsss(0) <='1';
          else
          cVar2S4S64N020P014P056nsss(0) <='0';
          end if;
        if(cVar1S5S64P018P069P011N029(0)='1' AND  B(19)='0' AND A(12)='0' AND E(10)='0' )then
          cVar2S5S64N020N014P063nsss(0) <='1';
          else
          cVar2S5S64N020N014P063nsss(0) <='0';
          end if;
        if(cVar1S6S64P018P069N011P029(0)='1' AND  D(14)='1' AND A(17)='1' AND A(16)='0' )then
          cVar2S6S64P045P004P006nsss(0) <='1';
          else
          cVar2S6S64P045P004P006nsss(0) <='0';
          end if;
        if(cVar1S7S64P018P069N011P029(0)='1' AND  D(14)='1' AND A(17)='0' )then
          cVar2S7S64P045N004psss(0) <='1';
          else
          cVar2S7S64P045N004psss(0) <='0';
          end if;
        if(cVar1S8S64P018P069N011P029(0)='1' AND  D(14)='0' AND D(15)='1' AND B(19)='1' )then
          cVar2S8S64N045P041P020nsss(0) <='1';
          else
          cVar2S8S64N045P041P020nsss(0) <='0';
          end if;
        if(cVar1S9S64P018P069N011P029(0)='1' AND  D(14)='0' AND D(15)='0' AND E(15)='0' )then
          cVar2S9S64N045N041P043nsss(0) <='1';
          else
          cVar2S9S64N045N041P043nsss(0) <='0';
          end if;
        if(cVar1S10S64P018P069N011P029(0)='1' AND  A( 5)='1' )then
          cVar2S10S64P009nsss(0) <='1';
          else
          cVar2S10S64P009nsss(0) <='0';
          end if;
        if(cVar1S11S64P018P069N011P029(0)='1' AND  A( 5)='0' AND A(14)='1' AND A( 0)='0' )then
          cVar2S11S64N009P010P019nsss(0) <='1';
          else
          cVar2S11S64N009P010P019nsss(0) <='0';
          end if;
        if(cVar1S12S64P018P069P019P067(0)='1' AND  D( 9)='1' )then
          cVar2S12S64P065nsss(0) <='1';
          else
          cVar2S12S64P065nsss(0) <='0';
          end if;
        if(cVar1S13S64P018P069P019P067(0)='1' AND  D( 9)='0' AND A( 1)='0' AND A( 3)='0' )then
          cVar2S13S64N065P017P013nsss(0) <='1';
          else
          cVar2S13S64N065P017P013nsss(0) <='0';
          end if;
        if(cVar1S14S64P018P069P019P067(0)='1' AND  D( 9)='0' AND A( 1)='1' AND B(11)='0' )then
          cVar2S14S64N065P017P036nsss(0) <='1';
          else
          cVar2S14S64N065P017P036nsss(0) <='0';
          end if;
        if(cVar1S15S64P018P069P019N067(0)='1' AND  E( 1)='1' AND B( 1)='0' )then
          cVar2S15S64P066P037nsss(0) <='1';
          else
          cVar2S15S64P066P037nsss(0) <='0';
          end if;
        if(cVar1S16S64P018P069N019P068(0)='1' AND  E(11)='1' )then
          cVar2S16S64P059nsss(0) <='1';
          else
          cVar2S16S64P059nsss(0) <='0';
          end if;
        if(cVar1S17S64P018P069N019P068(0)='1' AND  E(11)='0' AND D( 9)='0' )then
          cVar2S17S64N059P065nsss(0) <='1';
          else
          cVar2S17S64N059P065nsss(0) <='0';
          end if;
        if(cVar1S18S64P018P069N019N068(0)='1' AND  B( 2)='0' AND E( 9)='0' AND D( 4)='0' )then
          cVar2S18S64P035P067P052nsss(0) <='1';
          else
          cVar2S18S64P035P067P052nsss(0) <='0';
          end if;
        if(cVar1S19S64P018P069N019N068(0)='1' AND  B( 2)='1' AND A( 1)='1' AND D( 1)='1' )then
          cVar2S19S64P035P017P064nsss(0) <='1';
          else
          cVar2S19S64P035P017P064nsss(0) <='0';
          end if;
        if(cVar1S20S64P018P031P007P013(0)='1' AND  E( 4)='1' )then
          cVar2S20S64P054nsss(0) <='1';
          else
          cVar2S20S64P054nsss(0) <='0';
          end if;
        if(cVar1S21S64P018P031P007P013(0)='1' AND  E( 4)='0' AND D(11)='1' )then
          cVar2S21S64N054P057nsss(0) <='1';
          else
          cVar2S21S64N054P057nsss(0) <='0';
          end if;
        if(cVar1S22S64P018P031P007P013(0)='1' AND  E( 4)='0' AND D(11)='0' AND E( 3)='1' )then
          cVar2S22S64N054N057P058nsss(0) <='1';
          else
          cVar2S22S64N054N057P058nsss(0) <='0';
          end if;
        if(cVar1S23S64P018P031P007N013(0)='1' AND  D(11)='0' AND B( 1)='1' )then
          cVar2S23S64P057P037nsss(0) <='1';
          else
          cVar2S23S64P057P037nsss(0) <='0';
          end if;
        if(cVar1S24S64P018P031P007N013(0)='1' AND  D(11)='0' AND B( 1)='0' AND A(13)='1' )then
          cVar2S24S64P057N037P012nsss(0) <='1';
          else
          cVar2S24S64P057N037P012nsss(0) <='0';
          end if;
        if(cVar1S26S64P018N031P007N051(0)='1' AND  A( 3)='0' AND E(15)='1' )then
          cVar2S26S64P013P043nsss(0) <='1';
          else
          cVar2S26S64P013P043nsss(0) <='0';
          end if;
        if(cVar1S27S64P018N031P007N051(0)='1' AND  A( 3)='0' AND E(15)='0' AND B(12)='0' )then
          cVar2S27S64P013N043P034nsss(0) <='1';
          else
          cVar2S27S64P013N043P034nsss(0) <='0';
          end if;
        if(cVar1S28S64P018N031P007N051(0)='1' AND  A( 3)='1' AND D( 0)='1' )then
          cVar2S28S64P013P068nsss(0) <='1';
          else
          cVar2S28S64P013P068nsss(0) <='0';
          end if;
        if(cVar1S29S64P018N031N007P009(0)='1' AND  D( 0)='0' AND E( 2)='0' )then
          cVar2S29S64P068P062nsss(0) <='1';
          else
          cVar2S29S64P068P062nsss(0) <='0';
          end if;
        if(cVar1S30S64P018N031N007P009(0)='1' AND  D( 0)='0' AND E( 2)='1' AND B( 2)='1' )then
          cVar2S30S64P068P062P035nsss(0) <='1';
          else
          cVar2S30S64P068P062P035nsss(0) <='0';
          end if;
        if(cVar1S31S64P018N031N007N009(0)='1' AND  E( 1)='1' AND B(11)='1' AND E( 9)='0' )then
          cVar2S31S64P066P036P067nsss(0) <='1';
          else
          cVar2S31S64P066P036P067nsss(0) <='0';
          end if;
        if(cVar1S32S64P018N031N007N009(0)='1' AND  E( 1)='1' AND B(11)='0' AND B(15)='1' )then
          cVar2S32S64P066N036P028nsss(0) <='1';
          else
          cVar2S32S64P066N036P028nsss(0) <='0';
          end if;
        if(cVar1S33S64P018N031N007N009(0)='1' AND  E( 1)='0' AND B(11)='0' AND A(12)='1' )then
          cVar2S33S64N066P036P014nsss(0) <='1';
          else
          cVar2S33S64N066P036P014nsss(0) <='0';
          end if;
        if(cVar1S34S64P018N031N007N009(0)='1' AND  E( 1)='0' AND B(11)='1' AND E(11)='1' )then
          cVar2S34S64N066P036P059nsss(0) <='1';
          else
          cVar2S34S64N066P036P059nsss(0) <='0';
          end if;
        if(cVar1S0S65P018P014P042P068(0)='1' AND  B( 1)='0' AND B( 5)='0' AND A(13)='0' )then
          cVar2S0S65P037P029P012nsss(0) <='1';
          else
          cVar2S0S65P037P029P012nsss(0) <='0';
          end if;
        if(cVar1S1S65P018P014P042P068(0)='1' AND  B( 1)='1' AND B(17)='0' AND D( 3)='1' )then
          cVar2S1S65P037P024P056nsss(0) <='1';
          else
          cVar2S1S65P037P024P056nsss(0) <='0';
          end if;
        if(cVar1S2S65P018P014P042N068(0)='1' AND  A(13)='1' AND D( 9)='0' )then
          cVar2S2S65P012P065nsss(0) <='1';
          else
          cVar2S2S65P012P065nsss(0) <='0';
          end if;
        if(cVar1S3S65P018P014P042N068(0)='1' AND  A(13)='0' AND D( 3)='0' AND D( 2)='0' )then
          cVar2S3S65N012P056P060nsss(0) <='1';
          else
          cVar2S3S65N012P056P060nsss(0) <='0';
          end if;
        if(cVar1S5S65P018P014P042N004(0)='1' AND  A( 7)='1' )then
          cVar2S5S65P005nsss(0) <='1';
          else
          cVar2S5S65P005nsss(0) <='0';
          end if;
        if(cVar1S6S65P018P014P042N004(0)='1' AND  A( 7)='0' AND D( 8)='1' )then
          cVar2S6S65N005P069nsss(0) <='1';
          else
          cVar2S6S65N005P069nsss(0) <='0';
          end if;
        if(cVar1S9S65P018P014N045N046(0)='1' AND  B( 4)='1' AND B(11)='1' )then
          cVar2S9S65P031P036nsss(0) <='1';
          else
          cVar2S9S65P031P036nsss(0) <='0';
          end if;
        if(cVar1S10S65P018P014N045N046(0)='1' AND  B( 4)='1' AND B(11)='0' AND A( 0)='0' )then
          cVar2S10S65P031N036P019nsss(0) <='1';
          else
          cVar2S10S65P031N036P019nsss(0) <='0';
          end if;
        if(cVar1S11S65P018P014N045N046(0)='1' AND  B( 4)='0' AND B(13)='1' )then
          cVar2S11S65N031P032nsss(0) <='1';
          else
          cVar2S11S65N031P032nsss(0) <='0';
          end if;
        if(cVar1S12S65P018P014N045N046(0)='1' AND  B( 4)='0' AND B(13)='0' AND B(19)='1' )then
          cVar2S12S65N031N032P020nsss(0) <='1';
          else
          cVar2S12S65N031N032P020nsss(0) <='0';
          end if;
        if(cVar1S14S65N018P041P020N002(0)='1' AND  A( 8)='1' )then
          cVar2S14S65P003nsss(0) <='1';
          else
          cVar2S14S65P003nsss(0) <='0';
          end if;
        if(cVar1S15S65N018P041P020N002(0)='1' AND  A( 8)='0' AND A( 7)='1' )then
          cVar2S15S65N003P005nsss(0) <='1';
          else
          cVar2S15S65N003P005nsss(0) <='0';
          end if;
        if(cVar1S16S65N018P041N020P023(0)='1' AND  E( 7)='0' )then
          cVar2S16S65P042nsss(0) <='1';
          else
          cVar2S16S65P042nsss(0) <='0';
          end if;
        if(cVar1S17S65N018P041N020N023(0)='1' AND  A( 5)='0' AND B( 9)='1' )then
          cVar2S17S65P009P021nsss(0) <='1';
          else
          cVar2S17S65P009P021nsss(0) <='0';
          end if;
        if(cVar1S18S65N018P041N020N023(0)='1' AND  A( 5)='0' AND B( 9)='0' AND A(11)='1' )then
          cVar2S18S65P009N021P016nsss(0) <='1';
          else
          cVar2S18S65P009N021P016nsss(0) <='0';
          end if;
        if(cVar1S19S65N018N041P039P045(0)='1' AND  A(17)='1' AND A(11)='0' )then
          cVar2S19S65P004P016nsss(0) <='1';
          else
          cVar2S19S65P004P016nsss(0) <='0';
          end if;
        if(cVar1S20S65N018N041P039P045(0)='1' AND  A(17)='0' )then
          cVar2S20S65N004psss(0) <='1';
          else
          cVar2S20S65N004psss(0) <='0';
          end if;
        if(cVar1S21S65N018N041P039N045(0)='1' AND  A( 4)='1' AND B( 5)='1' AND A(14)='0' )then
          cVar2S21S65P011P029P010nsss(0) <='1';
          else
          cVar2S21S65P011P029P010nsss(0) <='0';
          end if;
        if(cVar1S22S65N018N041P039N045(0)='1' AND  A( 4)='1' AND B( 5)='0' AND A(12)='1' )then
          cVar2S22S65P011N029P014nsss(0) <='1';
          else
          cVar2S22S65P011N029P014nsss(0) <='0';
          end if;
        if(cVar1S23S65N018N041P039N045(0)='1' AND  A( 4)='0' AND B(19)='1' AND D( 7)='1' )then
          cVar2S23S65N011P020P040nsss(0) <='1';
          else
          cVar2S23S65N011P020P040nsss(0) <='0';
          end if;
        if(cVar1S25S65N018N041P039N049(0)='1' AND  A( 7)='1' )then
          cVar2S25S65P005nsss(0) <='1';
          else
          cVar2S25S65P005nsss(0) <='0';
          end if;
        if(cVar1S1S66P018P041P020N002(0)='1' AND  A( 8)='1' )then
          cVar2S1S66P003nsss(0) <='1';
          else
          cVar2S1S66P003nsss(0) <='0';
          end if;
        if(cVar1S2S66P018P041P020N002(0)='1' AND  A( 8)='0' AND A( 7)='1' )then
          cVar2S2S66N003P005nsss(0) <='1';
          else
          cVar2S2S66N003P005nsss(0) <='0';
          end if;
        if(cVar1S3S66P018P041N020P023(0)='1' AND  E( 7)='0' )then
          cVar2S3S66P042nsss(0) <='1';
          else
          cVar2S3S66P042nsss(0) <='0';
          end if;
        if(cVar1S4S66P018P041N020N023(0)='1' AND  A( 5)='0' AND B( 9)='1' )then
          cVar2S4S66P009P021nsss(0) <='1';
          else
          cVar2S4S66P009P021nsss(0) <='0';
          end if;
        if(cVar1S5S66P018P041N020N023(0)='1' AND  A( 5)='0' AND B( 9)='0' AND E(14)='1' )then
          cVar2S5S66P009N021P047nsss(0) <='1';
          else
          cVar2S5S66P009N021P047nsss(0) <='0';
          end if;
        if(cVar1S6S66P018N041P039P020(0)='1' AND  A( 5)='1' AND B( 6)='1' AND E( 1)='0' )then
          cVar2S6S66P009P027P066nsss(0) <='1';
          else
          cVar2S6S66P009P027P066nsss(0) <='0';
          end if;
        if(cVar1S7S66P018N041P039P020(0)='1' AND  A( 5)='1' AND B( 6)='0' AND D(13)='1' )then
          cVar2S7S66P009N027P049nsss(0) <='1';
          else
          cVar2S7S66P009N027P049nsss(0) <='0';
          end if;
        if(cVar1S8S66P018N041P039P020(0)='1' AND  A( 5)='0' AND B( 6)='0' AND A( 6)='0' )then
          cVar2S8S66N009P027P007nsss(0) <='1';
          else
          cVar2S8S66N009P027P007nsss(0) <='0';
          end if;
        if(cVar1S9S66P018N041P039P020(0)='1' AND  A( 5)='0' AND B( 6)='1' AND A( 6)='1' )then
          cVar2S9S66N009P027P007nsss(0) <='1';
          else
          cVar2S9S66N009P027P007nsss(0) <='0';
          end if;
        if(cVar1S10S66P018N041P039P020(0)='1' AND  A( 4)='1' )then
          cVar2S10S66P011nsss(0) <='1';
          else
          cVar2S10S66P011nsss(0) <='0';
          end if;
        if(cVar1S11S66P018N041P039P020(0)='1' AND  A( 4)='0' AND A( 6)='1' )then
          cVar2S11S66N011P007nsss(0) <='1';
          else
          cVar2S11S66N011P007nsss(0) <='0';
          end if;
        if(cVar1S12S66P018N041P039P020(0)='1' AND  A( 4)='0' AND A( 6)='0' AND D( 7)='1' )then
          cVar2S12S66N011N007P040nsss(0) <='1';
          else
          cVar2S12S66N011N007P040nsss(0) <='0';
          end if;
        if(cVar1S13S66P018N041P039P011(0)='1' AND  A( 7)='1' )then
          cVar2S13S66P005nsss(0) <='1';
          else
          cVar2S13S66P005nsss(0) <='0';
          end if;
        if(cVar1S15S66P018P068N057P063(0)='1' AND  D(15)='0' AND B(11)='1' AND B( 2)='0' )then
          cVar2S15S66P041P036P035nsss(0) <='1';
          else
          cVar2S15S66P041P036P035nsss(0) <='0';
          end if;
        if(cVar1S16S66P018P068N057P063(0)='1' AND  D(15)='0' AND B(11)='0' AND B(13)='0' )then
          cVar2S16S66P041N036P032nsss(0) <='1';
          else
          cVar2S16S66P041N036P032nsss(0) <='0';
          end if;
        if(cVar1S17S66P018P068N057P063(0)='1' AND  A( 1)='1' AND B(11)='0' )then
          cVar2S17S66P017P036nsss(0) <='1';
          else
          cVar2S17S66P017P036nsss(0) <='0';
          end if;
        if(cVar1S18S66P018P068N057P063(0)='1' AND  A( 1)='1' AND B(11)='1' AND A( 0)='1' )then
          cVar2S18S66P017P036P019nsss(0) <='1';
          else
          cVar2S18S66P017P036P019nsss(0) <='0';
          end if;
        if(cVar1S19S66P018P068N057P063(0)='1' AND  A( 1)='0' AND A(11)='1' )then
          cVar2S19S66N017P016nsss(0) <='1';
          else
          cVar2S19S66N017P016nsss(0) <='0';
          end if;
        if(cVar1S20S66P018N068P031P013(0)='1' AND  A(14)='0' )then
          cVar2S20S66P010nsss(0) <='1';
          else
          cVar2S20S66P010nsss(0) <='0';
          end if;
        if(cVar1S21S66P018N068P031N013(0)='1' AND  D(11)='0' AND A(13)='1' )then
          cVar2S21S66P057P012nsss(0) <='1';
          else
          cVar2S21S66P057P012nsss(0) <='0';
          end if;
        if(cVar1S22S66P018N068P031N013(0)='1' AND  D(11)='0' AND A(13)='0' AND A(12)='1' )then
          cVar2S22S66P057N012P014nsss(0) <='1';
          else
          cVar2S22S66P057N012P014nsss(0) <='0';
          end if;
        if(cVar1S23S66P018N068N031P005(0)='1' AND  D( 8)='0' AND E(10)='0' AND E( 6)='0' )then
          cVar2S23S66P069P063P046nsss(0) <='1';
          else
          cVar2S23S66P069P063P046nsss(0) <='0';
          end if;
        if(cVar1S24S66P018N068N031N005(0)='1' AND  A(18)='1' AND B(12)='1' )then
          cVar2S24S66P002P034nsss(0) <='1';
          else
          cVar2S24S66P002P034nsss(0) <='0';
          end if;
        if(cVar1S25S66P018N068N031N005(0)='1' AND  A(18)='1' AND B(12)='0' AND A( 3)='0' )then
          cVar2S25S66P002N034P013nsss(0) <='1';
          else
          cVar2S25S66P002N034P013nsss(0) <='0';
          end if;
        if(cVar1S26S66P018N068N031N005(0)='1' AND  A(18)='0' AND B(10)='0' AND B( 6)='1' )then
          cVar2S26S66N002P038P027nsss(0) <='1';
          else
          cVar2S26S66N002P038P027nsss(0) <='0';
          end if;
        if(cVar1S1S67P009P027P063P018(0)='1' AND  A( 0)='1' )then
          cVar2S1S67P019nsss(0) <='1';
          else
          cVar2S1S67P019nsss(0) <='0';
          end if;
        if(cVar1S2S67P009P027P063P018(0)='1' AND  A( 0)='0' AND D( 4)='0' AND D( 5)='0' )then
          cVar2S2S67N019P052P048nsss(0) <='1';
          else
          cVar2S2S67N019P052P048nsss(0) <='0';
          end if;
        if(cVar1S4S67P009N027P049N026(0)='1' AND  B( 7)='1' )then
          cVar2S4S67P025nsss(0) <='1';
          else
          cVar2S4S67P025nsss(0) <='0';
          end if;
        if(cVar1S5S67P009N027P049N026(0)='1' AND  B( 7)='0' AND B(17)='1' )then
          cVar2S5S67N025P024nsss(0) <='1';
          else
          cVar2S5S67N025P024nsss(0) <='0';
          end if;
        if(cVar1S6S67P009N027N049P014(0)='1' AND  A( 9)='1' )then
          cVar2S6S67P001nsss(0) <='1';
          else
          cVar2S6S67P001nsss(0) <='0';
          end if;
        if(cVar1S7S67P009N027N049P014(0)='1' AND  A( 9)='0' AND A(19)='0' )then
          cVar2S7S67N001P000nsss(0) <='1';
          else
          cVar2S7S67N001P000nsss(0) <='0';
          end if;
        if(cVar1S8S67P009N027N049N014(0)='1' AND  A(13)='1' AND D( 9)='1' )then
          cVar2S8S67P012P065nsss(0) <='1';
          else
          cVar2S8S67P012P065nsss(0) <='0';
          end if;
        if(cVar1S9S67P009N027N049N014(0)='1' AND  A(13)='1' AND D( 9)='0' AND A(16)='0' )then
          cVar2S9S67P012N065P006nsss(0) <='1';
          else
          cVar2S9S67P012N065P006nsss(0) <='0';
          end if;
        if(cVar1S10S67P009N027N049N014(0)='1' AND  A(13)='0' AND A( 1)='1' AND E( 5)='0' )then
          cVar2S10S67N012P017P050nsss(0) <='1';
          else
          cVar2S10S67N012P017P050nsss(0) <='0';
          end if;
        if(cVar1S13S67N009P041N020N021(0)='1' AND  A(10)='0' AND A( 6)='1' )then
          cVar2S13S67P018P007nsss(0) <='1';
          else
          cVar2S13S67P018P007nsss(0) <='0';
          end if;
        if(cVar1S14S67N009P041N020N021(0)='1' AND  A(10)='0' AND A( 6)='0' AND D( 0)='0' )then
          cVar2S14S67P018N007P068nsss(0) <='1';
          else
          cVar2S14S67P018N007P068nsss(0) <='0';
          end if;
        if(cVar1S15S67N009P041N020N021(0)='1' AND  A(10)='1' AND A(13)='0' AND E(15)='1' )then
          cVar2S15S67P018P012P043nsss(0) <='1';
          else
          cVar2S15S67P018P012P043nsss(0) <='0';
          end if;
        if(cVar1S16S67N009N041P018P000(0)='1' AND  A( 8)='0' AND B(11)='0' AND E( 9)='0' )then
          cVar2S16S67P003P036P067nsss(0) <='1';
          else
          cVar2S16S67P003P036P067nsss(0) <='0';
          end if;
        if(cVar1S17S67N009N041P018P000(0)='1' AND  A( 8)='0' AND B(11)='1' AND A( 0)='1' )then
          cVar2S17S67P003P036P019nsss(0) <='1';
          else
          cVar2S17S67P003P036P019nsss(0) <='0';
          end if;
        if(cVar1S18S67N009N041P018N000(0)='1' AND  B( 4)='1' AND A( 3)='1' AND D( 0)='0' )then
          cVar2S18S67P031P013P068nsss(0) <='1';
          else
          cVar2S18S67P031P013P068nsss(0) <='0';
          end if;
        if(cVar1S19S67N009N041P018N000(0)='1' AND  B( 4)='1' AND A( 3)='0' AND D(11)='0' )then
          cVar2S19S67P031N013P057nsss(0) <='1';
          else
          cVar2S19S67P031N013P057nsss(0) <='0';
          end if;
        if(cVar1S20S67N009N041P018N000(0)='1' AND  B( 4)='0' AND A(17)='0' AND B(10)='0' )then
          cVar2S20S67N031P004P038nsss(0) <='1';
          else
          cVar2S20S67N031P004P038nsss(0) <='0';
          end if;
        if(cVar1S21S67N009N041P018N000(0)='1' AND  B( 4)='0' AND A(17)='1' AND A( 1)='1' )then
          cVar2S21S67N031P004P017nsss(0) <='1';
          else
          cVar2S21S67N031P004P017nsss(0) <='0';
          end if;
        if(cVar1S22S67N009N041N018P039(0)='1' AND  B(19)='0' AND A( 2)='1' AND A(15)='0' )then
          cVar2S22S67P020P015P008nsss(0) <='1';
          else
          cVar2S22S67P020P015P008nsss(0) <='0';
          end if;
        if(cVar1S23S67N009N041N018P039(0)='1' AND  B(19)='0' AND A( 2)='0' AND A(11)='1' )then
          cVar2S23S67P020N015P016nsss(0) <='1';
          else
          cVar2S23S67P020N015P016nsss(0) <='0';
          end if;
        if(cVar1S24S67N009N041N018P039(0)='1' AND  B(19)='1' AND A( 0)='1' AND A( 2)='0' )then
          cVar2S24S67P020P019P015nsss(0) <='1';
          else
          cVar2S24S67P020P019P015nsss(0) <='0';
          end if;
        if(cVar1S25S67N009N041N018P039(0)='1' AND  B(19)='1' AND A( 0)='0' AND A( 4)='1' )then
          cVar2S25S67P020N019P011nsss(0) <='1';
          else
          cVar2S25S67P020N019P011nsss(0) <='0';
          end if;
        if(cVar1S26S67N009N041N018P039(0)='1' AND  A( 4)='0' AND A( 7)='1' )then
          cVar2S26S67P011P005nsss(0) <='1';
          else
          cVar2S26S67P011P005nsss(0) <='0';
          end if;
        if(cVar1S1S68P009P027P063P018(0)='1' AND  A( 0)='1' )then
          cVar2S1S68P019nsss(0) <='1';
          else
          cVar2S1S68P019nsss(0) <='0';
          end if;
        if(cVar1S3S68P009N027P049N026(0)='1' AND  B( 7)='1' )then
          cVar2S3S68P025nsss(0) <='1';
          else
          cVar2S3S68P025nsss(0) <='0';
          end if;
        if(cVar1S4S68P009N027P049N026(0)='1' AND  B( 7)='0' AND A( 0)='0' AND B(17)='1' )then
          cVar2S4S68N025P019P024nsss(0) <='1';
          else
          cVar2S4S68N025P019P024nsss(0) <='0';
          end if;
        if(cVar1S5S68P009N027N049P053(0)='1' AND  B( 5)='1' )then
          cVar2S5S68P029nsss(0) <='1';
          else
          cVar2S5S68P029nsss(0) <='0';
          end if;
        if(cVar1S6S68P009N027N049P053(0)='1' AND  B( 5)='0' AND E(13)='1' AND A( 2)='0' )then
          cVar2S6S68N029P051P015nsss(0) <='1';
          else
          cVar2S6S68N029P051P015nsss(0) <='0';
          end if;
        if(cVar1S7S68P009N027N049N053(0)='1' AND  A( 2)='1' AND D( 1)='0' AND B( 3)='0' )then
          cVar2S7S68P015P064P033nsss(0) <='1';
          else
          cVar2S7S68P015P064P033nsss(0) <='0';
          end if;
        if(cVar1S8S68P009N027N049N053(0)='1' AND  A( 2)='1' AND D( 1)='1' AND E(10)='1' )then
          cVar2S8S68P015P064P063nsss(0) <='1';
          else
          cVar2S8S68P015P064P063nsss(0) <='0';
          end if;
        if(cVar1S9S68P009N027N049N053(0)='1' AND  A( 2)='0' AND B(12)='1' )then
          cVar2S9S68N015P034nsss(0) <='1';
          else
          cVar2S9S68N015P034nsss(0) <='0';
          end if;
        if(cVar1S10S68P009N027N049N053(0)='1' AND  A( 2)='0' AND B(12)='0' AND B( 8)='1' )then
          cVar2S10S68N015N034P023nsss(0) <='1';
          else
          cVar2S10S68N015N034P023nsss(0) <='0';
          end if;
        if(cVar1S12S68N009P041P020N003(0)='1' AND  A(18)='1' )then
          cVar2S12S68P002nsss(0) <='1';
          else
          cVar2S12S68P002nsss(0) <='0';
          end if;
        if(cVar1S13S68N009P041P020N003(0)='1' AND  A(18)='0' AND A(17)='1' )then
          cVar2S13S68N002P004nsss(0) <='1';
          else
          cVar2S13S68N002P004nsss(0) <='0';
          end if;
        if(cVar1S14S68N009P041P020N003(0)='1' AND  A(18)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S14S68N002N004P005nsss(0) <='1';
          else
          cVar2S14S68N002N004P005nsss(0) <='0';
          end if;
        if(cVar1S15S68N009P041N020P021(0)='1' AND  B(10)='1' )then
          cVar2S15S68P038nsss(0) <='1';
          else
          cVar2S15S68P038nsss(0) <='0';
          end if;
        if(cVar1S16S68N009P041N020P021(0)='1' AND  B(10)='0' AND E( 7)='0' )then
          cVar2S16S68N038P042nsss(0) <='1';
          else
          cVar2S16S68N038P042nsss(0) <='0';
          end if;
        if(cVar1S17S68N009P041N020N021(0)='1' AND  A(10)='0' AND A( 6)='1' )then
          cVar2S17S68P018P007nsss(0) <='1';
          else
          cVar2S17S68P018P007nsss(0) <='0';
          end if;
        if(cVar1S18S68N009P041N020N021(0)='1' AND  A(10)='0' AND A( 6)='0' AND E(14)='1' )then
          cVar2S18S68P018N007P047nsss(0) <='1';
          else
          cVar2S18S68P018N007P047nsss(0) <='0';
          end if;
        if(cVar1S19S68N009P041N020N021(0)='1' AND  A(10)='1' AND A(13)='0' AND E(15)='1' )then
          cVar2S19S68P018P012P043nsss(0) <='1';
          else
          cVar2S19S68P018P012P043nsss(0) <='0';
          end if;
        if(cVar1S20S68N009N041P016P031(0)='1' AND  E( 4)='1' AND A( 3)='1' )then
          cVar2S20S68P054P013nsss(0) <='1';
          else
          cVar2S20S68P054P013nsss(0) <='0';
          end if;
        if(cVar1S21S68N009N041P016P031(0)='1' AND  E( 4)='1' AND A( 3)='0' AND A( 0)='0' )then
          cVar2S21S68P054N013P019nsss(0) <='1';
          else
          cVar2S21S68P054N013P019nsss(0) <='0';
          end if;
        if(cVar1S22S68N009N041P016P031(0)='1' AND  E( 4)='0' AND A( 3)='1' )then
          cVar2S22S68N054P013nsss(0) <='1';
          else
          cVar2S22S68N054P013nsss(0) <='0';
          end if;
        if(cVar1S23S68N009N041P016P031(0)='1' AND  E( 4)='0' AND A( 3)='0' AND A( 4)='1' )then
          cVar2S23S68N054N013P011nsss(0) <='1';
          else
          cVar2S23S68N054N013P011nsss(0) <='0';
          end if;
        if(cVar1S24S68N009N041P016N031(0)='1' AND  B(19)='0' AND B( 0)='0' )then
          cVar2S24S68P020P039nsss(0) <='1';
          else
          cVar2S24S68P020P039nsss(0) <='0';
          end if;
        if(cVar1S25S68N009N041P016N031(0)='1' AND  B(19)='0' AND B( 0)='1' AND D(14)='1' )then
          cVar2S25S68P020P039P045nsss(0) <='1';
          else
          cVar2S25S68P020P039P045nsss(0) <='0';
          end if;
        if(cVar1S26S68N009N041P016N031(0)='1' AND  B(19)='1' AND E( 5)='0' AND A( 8)='1' )then
          cVar2S26S68P020P050P003nsss(0) <='1';
          else
          cVar2S26S68P020P050P003nsss(0) <='0';
          end if;
        if(cVar1S27S68N009N041P016P059(0)='1' AND  B( 2)='0' AND D(12)='0' AND B(14)='1' )then
          cVar2S27S68P035P053P030nsss(0) <='1';
          else
          cVar2S27S68P035P053P030nsss(0) <='0';
          end if;
        if(cVar1S28S68N009N041P016P059(0)='1' AND  B( 2)='1' AND B( 5)='0' AND B( 1)='1' )then
          cVar2S28S68P035P029P037nsss(0) <='1';
          else
          cVar2S28S68P035P029P037nsss(0) <='0';
          end if;
        if(cVar1S29S68N009N041P016P059(0)='1' AND  A(10)='1' AND A(12)='0' )then
          cVar2S29S68P018P014nsss(0) <='1';
          else
          cVar2S29S68P018P014nsss(0) <='0';
          end if;
        if(cVar1S30S68N009N041P016P059(0)='1' AND  A(10)='1' AND A(12)='1' AND A( 1)='1' )then
          cVar2S30S68P018P014P017nsss(0) <='1';
          else
          cVar2S30S68P018P014P017nsss(0) <='0';
          end if;
        if(cVar1S31S68N009N041P016P059(0)='1' AND  A(10)='0' AND D( 8)='1' AND A( 0)='0' )then
          cVar2S31S68N018P069P019nsss(0) <='1';
          else
          cVar2S31S68N018P069P019nsss(0) <='0';
          end if;
        if(cVar1S0S69P009P049P060P067(0)='1' AND  A( 3)='0' AND E(13)='0' )then
          cVar2S0S69P013P051nsss(0) <='1';
          else
          cVar2S0S69P013P051nsss(0) <='0';
          end if;
        if(cVar1S1S69P009P049P060P067(0)='1' AND  A( 3)='0' AND E(13)='1' AND E(14)='0' )then
          cVar2S1S69P013P051P047nsss(0) <='1';
          else
          cVar2S1S69P013P051P047nsss(0) <='0';
          end if;
        if(cVar1S2S69P009P049P060P067(0)='1' AND  A( 3)='1' )then
          cVar2S2S69P013psss(0) <='1';
          else
          cVar2S2S69P013psss(0) <='0';
          end if;
        if(cVar1S4S69P009N049P053N029(0)='1' AND  E(13)='1' AND A( 6)='0' )then
          cVar2S4S69P051P007nsss(0) <='1';
          else
          cVar2S4S69P051P007nsss(0) <='0';
          end if;
        if(cVar1S5S69P009N049P053N029(0)='1' AND  E(13)='0' AND A( 0)='1' )then
          cVar2S5S69N051P019nsss(0) <='1';
          else
          cVar2S5S69N051P019nsss(0) <='0';
          end if;
        if(cVar1S6S69P009N049N053P050(0)='1' AND  B( 6)='1' AND A( 3)='0' )then
          cVar2S6S69P027P013nsss(0) <='1';
          else
          cVar2S6S69P027P013nsss(0) <='0';
          end if;
        if(cVar1S7S69P009N049N053P050(0)='1' AND  B( 6)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar2S7S69N027P029P011nsss(0) <='1';
          else
          cVar2S7S69N027P029P011nsss(0) <='0';
          end if;
        if(cVar1S8S69P009N049N053P050(0)='1' AND  B( 6)='0' AND B( 5)='0' AND A( 2)='1' )then
          cVar2S8S69N027N029P015nsss(0) <='1';
          else
          cVar2S8S69N027N029P015nsss(0) <='0';
          end if;
        if(cVar1S9S69P009N049N053N050(0)='1' AND  E(13)='0' AND A( 0)='1' AND A(18)='0' )then
          cVar2S9S69P051P019P002nsss(0) <='1';
          else
          cVar2S9S69P051P019P002nsss(0) <='0';
          end if;
        if(cVar1S10S69P009N049N053N050(0)='1' AND  E(13)='0' AND A( 0)='0' AND E( 1)='0' )then
          cVar2S10S69P051N019P066nsss(0) <='1';
          else
          cVar2S10S69P051N019P066nsss(0) <='0';
          end if;
        if(cVar1S12S69N009P041P020N003(0)='1' AND  A(18)='1' )then
          cVar2S12S69P002nsss(0) <='1';
          else
          cVar2S12S69P002nsss(0) <='0';
          end if;
        if(cVar1S13S69N009P041P020N003(0)='1' AND  A(18)='0' AND A(17)='1' )then
          cVar2S13S69N002P004nsss(0) <='1';
          else
          cVar2S13S69N002P004nsss(0) <='0';
          end if;
        if(cVar1S14S69N009P041P020N003(0)='1' AND  A(18)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S14S69N002N004P005nsss(0) <='1';
          else
          cVar2S14S69N002N004P005nsss(0) <='0';
          end if;
        if(cVar1S16S69N009P041N020N001(0)='1' AND  B( 9)='1' AND D( 7)='0' )then
          cVar2S16S69P021P040nsss(0) <='1';
          else
          cVar2S16S69P021P040nsss(0) <='0';
          end if;
        if(cVar1S17S69N009P041N020N001(0)='1' AND  B( 9)='1' AND D( 7)='1' AND E( 7)='0' )then
          cVar2S17S69P021P040P042nsss(0) <='1';
          else
          cVar2S17S69P021P040P042nsss(0) <='0';
          end if;
        if(cVar1S18S69N009P041N020N001(0)='1' AND  B( 9)='0' AND B( 0)='0' AND E(15)='1' )then
          cVar2S18S69N021P039P043nsss(0) <='1';
          else
          cVar2S18S69N021P039P043nsss(0) <='0';
          end if;
        if(cVar1S19S69N009N041P031P013(0)='1' AND  E( 4)='1' AND A(13)='0' AND D( 9)='0' )then
          cVar2S19S69P054P012P065nsss(0) <='1';
          else
          cVar2S19S69P054P012P065nsss(0) <='0';
          end if;
        if(cVar1S20S69N009N041P031P013(0)='1' AND  E( 4)='1' AND A(13)='1' )then
          cVar2S20S69P054P012psss(0) <='1';
          else
          cVar2S20S69P054P012psss(0) <='0';
          end if;
        if(cVar1S21S69N009N041P031P013(0)='1' AND  E( 4)='0' AND D(11)='1' )then
          cVar2S21S69N054P057nsss(0) <='1';
          else
          cVar2S21S69N054P057nsss(0) <='0';
          end if;
        if(cVar1S22S69N009N041P031P013(0)='1' AND  E( 4)='0' AND D(11)='0' AND E( 3)='1' )then
          cVar2S22S69N054N057P058nsss(0) <='1';
          else
          cVar2S22S69N054N057P058nsss(0) <='0';
          end if;
        if(cVar1S23S69N009N041P031N013(0)='1' AND  E( 4)='1' AND A(11)='0' )then
          cVar2S23S69P054P016nsss(0) <='1';
          else
          cVar2S23S69P054P016nsss(0) <='0';
          end if;
        if(cVar1S24S69N009N041P031N013(0)='1' AND  E( 4)='0' AND A(10)='1' AND A(13)='1' )then
          cVar2S24S69N054P018P012nsss(0) <='1';
          else
          cVar2S24S69N054P018P012nsss(0) <='0';
          end if;
        if(cVar1S25S69N009N041N031P054(0)='1' AND  B( 0)='0' AND A(11)='1' AND E(11)='0' )then
          cVar2S25S69P039P016P059nsss(0) <='1';
          else
          cVar2S25S69P039P016P059nsss(0) <='0';
          end if;
        if(cVar1S26S69N009N041N031P054(0)='1' AND  B( 0)='0' AND A(11)='0' AND B( 7)='1' )then
          cVar2S26S69P039N016P025nsss(0) <='1';
          else
          cVar2S26S69P039N016P025nsss(0) <='0';
          end if;
        if(cVar1S27S69N009N041N031P054(0)='1' AND  B( 0)='1' AND A( 4)='0' AND D( 1)='1' )then
          cVar2S27S69P039P011P064nsss(0) <='1';
          else
          cVar2S27S69P039P011P064nsss(0) <='0';
          end if;
        if(cVar1S28S69N009N041N031P054(0)='1' AND  A( 4)='1' AND B( 5)='1' )then
          cVar2S28S69P011P029nsss(0) <='1';
          else
          cVar2S28S69P011P029nsss(0) <='0';
          end if;
        if(cVar1S29S69N009N041N031P054(0)='1' AND  A( 4)='1' AND B( 5)='0' AND A(13)='1' )then
          cVar2S29S69P011N029P012nsss(0) <='1';
          else
          cVar2S29S69P011N029P012nsss(0) <='0';
          end if;
        if(cVar1S30S69N009N041N031P054(0)='1' AND  A( 4)='0' AND A(14)='1' )then
          cVar2S30S69N011P010nsss(0) <='1';
          else
          cVar2S30S69N011P010nsss(0) <='0';
          end if;
        if(cVar1S31S69N009N041N031P054(0)='1' AND  A( 4)='0' AND A(14)='0' AND B(14)='1' )then
          cVar2S31S69N011N010P030nsss(0) <='1';
          else
          cVar2S31S69N011N010P030nsss(0) <='0';
          end if;
        if(cVar1S0S70P016P018P036P053(0)='1' AND  A(12)='0' AND B(15)='1' AND A( 2)='0' )then
          cVar2S0S70P014P028P015nsss(0) <='1';
          else
          cVar2S0S70P014P028P015nsss(0) <='0';
          end if;
        if(cVar1S1S70P016P018P036P053(0)='1' AND  A(12)='0' AND B(15)='0' )then
          cVar2S1S70P014N028psss(0) <='1';
          else
          cVar2S1S70P014N028psss(0) <='0';
          end if;
        if(cVar1S2S70P016P018P036P053(0)='1' AND  A(12)='1' AND A( 5)='1' )then
          cVar2S2S70P014P009nsss(0) <='1';
          else
          cVar2S2S70P014P009nsss(0) <='0';
          end if;
        if(cVar1S3S70P016P018P036N053(0)='1' AND  B( 8)='1' AND A( 7)='1' )then
          cVar2S3S70P023P005nsss(0) <='1';
          else
          cVar2S3S70P023P005nsss(0) <='0';
          end if;
        if(cVar1S4S70P016P018P036N053(0)='1' AND  B( 8)='1' AND A( 7)='0' AND A( 1)='0' )then
          cVar2S4S70P023N005P017nsss(0) <='1';
          else
          cVar2S4S70P023N005P017nsss(0) <='0';
          end if;
        if(cVar1S5S70P016P018P036N053(0)='1' AND  B( 8)='0' AND D(13)='1' AND B(16)='1' )then
          cVar2S5S70N023P049P026nsss(0) <='1';
          else
          cVar2S5S70N023P049P026nsss(0) <='0';
          end if;
        if(cVar1S6S70P016P018P036N053(0)='1' AND  B( 8)='0' AND D(13)='0' AND E(14)='0' )then
          cVar2S6S70N023N049P047nsss(0) <='1';
          else
          cVar2S6S70N023N049P047nsss(0) <='0';
          end if;
        if(cVar1S7S70P016P018P036P017(0)='1' AND  B( 1)='0' AND D( 3)='0' )then
          cVar2S7S70P037P056nsss(0) <='1';
          else
          cVar2S7S70P037P056nsss(0) <='0';
          end if;
        if(cVar1S8S70P016P018P036P017(0)='1' AND  B( 1)='1' AND A( 0)='0' )then
          cVar2S8S70P037P019nsss(0) <='1';
          else
          cVar2S8S70P037P019nsss(0) <='0';
          end if;
        if(cVar1S9S70P016P018P036N017(0)='1' AND  A( 0)='1' AND D( 9)='1' )then
          cVar2S9S70P019P065nsss(0) <='1';
          else
          cVar2S9S70P019P065nsss(0) <='0';
          end if;
        if(cVar1S10S70P016P018P036N017(0)='1' AND  A( 0)='1' AND D( 9)='0' AND A( 2)='0' )then
          cVar2S10S70P019N065P015nsss(0) <='1';
          else
          cVar2S10S70P019N065P015nsss(0) <='0';
          end if;
        if(cVar1S11S70P016P018P036N017(0)='1' AND  A( 0)='0' AND D( 9)='0' AND A( 4)='1' )then
          cVar2S11S70N019P065P011nsss(0) <='1';
          else
          cVar2S11S70N019P065P011nsss(0) <='0';
          end if;
        if(cVar1S12S70P016P018P045P017(0)='1' AND  A( 3)='0' )then
          cVar2S12S70P013nsss(0) <='1';
          else
          cVar2S12S70P013nsss(0) <='0';
          end if;
        if(cVar1S13S70P016P018N045P026(0)='1' AND  E(14)='0' AND A( 5)='0' )then
          cVar2S13S70P047P009nsss(0) <='1';
          else
          cVar2S13S70P047P009nsss(0) <='0';
          end if;
        if(cVar1S14S70P016P018N045P026(0)='1' AND  E(14)='1' AND A( 5)='1' )then
          cVar2S14S70P047P009nsss(0) <='1';
          else
          cVar2S14S70P047P009nsss(0) <='0';
          end if;
        if(cVar1S15S70P016P018N045P026(0)='1' AND  E(14)='1' AND A( 5)='0' AND A( 1)='1' )then
          cVar2S15S70P047N009P017nsss(0) <='1';
          else
          cVar2S15S70P047N009P017nsss(0) <='0';
          end if;
        if(cVar1S16S70P016P018N045P026(0)='1' AND  D(13)='1' )then
          cVar2S16S70P049nsss(0) <='1';
          else
          cVar2S16S70P049nsss(0) <='0';
          end if;
        if(cVar1S17S70P016P018N045P026(0)='1' AND  D(13)='0' AND D( 4)='1' )then
          cVar2S17S70N049P052nsss(0) <='1';
          else
          cVar2S17S70N049P052nsss(0) <='0';
          end if;
        if(cVar1S18S70P016P035P053P041(0)='1' AND  D( 7)='1' )then
          cVar2S18S70P040nsss(0) <='1';
          else
          cVar2S18S70P040nsss(0) <='0';
          end if;
        if(cVar1S19S70P016P035P053P041(0)='1' AND  D( 7)='0' AND A(13)='0' )then
          cVar2S19S70N040P012nsss(0) <='1';
          else
          cVar2S19S70N040P012nsss(0) <='0';
          end if;
        if(cVar1S20S70P016P035P053N041(0)='1' AND  E( 7)='0' AND E(14)='1' AND D( 0)='1' )then
          cVar2S20S70P042P047P068nsss(0) <='1';
          else
          cVar2S20S70P042P047P068nsss(0) <='0';
          end if;
        if(cVar1S21S70P016P035P053N041(0)='1' AND  E( 7)='1' AND A( 7)='1' )then
          cVar2S21S70P042P005nsss(0) <='1';
          else
          cVar2S21S70P042P005nsss(0) <='0';
          end if;
        if(cVar1S22S70P016P035P053N041(0)='1' AND  E( 7)='1' AND A( 7)='0' AND A(13)='1' )then
          cVar2S22S70P042N005P012nsss(0) <='1';
          else
          cVar2S22S70P042N005P012nsss(0) <='0';
          end if;
        if(cVar1S23S70P016P035P053P037(0)='1' AND  A( 0)='1' )then
          cVar2S23S70P019nsss(0) <='1';
          else
          cVar2S23S70P019nsss(0) <='0';
          end if;
        if(cVar1S24S70P016P035P053N037(0)='1' AND  B(11)='0' AND A( 2)='1' AND A( 0)='1' )then
          cVar2S24S70P036P015P019nsss(0) <='1';
          else
          cVar2S24S70P036P015P019nsss(0) <='0';
          end if;
        if(cVar1S25S70P016P035P053N037(0)='1' AND  B(11)='0' AND A( 2)='0' AND A( 5)='1' )then
          cVar2S25S70P036N015P009nsss(0) <='1';
          else
          cVar2S25S70P036N015P009nsss(0) <='0';
          end if;
        if(cVar1S27S70P016P035N032P034(0)='1' AND  A(14)='0' AND A( 5)='1' AND A( 2)='0' )then
          cVar2S27S70P010P009P015nsss(0) <='1';
          else
          cVar2S27S70P010P009P015nsss(0) <='0';
          end if;
        if(cVar1S2S71P041P020N003N002(0)='1' AND  A(17)='1' )then
          cVar2S2S71P004nsss(0) <='1';
          else
          cVar2S2S71P004nsss(0) <='0';
          end if;
        if(cVar1S3S71P041P020N003N002(0)='1' AND  A(17)='0' AND A( 7)='1' )then
          cVar2S3S71N004P005nsss(0) <='1';
          else
          cVar2S3S71N004P005nsss(0) <='0';
          end if;
        if(cVar1S5S71P041N020N001P005(0)='1' AND  B( 9)='1' AND D( 7)='0' )then
          cVar2S5S71P021P040nsss(0) <='1';
          else
          cVar2S5S71P021P040nsss(0) <='0';
          end if;
        if(cVar1S6S71P041N020N001P005(0)='1' AND  B( 9)='0' AND B(18)='1' )then
          cVar2S6S71N021P022nsss(0) <='1';
          else
          cVar2S6S71N021P022nsss(0) <='0';
          end if;
        if(cVar1S7S71P041N020N001P005(0)='1' AND  B( 9)='0' AND B(18)='0' AND E( 7)='1' )then
          cVar2S7S71N021N022P042nsss(0) <='1';
          else
          cVar2S7S71N021N022P042nsss(0) <='0';
          end if;
        if(cVar1S8S71P041N020N001N005(0)='1' AND  B( 0)='0' AND E( 9)='1' )then
          cVar2S8S71P039P067nsss(0) <='1';
          else
          cVar2S8S71P039P067nsss(0) <='0';
          end if;
        if(cVar1S9S71P041N020N001N005(0)='1' AND  B( 0)='0' AND E( 9)='0' AND B(18)='1' )then
          cVar2S9S71P039N067P022nsss(0) <='1';
          else
          cVar2S9S71P039N067P022nsss(0) <='0';
          end if;
        if(cVar1S10S71P041N020N001N005(0)='1' AND  B( 0)='1' AND A( 1)='0' AND B( 9)='1' )then
          cVar2S10S71P039P017P021nsss(0) <='1';
          else
          cVar2S10S71P039P017P021nsss(0) <='0';
          end if;
        if(cVar1S11S71N041P049P026P033(0)='1' AND  B(17)='0' )then
          cVar2S11S71P024nsss(0) <='1';
          else
          cVar2S11S71P024nsss(0) <='0';
          end if;
        if(cVar1S12S71N041P049N026P024(0)='1' AND  A(16)='1' )then
          cVar2S12S71P006nsss(0) <='1';
          else
          cVar2S12S71P006nsss(0) <='0';
          end if;
        if(cVar1S13S71N041P049N026P024(0)='1' AND  A(16)='0' AND A(11)='0' )then
          cVar2S13S71N006P016nsss(0) <='1';
          else
          cVar2S13S71N006P016nsss(0) <='0';
          end if;
        if(cVar1S14S71N041P049N026N024(0)='1' AND  B( 6)='1' AND D( 5)='0' )then
          cVar2S14S71P027P048nsss(0) <='1';
          else
          cVar2S14S71P027P048nsss(0) <='0';
          end if;
        if(cVar1S15S71N041P049N026N024(0)='1' AND  B( 6)='1' AND D( 5)='1' AND E(14)='0' )then
          cVar2S15S71P027P048P047nsss(0) <='1';
          else
          cVar2S15S71P027P048P047nsss(0) <='0';
          end if;
        if(cVar1S16S71N041P049N026N024(0)='1' AND  B( 6)='0' AND B( 7)='1' )then
          cVar2S16S71N027P025nsss(0) <='1';
          else
          cVar2S16S71N027P025nsss(0) <='0';
          end if;
        if(cVar1S17S71N041N049P039P045(0)='1' AND  A( 6)='1' AND B( 1)='0' )then
          cVar2S17S71P007P037nsss(0) <='1';
          else
          cVar2S17S71P007P037nsss(0) <='0';
          end if;
        if(cVar1S18S71N041N049P039P045(0)='1' AND  A( 6)='0' AND A(17)='1' AND A( 3)='0' )then
          cVar2S18S71N007P004P013nsss(0) <='1';
          else
          cVar2S18S71N007P004P013nsss(0) <='0';
          end if;
        if(cVar1S19S71N041N049P039P045(0)='1' AND  A( 6)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S19S71N007N004P005nsss(0) <='1';
          else
          cVar2S19S71N007N004P005nsss(0) <='0';
          end if;
        if(cVar1S20S71N041N049P039N045(0)='1' AND  E(14)='0' AND A(11)='1' AND B( 2)='0' )then
          cVar2S20S71P047P016P035nsss(0) <='1';
          else
          cVar2S20S71P047P016P035nsss(0) <='0';
          end if;
        if(cVar1S21S71N041N049P039N045(0)='1' AND  E(14)='0' AND A(11)='0' AND D(12)='1' )then
          cVar2S21S71P047N016P053nsss(0) <='1';
          else
          cVar2S21S71P047N016P053nsss(0) <='0';
          end if;
        if(cVar1S22S71N041N049P039N045(0)='1' AND  E(14)='1' AND D( 8)='1' )then
          cVar2S22S71P047P069nsss(0) <='1';
          else
          cVar2S22S71P047P069nsss(0) <='0';
          end if;
        if(cVar1S23S71N041N049P039N045(0)='1' AND  E(14)='1' AND D( 8)='0' AND A(15)='1' )then
          cVar2S23S71P047N069P008nsss(0) <='1';
          else
          cVar2S23S71P047N069P008nsss(0) <='0';
          end if;
        if(cVar1S25S71N041N049P039N036(0)='1' AND  A( 4)='0' AND B(19)='1' )then
          cVar2S25S71P011P020nsss(0) <='1';
          else
          cVar2S25S71P011P020nsss(0) <='0';
          end if;
        if(cVar1S26S71N041N049P039N036(0)='1' AND  A( 4)='0' AND B(19)='0' AND A( 3)='1' )then
          cVar2S26S71P011N020P013nsss(0) <='1';
          else
          cVar2S26S71P011N020P013nsss(0) <='0';
          end if;
        if(cVar1S1S72P016P018P023N042(0)='1' AND  E(15)='1' )then
          cVar2S1S72P043nsss(0) <='1';
          else
          cVar2S1S72P043nsss(0) <='0';
          end if;
        if(cVar1S2S72P016P018P023N042(0)='1' AND  E(15)='0' AND A( 1)='0' AND A( 0)='1' )then
          cVar2S2S72N043P017P019nsss(0) <='1';
          else
          cVar2S2S72N043P017P019nsss(0) <='0';
          end if;
        if(cVar1S3S72P016P018N023P047(0)='1' AND  A(16)='1' )then
          cVar2S3S72P006nsss(0) <='1';
          else
          cVar2S3S72P006nsss(0) <='0';
          end if;
        if(cVar1S4S72P016P018N023P047(0)='1' AND  A(16)='0' AND A(15)='1' )then
          cVar2S4S72N006P008nsss(0) <='1';
          else
          cVar2S4S72N006P008nsss(0) <='0';
          end if;
        if(cVar1S5S72P016P018N023P047(0)='1' AND  A(16)='0' AND A(15)='0' AND A( 6)='1' )then
          cVar2S5S72N006N008P007nsss(0) <='1';
          else
          cVar2S5S72N006N008P007nsss(0) <='0';
          end if;
        if(cVar1S6S72P016P018N023N047(0)='1' AND  B(15)='1' AND B(13)='0' )then
          cVar2S6S72P028P032nsss(0) <='1';
          else
          cVar2S6S72P028P032nsss(0) <='0';
          end if;
        if(cVar1S7S72P016P018N023N047(0)='1' AND  B(15)='0' AND B( 4)='1' AND E( 4)='1' )then
          cVar2S7S72N028P031P054nsss(0) <='1';
          else
          cVar2S7S72N028P031P054nsss(0) <='0';
          end if;
        if(cVar1S8S72P016P018N023N047(0)='1' AND  B(15)='0' AND B( 4)='0' AND E( 4)='0' )then
          cVar2S8S72N028N031P054nsss(0) <='1';
          else
          cVar2S8S72N028N031P054nsss(0) <='0';
          end if;
        if(cVar1S10S72P016P018P045N015(0)='1' AND  A( 1)='0' )then
          cVar2S10S72P017nsss(0) <='1';
          else
          cVar2S10S72P017nsss(0) <='0';
          end if;
        if(cVar1S11S72P016P018N045P013(0)='1' AND  E(14)='0' AND B(15)='1' )then
          cVar2S11S72P047P028nsss(0) <='1';
          else
          cVar2S11S72P047P028nsss(0) <='0';
          end if;
        if(cVar1S12S72P016P018N045P013(0)='1' AND  E(14)='0' AND B(15)='0' AND E( 4)='0' )then
          cVar2S12S72P047N028P054nsss(0) <='1';
          else
          cVar2S12S72P047N028P054nsss(0) <='0';
          end if;
        if(cVar1S13S72P016P018N045P013(0)='1' AND  E(14)='1' AND A( 5)='1' )then
          cVar2S13S72P047P009nsss(0) <='1';
          else
          cVar2S13S72P047P009nsss(0) <='0';
          end if;
        if(cVar1S14S72P016P018N045P013(0)='1' AND  E(14)='1' AND A( 5)='0' AND A( 1)='1' )then
          cVar2S14S72P047N009P017nsss(0) <='1';
          else
          cVar2S14S72P047N009P017nsss(0) <='0';
          end if;
        if(cVar1S15S72P016P018N045P013(0)='1' AND  B( 4)='1' )then
          cVar2S15S72P031nsss(0) <='1';
          else
          cVar2S15S72P031nsss(0) <='0';
          end if;
        if(cVar1S16S72P016P018N045P013(0)='1' AND  B( 4)='0' AND E( 6)='1' )then
          cVar2S16S72N031P046nsss(0) <='1';
          else
          cVar2S16S72N031P046nsss(0) <='0';
          end if;
        if(cVar1S17S72P016P018N045P013(0)='1' AND  B( 4)='0' AND E( 6)='0' AND B( 5)='1' )then
          cVar2S17S72N031N046P029nsss(0) <='1';
          else
          cVar2S17S72N031N046P029nsss(0) <='0';
          end if;
        if(cVar1S18S72P016P033P041P011(0)='1' AND  A( 0)='0' AND B(19)='0' )then
          cVar2S18S72P019P020nsss(0) <='1';
          else
          cVar2S18S72P019P020nsss(0) <='0';
          end if;
        if(cVar1S19S72P016P033P041P011(0)='1' AND  A( 0)='1' AND B( 0)='0' )then
          cVar2S19S72P019P039nsss(0) <='1';
          else
          cVar2S19S72P019P039nsss(0) <='0';
          end if;
        if(cVar1S20S72P016P033N041P009(0)='1' AND  B( 5)='1' )then
          cVar2S20S72P029nsss(0) <='1';
          else
          cVar2S20S72P029nsss(0) <='0';
          end if;
        if(cVar1S21S72P016P033N041P009(0)='1' AND  B( 5)='0' AND A( 6)='0' )then
          cVar2S21S72N029P007nsss(0) <='1';
          else
          cVar2S21S72N029P007nsss(0) <='0';
          end if;
        if(cVar1S22S72P016P033N041P009(0)='1' AND  B( 5)='0' AND A( 6)='1' AND A(12)='1' )then
          cVar2S22S72N029P007P014nsss(0) <='1';
          else
          cVar2S22S72N029P007P014nsss(0) <='0';
          end if;
        if(cVar1S23S72P016P033N041N009(0)='1' AND  D(12)='0' AND A(17)='1' )then
          cVar2S23S72P053P004nsss(0) <='1';
          else
          cVar2S23S72P053P004nsss(0) <='0';
          end if;
        if(cVar1S24S72P016P033N041N009(0)='1' AND  D(12)='1' AND A( 4)='1' AND A( 0)='1' )then
          cVar2S24S72P053P011P019nsss(0) <='1';
          else
          cVar2S24S72P053P011P019nsss(0) <='0';
          end if;
        if(cVar1S25S72P016P033P069P068(0)='1' AND  A( 3)='1' )then
          cVar2S25S72P013nsss(0) <='1';
          else
          cVar2S25S72P013nsss(0) <='0';
          end if;
        if(cVar1S26S72P016P033P069P068(0)='1' AND  A( 3)='0' AND A( 2)='1' )then
          cVar2S26S72N013P015nsss(0) <='1';
          else
          cVar2S26S72N013P015nsss(0) <='0';
          end if;
        if(cVar1S27S72P016P033P069N068(0)='1' AND  A( 6)='1' )then
          cVar2S27S72P007nsss(0) <='1';
          else
          cVar2S27S72P007nsss(0) <='0';
          end if;
        if(cVar1S28S72P016P033P069N068(0)='1' AND  A( 6)='0' AND A(10)='1' AND A( 8)='0' )then
          cVar2S28S72N007P018P003nsss(0) <='1';
          else
          cVar2S28S72N007P018P003nsss(0) <='0';
          end if;
        if(cVar1S29S72P016P033P069N068(0)='1' AND  A( 6)='0' AND A(10)='0' AND B( 1)='1' )then
          cVar2S29S72N007N018P037nsss(0) <='1';
          else
          cVar2S29S72N007N018P037nsss(0) <='0';
          end if;
        if(cVar1S30S72P016P033P069P067(0)='1' AND  B(11)='1' )then
          cVar2S30S72P036nsss(0) <='1';
          else
          cVar2S30S72P036nsss(0) <='0';
          end if;
        if(cVar1S3S73P047N006P008N026(0)='1' AND  D(13)='1' )then
          cVar2S3S73P049nsss(0) <='1';
          else
          cVar2S3S73P049nsss(0) <='0';
          end if;
        if(cVar1S4S73P047N006N008P007(0)='1' AND  A( 2)='0' AND D( 0)='0' )then
          cVar2S4S73P015P068nsss(0) <='1';
          else
          cVar2S4S73P015P068nsss(0) <='0';
          end if;
        if(cVar1S5S73P047N006N008N007(0)='1' AND  A( 5)='1' AND A( 1)='0' )then
          cVar2S5S73P009P017nsss(0) <='1';
          else
          cVar2S5S73P009P017nsss(0) <='0';
          end if;
        if(cVar1S6S73P047N006N008N007(0)='1' AND  A( 5)='0' AND A( 7)='1' )then
          cVar2S6S73N009P005nsss(0) <='1';
          else
          cVar2S6S73N009P005nsss(0) <='0';
          end if;
        if(cVar1S7S73P047N006N008N007(0)='1' AND  A( 5)='0' AND A( 7)='0' AND D( 8)='1' )then
          cVar2S7S73N009N005P069nsss(0) <='1';
          else
          cVar2S7S73N009N005P069nsss(0) <='0';
          end if;
        if(cVar1S8S73N047P031P013P056(0)='1' AND  A(13)='0' )then
          cVar2S8S73P012nsss(0) <='1';
          else
          cVar2S8S73P012nsss(0) <='0';
          end if;
        if(cVar1S9S73N047P031P013P056(0)='1' AND  A(13)='1' AND A( 1)='0' )then
          cVar2S9S73P012P017nsss(0) <='1';
          else
          cVar2S9S73P012P017nsss(0) <='0';
          end if;
        if(cVar1S10S73N047P031P013N056(0)='1' AND  D(11)='1' )then
          cVar2S10S73P057nsss(0) <='1';
          else
          cVar2S10S73P057nsss(0) <='0';
          end if;
        if(cVar1S11S73N047P031P013N056(0)='1' AND  D(11)='0' AND D( 2)='1' AND A( 2)='0' )then
          cVar2S11S73N057P060P015nsss(0) <='1';
          else
          cVar2S11S73N057P060P015nsss(0) <='0';
          end if;
        if(cVar1S12S73N047P031P013N056(0)='1' AND  D(11)='0' AND D( 2)='0' AND A(11)='1' )then
          cVar2S12S73N057N060P016nsss(0) <='1';
          else
          cVar2S12S73N057N060P016nsss(0) <='0';
          end if;
        if(cVar1S13S73N047P031N013P011(0)='1' AND  A(15)='0' AND E(12)='1' )then
          cVar2S13S73P008P055nsss(0) <='1';
          else
          cVar2S13S73P008P055nsss(0) <='0';
          end if;
        if(cVar1S14S73N047P031N013P011(0)='1' AND  A(15)='0' AND E(12)='0' AND A(11)='0' )then
          cVar2S14S73P008N055P016nsss(0) <='1';
          else
          cVar2S14S73P008N055P016nsss(0) <='0';
          end if;
        if(cVar1S15S73N047P031N013N011(0)='1' AND  E(12)='0' AND A(13)='1' )then
          cVar2S15S73P055P012nsss(0) <='1';
          else
          cVar2S15S73P055P012nsss(0) <='0';
          end if;
        if(cVar1S16S73N047P031N013N011(0)='1' AND  E(12)='0' AND A(13)='0' AND A(10)='1' )then
          cVar2S16S73P055N012P018nsss(0) <='1';
          else
          cVar2S16S73P055N012P018nsss(0) <='0';
          end if;
        if(cVar1S17S73N047N031P030P012(0)='1' AND  D( 3)='1' )then
          cVar2S17S73P056nsss(0) <='1';
          else
          cVar2S17S73P056nsss(0) <='0';
          end if;
        if(cVar1S18S73N047N031P030P012(0)='1' AND  D( 3)='0' AND D(11)='1' AND D( 9)='0' )then
          cVar2S18S73N056P057P065nsss(0) <='1';
          else
          cVar2S18S73N056P057P065nsss(0) <='0';
          end if;
        if(cVar1S19S73N047N031P030P012(0)='1' AND  D( 3)='0' AND D(11)='0' AND E(11)='1' )then
          cVar2S19S73N056N057P059nsss(0) <='1';
          else
          cVar2S19S73N056N057P059nsss(0) <='0';
          end if;
        if(cVar1S20S73N047N031P030N012(0)='1' AND  A(14)='1' AND D(11)='1' )then
          cVar2S20S73P010P057nsss(0) <='1';
          else
          cVar2S20S73P010P057nsss(0) <='0';
          end if;
        if(cVar1S21S73N047N031P030N012(0)='1' AND  A(14)='1' AND D(11)='0' AND A( 1)='1' )then
          cVar2S21S73P010N057P017nsss(0) <='1';
          else
          cVar2S21S73P010N057P017nsss(0) <='0';
          end if;
        if(cVar1S22S73N047N031P030N012(0)='1' AND  A(14)='0' AND A( 3)='1' AND D(11)='1' )then
          cVar2S22S73N010P013P057nsss(0) <='1';
          else
          cVar2S22S73N010P013P057nsss(0) <='0';
          end if;
        if(cVar1S23S73N047N031N030P057(0)='1' AND  A( 0)='1' AND E( 1)='1' AND D( 9)='0' )then
          cVar2S23S73P019P066P065nsss(0) <='1';
          else
          cVar2S23S73P019P066P065nsss(0) <='0';
          end if;
        if(cVar1S24S73N047N031N030P057(0)='1' AND  A( 0)='1' AND E( 1)='0' AND A( 3)='1' )then
          cVar2S24S73P019N066P013nsss(0) <='1';
          else
          cVar2S24S73P019N066P013nsss(0) <='0';
          end if;
        if(cVar1S25S73N047N031N030P057(0)='1' AND  A( 0)='0' AND D( 0)='0' AND D( 1)='1' )then
          cVar2S25S73N019P068P064nsss(0) <='1';
          else
          cVar2S25S73N019P068P064nsss(0) <='0';
          end if;
        if(cVar1S26S73N047N031N030P057(0)='1' AND  B(13)='1' )then
          cVar2S26S73P032nsss(0) <='1';
          else
          cVar2S26S73P032nsss(0) <='0';
          end if;
        if(cVar1S27S73N047N031N030P057(0)='1' AND  B(13)='0' AND B(15)='1' AND A(14)='1' )then
          cVar2S27S73N032P028P010nsss(0) <='1';
          else
          cVar2S27S73N032P028P010nsss(0) <='0';
          end if;
        if(cVar1S28S73N047N031N030P057(0)='1' AND  B(13)='0' AND B(15)='0' AND D( 0)='1' )then
          cVar2S28S73N032N028P068nsss(0) <='1';
          else
          cVar2S28S73N032N028P068nsss(0) <='0';
          end if;
        if(cVar1S0S74P064P066P027P009(0)='1' AND  A( 1)='0' AND A( 2)='0' )then
          cVar2S0S74P017P015nsss(0) <='1';
          else
          cVar2S0S74P017P015nsss(0) <='0';
          end if;
        if(cVar1S1S74P064P066P027P009(0)='1' AND  A( 1)='0' AND A( 2)='1' AND D( 5)='1' )then
          cVar2S1S74P017P015P048nsss(0) <='1';
          else
          cVar2S1S74P017P015P048nsss(0) <='0';
          end if;
        if(cVar1S2S74P064P066P027P009(0)='1' AND  A( 1)='1' AND D( 4)='1' )then
          cVar2S2S74P017P052nsss(0) <='1';
          else
          cVar2S2S74P017P052nsss(0) <='0';
          end if;
        if(cVar1S3S74P064P066P027P009(0)='1' AND  A( 1)='1' AND D( 4)='0' AND A( 0)='1' )then
          cVar2S3S74P017N052P019nsss(0) <='1';
          else
          cVar2S3S74P017N052P019nsss(0) <='0';
          end if;
        if(cVar1S4S74P064P066P027N009(0)='1' AND  A( 6)='1' )then
          cVar2S4S74P007nsss(0) <='1';
          else
          cVar2S4S74P007nsss(0) <='0';
          end if;
        if(cVar1S5S74P064P066P027N009(0)='1' AND  A( 6)='0' AND A(15)='1' )then
          cVar2S5S74N007P008nsss(0) <='1';
          else
          cVar2S5S74N007P008nsss(0) <='0';
          end if;
        if(cVar1S6S74P064P066P027N009(0)='1' AND  A( 6)='0' AND A(15)='0' AND A( 4)='1' )then
          cVar2S6S74N007N008P011nsss(0) <='1';
          else
          cVar2S6S74N007N008P011nsss(0) <='0';
          end if;
        if(cVar1S7S74P064P066N027P041(0)='1' AND  B(19)='1' AND A( 8)='1' )then
          cVar2S7S74P020P003nsss(0) <='1';
          else
          cVar2S7S74P020P003nsss(0) <='0';
          end if;
        if(cVar1S8S74P064P066N027P041(0)='1' AND  B(19)='1' AND A( 8)='0' AND A(18)='1' )then
          cVar2S8S74P020N003P002nsss(0) <='1';
          else
          cVar2S8S74P020N003P002nsss(0) <='0';
          end if;
        if(cVar1S9S74P064P066N027P041(0)='1' AND  B(19)='0' AND A( 7)='1' )then
          cVar2S9S74N020P005nsss(0) <='1';
          else
          cVar2S9S74N020P005nsss(0) <='0';
          end if;
        if(cVar1S10S74P064P066N027P041(0)='1' AND  B(19)='0' AND A( 7)='0' AND A(13)='0' )then
          cVar2S10S74N020N005P012nsss(0) <='1';
          else
          cVar2S10S74N020N005P012nsss(0) <='0';
          end if;
        if(cVar1S11S74P064P066N027N041(0)='1' AND  B( 5)='1' AND A( 4)='1' AND A(15)='0' )then
          cVar2S11S74P029P011P008nsss(0) <='1';
          else
          cVar2S11S74P029P011P008nsss(0) <='0';
          end if;
        if(cVar1S12S74P064P066N027N041(0)='1' AND  B( 5)='1' AND A( 4)='0' AND A( 5)='1' )then
          cVar2S12S74P029N011P009nsss(0) <='1';
          else
          cVar2S12S74P029N011P009nsss(0) <='0';
          end if;
        if(cVar1S13S74P064P066N027N041(0)='1' AND  B( 5)='0' AND B(15)='1' )then
          cVar2S13S74N029P028nsss(0) <='1';
          else
          cVar2S13S74N029P028nsss(0) <='0';
          end if;
        if(cVar1S14S74P064P066N027N041(0)='1' AND  B( 5)='0' AND B(15)='0' AND D(12)='0' )then
          cVar2S14S74N029N028P053nsss(0) <='1';
          else
          cVar2S14S74N029N028P053nsss(0) <='0';
          end if;
        if(cVar1S15S74P064P066P006P059(0)='1' AND  B( 8)='0' AND E( 7)='0' AND A(13)='0' )then
          cVar2S15S74P023P042P012nsss(0) <='1';
          else
          cVar2S15S74P023P042P012nsss(0) <='0';
          end if;
        if(cVar1S16S74P064P066P006P059(0)='1' AND  B( 8)='1' AND E( 7)='1' )then
          cVar2S16S74P023P042nsss(0) <='1';
          else
          cVar2S16S74P023P042nsss(0) <='0';
          end if;
        if(cVar1S17S74P064P066P006P059(0)='1' AND  D( 0)='1' AND A( 3)='1' )then
          cVar2S17S74P068P013nsss(0) <='1';
          else
          cVar2S17S74P068P013nsss(0) <='0';
          end if;
        if(cVar1S18S74P064P066P006P035(0)='1' AND  A(13)='1' AND A(10)='0' )then
          cVar2S18S74P012P018nsss(0) <='1';
          else
          cVar2S18S74P012P018nsss(0) <='0';
          end if;
        if(cVar1S19S74P064P066P006P035(0)='1' AND  A(13)='0' AND A( 4)='1' )then
          cVar2S19S74N012P011nsss(0) <='1';
          else
          cVar2S19S74N012P011nsss(0) <='0';
          end if;
        if(cVar1S21S74P064P011N042P003(0)='1' AND  B( 5)='0' AND A( 5)='0' AND E( 9)='0' )then
          cVar2S21S74P029P009P067nsss(0) <='1';
          else
          cVar2S21S74P029P009P067nsss(0) <='0';
          end if;
        if(cVar1S22S74P064P011N042P003(0)='1' AND  B( 5)='0' AND A( 5)='1' AND B( 6)='1' )then
          cVar2S22S74P029P009P027nsss(0) <='1';
          else
          cVar2S22S74P029P009P027nsss(0) <='0';
          end if;
        if(cVar1S23S74P064P011N042P003(0)='1' AND  A(14)='1' )then
          cVar2S23S74P010nsss(0) <='1';
          else
          cVar2S23S74P010nsss(0) <='0';
          end if;
        if(cVar1S24S74P064P011N042P003(0)='1' AND  A(14)='0' AND A( 5)='1' )then
          cVar2S24S74N010P009nsss(0) <='1';
          else
          cVar2S24S74N010P009nsss(0) <='0';
          end if;
        if(cVar1S26S74P064P011P017N054(0)='1' AND  B( 3)='0' AND E( 2)='1' AND A(10)='1' )then
          cVar2S26S74P033P062P018nsss(0) <='1';
          else
          cVar2S26S74P033P062P018nsss(0) <='0';
          end if;
        if(cVar1S27S74P064P011P017N054(0)='1' AND  B( 3)='0' AND E( 2)='0' AND E( 1)='1' )then
          cVar2S27S74P033N062P066nsss(0) <='1';
          else
          cVar2S27S74P033N062P066nsss(0) <='0';
          end if;
        if(cVar1S28S74P064P011N017P009(0)='1' AND  A(12)='1' )then
          cVar2S28S74P014nsss(0) <='1';
          else
          cVar2S28S74P014nsss(0) <='0';
          end if;
        if(cVar1S29S74P064P011N017N009(0)='1' AND  A(11)='1' AND E( 1)='1' )then
          cVar2S29S74P016P066nsss(0) <='1';
          else
          cVar2S29S74P016P066nsss(0) <='0';
          end if;
        if(cVar1S1S75P029P011N051P054(0)='1' AND  E( 5)='0' AND D(11)='0' )then
          cVar2S1S75P050P057nsss(0) <='1';
          else
          cVar2S1S75P050P057nsss(0) <='0';
          end if;
        if(cVar1S2S75P029P011N051P054(0)='1' AND  E( 5)='1' AND D( 3)='1' )then
          cVar2S2S75P050P056nsss(0) <='1';
          else
          cVar2S2S75P050P056nsss(0) <='0';
          end if;
        if(cVar1S3S75P029P011N051N054(0)='1' AND  A(15)='0' AND D( 0)='0' )then
          cVar2S3S75P008P068nsss(0) <='1';
          else
          cVar2S3S75P008P068nsss(0) <='0';
          end if;
        if(cVar1S5S75P029N011P010N052(0)='1' AND  E( 4)='1' )then
          cVar2S5S75P054nsss(0) <='1';
          else
          cVar2S5S75P054nsss(0) <='0';
          end if;
        if(cVar1S6S75P029N011N010P009(0)='1' AND  E( 5)='1' )then
          cVar2S6S75P050nsss(0) <='1';
          else
          cVar2S6S75P050nsss(0) <='0';
          end if;
        if(cVar1S7S75P029N011N010P009(0)='1' AND  E( 5)='0' AND D(12)='1' )then
          cVar2S7S75N050P053nsss(0) <='1';
          else
          cVar2S7S75N050P053nsss(0) <='0';
          end if;
        if(cVar1S8S75P029N011N010P009(0)='1' AND  E( 5)='0' AND D(12)='0' AND E( 4)='1' )then
          cVar2S8S75N050N053P054nsss(0) <='1';
          else
          cVar2S8S75N050N053P054nsss(0) <='0';
          end if;
        if(cVar1S9S75P029N011N010N009(0)='1' AND  A( 2)='1' AND A( 0)='0' )then
          cVar2S9S75P015P019nsss(0) <='1';
          else
          cVar2S9S75P015P019nsss(0) <='0';
          end if;
        if(cVar1S10S75P029N011N010N009(0)='1' AND  A( 2)='0' AND A( 3)='1' )then
          cVar2S10S75N015P013nsss(0) <='1';
          else
          cVar2S10S75N015P013nsss(0) <='0';
          end if;
        if(cVar1S12S75N029P041P020N003(0)='1' AND  A(18)='1' )then
          cVar2S12S75P002nsss(0) <='1';
          else
          cVar2S12S75P002nsss(0) <='0';
          end if;
        if(cVar1S13S75N029P041P020N003(0)='1' AND  A(18)='0' AND A(17)='1' )then
          cVar2S13S75N002P004nsss(0) <='1';
          else
          cVar2S13S75N002P004nsss(0) <='0';
          end if;
        if(cVar1S14S75N029P041P020N003(0)='1' AND  A(18)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S14S75N002N004P005nsss(0) <='1';
          else
          cVar2S14S75N002N004P005nsss(0) <='0';
          end if;
        if(cVar1S15S75N029P041N020P005(0)='1' AND  B( 9)='1' AND D( 7)='0' )then
          cVar2S15S75P021P040nsss(0) <='1';
          else
          cVar2S15S75P021P040nsss(0) <='0';
          end if;
        if(cVar1S16S75N029P041N020P005(0)='1' AND  B( 9)='0' AND B(18)='1' )then
          cVar2S16S75N021P022nsss(0) <='1';
          else
          cVar2S16S75N021P022nsss(0) <='0';
          end if;
        if(cVar1S17S75N029P041N020P005(0)='1' AND  B( 9)='0' AND B(18)='0' AND E( 7)='1' )then
          cVar2S17S75N021N022P042nsss(0) <='1';
          else
          cVar2S17S75N021N022P042nsss(0) <='0';
          end if;
        if(cVar1S18S75N029P041N020N005(0)='1' AND  A( 9)='1' )then
          cVar2S18S75P001nsss(0) <='1';
          else
          cVar2S18S75P001nsss(0) <='0';
          end if;
        if(cVar1S19S75N029P041N020N005(0)='1' AND  A( 9)='0' AND B( 0)='0' AND B( 3)='1' )then
          cVar2S19S75N001P039P033nsss(0) <='1';
          else
          cVar2S19S75N001P039P033nsss(0) <='0';
          end if;
        if(cVar1S21S75N029N041P045N023(0)='1' AND  B(18)='1' )then
          cVar2S21S75P022nsss(0) <='1';
          else
          cVar2S21S75P022nsss(0) <='0';
          end if;
        if(cVar1S22S75N029N041P045N023(0)='1' AND  B(18)='0' AND B(17)='1' )then
          cVar2S22S75N022P024nsss(0) <='1';
          else
          cVar2S22S75N022P024nsss(0) <='0';
          end if;
        if(cVar1S23S75N029N041P045N023(0)='1' AND  B(18)='0' AND B(17)='0' AND B(11)='1' )then
          cVar2S23S75N022N024P036nsss(0) <='1';
          else
          cVar2S23S75N022N024P036nsss(0) <='0';
          end if;
        if(cVar1S24S75N029N041N045P027(0)='1' AND  D(13)='1' )then
          cVar2S24S75P049nsss(0) <='1';
          else
          cVar2S24S75P049nsss(0) <='0';
          end if;
        if(cVar1S25S75N029N041N045P027(0)='1' AND  D(13)='0' AND E( 1)='0' AND A( 5)='1' )then
          cVar2S25S75N049P066P009nsss(0) <='1';
          else
          cVar2S25S75N049P066P009nsss(0) <='0';
          end if;
        if(cVar1S26S75N029N041N045N027(0)='1' AND  B(15)='1' AND A(14)='1' AND B( 4)='0' )then
          cVar2S26S75P028P010P031nsss(0) <='1';
          else
          cVar2S26S75P028P010P031nsss(0) <='0';
          end if;
        if(cVar1S27S75N029N041N045N027(0)='1' AND  B(15)='0' AND D( 7)='1' AND B( 9)='1' )then
          cVar2S27S75N028P040P021nsss(0) <='1';
          else
          cVar2S27S75N028P040P021nsss(0) <='0';
          end if;
        if(cVar1S0S76P064P027P066P009(0)='1' AND  E( 5)='1' AND A( 3)='0' )then
          cVar2S0S76P050P013nsss(0) <='1';
          else
          cVar2S0S76P050P013nsss(0) <='0';
          end if;
        if(cVar1S1S76P064P027P066P009(0)='1' AND  E( 5)='0' AND A( 1)='0' )then
          cVar2S1S76N050P017nsss(0) <='1';
          else
          cVar2S1S76N050P017nsss(0) <='0';
          end if;
        if(cVar1S2S76P064P027P066N009(0)='1' AND  B( 3)='0' )then
          cVar2S2S76P033nsss(0) <='1';
          else
          cVar2S2S76P033nsss(0) <='0';
          end if;
        if(cVar1S4S76P064P027P066P068(0)='1' AND  A( 3)='1' )then
          cVar2S4S76P013nsss(0) <='1';
          else
          cVar2S4S76P013nsss(0) <='0';
          end if;
        if(cVar1S5S76P064P027P066P068(0)='1' AND  A( 3)='0' AND E( 5)='1' )then
          cVar2S5S76N013P050nsss(0) <='1';
          else
          cVar2S5S76N013P050nsss(0) <='0';
          end if;
        if(cVar1S6S76P064N027P041P020(0)='1' AND  A( 8)='1' )then
          cVar2S6S76P003nsss(0) <='1';
          else
          cVar2S6S76P003nsss(0) <='0';
          end if;
        if(cVar1S7S76P064N027P041P020(0)='1' AND  A( 8)='0' AND A(18)='1' )then
          cVar2S7S76N003P002nsss(0) <='1';
          else
          cVar2S7S76N003P002nsss(0) <='0';
          end if;
        if(cVar1S8S76P064N027P041P020(0)='1' AND  A( 8)='0' AND A(18)='0' AND A( 0)='0' )then
          cVar2S8S76N003N002P019nsss(0) <='1';
          else
          cVar2S8S76N003N002P019nsss(0) <='0';
          end if;
        if(cVar1S9S76P064N027P041N020(0)='1' AND  A( 7)='1' AND D( 7)='0' )then
          cVar2S9S76P005P040nsss(0) <='1';
          else
          cVar2S9S76P005P040nsss(0) <='0';
          end if;
        if(cVar1S10S76P064N027P041N020(0)='1' AND  A( 7)='0' AND A( 9)='1' )then
          cVar2S10S76N005P001nsss(0) <='1';
          else
          cVar2S10S76N005P001nsss(0) <='0';
          end if;
        if(cVar1S11S76P064N027P041N020(0)='1' AND  A( 7)='0' AND A( 9)='0' AND B(18)='1' )then
          cVar2S11S76N005N001P022nsss(0) <='1';
          else
          cVar2S11S76N005N001P022nsss(0) <='0';
          end if;
        if(cVar1S12S76P064N027N041P039(0)='1' AND  B(12)='1' AND E(10)='1' AND A(16)='0' )then
          cVar2S12S76P034P063P006nsss(0) <='1';
          else
          cVar2S12S76P034P063P006nsss(0) <='0';
          end if;
        if(cVar1S13S76P064N027N041P039(0)='1' AND  B(12)='1' AND E(10)='0' AND E( 2)='1' )then
          cVar2S13S76P034N063P062nsss(0) <='1';
          else
          cVar2S13S76P034N063P062nsss(0) <='0';
          end if;
        if(cVar1S14S76P064N027N041P039(0)='1' AND  B(12)='0' AND E(10)='0' AND A( 1)='0' )then
          cVar2S14S76N034P063P017nsss(0) <='1';
          else
          cVar2S14S76N034P063P017nsss(0) <='0';
          end if;
        if(cVar1S15S76P064N027N041P039(0)='1' AND  B(12)='0' AND E(10)='1' AND B(11)='1' )then
          cVar2S15S76N034P063P036nsss(0) <='1';
          else
          cVar2S15S76N034P063P036nsss(0) <='0';
          end if;
        if(cVar1S16S76P064N027N041P039(0)='1' AND  E( 7)='1' )then
          cVar2S16S76P042nsss(0) <='1';
          else
          cVar2S16S76P042nsss(0) <='0';
          end if;
        if(cVar1S17S76P064N027N041P039(0)='1' AND  E( 7)='0' AND B( 3)='1' )then
          cVar2S17S76N042P033nsss(0) <='1';
          else
          cVar2S17S76N042P033nsss(0) <='0';
          end if;
        if(cVar1S19S76P064N042P008P027(0)='1' AND  E( 6)='1' )then
          cVar2S19S76P046nsss(0) <='1';
          else
          cVar2S19S76P046nsss(0) <='0';
          end if;
        if(cVar1S20S76P064N042P008P027(0)='1' AND  E( 6)='0' AND B(12)='0' AND D( 0)='0' )then
          cVar2S20S76N046P034P068nsss(0) <='1';
          else
          cVar2S20S76N046P034P068nsss(0) <='0';
          end if;
        if(cVar1S21S76P064N042P008P027(0)='1' AND  E( 6)='0' AND B(12)='1' AND A(12)='1' )then
          cVar2S21S76N046P034P014nsss(0) <='1';
          else
          cVar2S21S76N046P034P014nsss(0) <='0';
          end if;
        if(cVar1S22S76P064N042P008P027(0)='1' AND  A(12)='1' )then
          cVar2S22S76P014nsss(0) <='1';
          else
          cVar2S22S76P014nsss(0) <='0';
          end if;
        if(cVar1S23S76P064N042P008P010(0)='1' AND  A( 0)='1' AND A(11)='0' )then
          cVar2S23S76P019P016nsss(0) <='1';
          else
          cVar2S23S76P019P016nsss(0) <='0';
          end if;
        if(cVar1S24S76P064N042P008P010(0)='1' AND  A( 0)='0' AND D( 0)='1' )then
          cVar2S24S76N019P068nsss(0) <='1';
          else
          cVar2S24S76N019P068nsss(0) <='0';
          end if;
        if(cVar1S0S77P017P064P034P035(0)='1' AND  D(11)='0' AND D( 0)='0' AND A( 3)='0' )then
          cVar2S0S77P057P068P013nsss(0) <='1';
          else
          cVar2S0S77P057P068P013nsss(0) <='0';
          end if;
        if(cVar1S1S77P017P064P034P035(0)='1' AND  D(11)='0' AND D( 0)='1' AND A( 3)='1' )then
          cVar2S1S77P057P068P013nsss(0) <='1';
          else
          cVar2S1S77P057P068P013nsss(0) <='0';
          end if;
        if(cVar1S2S77P017P064P034P035(0)='1' AND  A(10)='1' )then
          cVar2S2S77P018nsss(0) <='1';
          else
          cVar2S2S77P018nsss(0) <='0';
          end if;
        if(cVar1S3S77P017P064N034P020(0)='1' AND  E( 9)='1' )then
          cVar2S3S77P067nsss(0) <='1';
          else
          cVar2S3S77P067nsss(0) <='0';
          end if;
        if(cVar1S4S77P017P064N034P020(0)='1' AND  E( 9)='0' AND A( 8)='1' )then
          cVar2S4S77N067P003nsss(0) <='1';
          else
          cVar2S4S77N067P003nsss(0) <='0';
          end if;
        if(cVar1S5S77P017P064N034P020(0)='1' AND  E( 9)='0' AND A( 8)='0' AND B( 1)='0' )then
          cVar2S5S77N067N003P037nsss(0) <='1';
          else
          cVar2S5S77N067N003P037nsss(0) <='0';
          end if;
        if(cVar1S6S77P017P064N034N020(0)='1' AND  B( 0)='0' AND A(11)='1' AND E(10)='0' )then
          cVar2S6S77P039P016P063nsss(0) <='1';
          else
          cVar2S6S77P039P016P063nsss(0) <='0';
          end if;
        if(cVar1S7S77P017P064N034N020(0)='1' AND  B( 0)='0' AND A(11)='0' AND A(18)='0' )then
          cVar2S7S77P039N016P002nsss(0) <='1';
          else
          cVar2S7S77P039N016P002nsss(0) <='0';
          end if;
        if(cVar1S8S77P017P064N034N020(0)='1' AND  B( 0)='1' AND A( 2)='1' )then
          cVar2S8S77P039P015nsss(0) <='1';
          else
          cVar2S8S77P039P015nsss(0) <='0';
          end if;
        if(cVar1S10S77P017P064N050P020(0)='1' AND  A( 2)='0' AND D( 4)='0' AND E(12)='0' )then
          cVar2S10S77P015P052P055nsss(0) <='1';
          else
          cVar2S10S77P015P052P055nsss(0) <='0';
          end if;
        if(cVar1S11S77P017P064N050P020(0)='1' AND  A( 2)='1' AND A(10)='1' AND D( 9)='1' )then
          cVar2S11S77P015P018P065nsss(0) <='1';
          else
          cVar2S11S77P015P018P065nsss(0) <='0';
          end if;
        if(cVar1S12S77P017P064N050P020(0)='1' AND  A( 2)='1' AND A(10)='0' AND B( 3)='1' )then
          cVar2S12S77P015N018P033nsss(0) <='1';
          else
          cVar2S12S77P015N018P033nsss(0) <='0';
          end if;
        if(cVar1S14S77N017P041P020N003(0)='1' AND  A(18)='1' )then
          cVar2S14S77P002nsss(0) <='1';
          else
          cVar2S14S77P002nsss(0) <='0';
          end if;
        if(cVar1S15S77N017P041P020N003(0)='1' AND  A(18)='0' AND A(17)='1' )then
          cVar2S15S77N002P004nsss(0) <='1';
          else
          cVar2S15S77N002P004nsss(0) <='0';
          end if;
        if(cVar1S16S77N017P041N020P015(0)='1' AND  B( 0)='1' )then
          cVar2S16S77P039nsss(0) <='1';
          else
          cVar2S16S77P039nsss(0) <='0';
          end if;
        if(cVar1S17S77N017P041N020P015(0)='1' AND  B( 0)='0' AND E(15)='1' )then
          cVar2S17S77N039P043nsss(0) <='1';
          else
          cVar2S17S77N039P043nsss(0) <='0';
          end if;
        if(cVar1S18S77N017P041N020P015(0)='1' AND  B( 0)='0' AND E(15)='0' AND A(11)='1' )then
          cVar2S18S77N039N043P016nsss(0) <='1';
          else
          cVar2S18S77N039N043P016nsss(0) <='0';
          end if;
        if(cVar1S19S77N017P041N020P015(0)='1' AND  A( 0)='1' )then
          cVar2S19S77P019nsss(0) <='1';
          else
          cVar2S19S77P019nsss(0) <='0';
          end if;
        if(cVar1S20S77N017N041P062P027(0)='1' AND  A( 5)='1' )then
          cVar2S20S77P009nsss(0) <='1';
          else
          cVar2S20S77P009nsss(0) <='0';
          end if;
        if(cVar1S21S77N017N041P062P027(0)='1' AND  A( 5)='0' AND A(15)='1' )then
          cVar2S21S77N009P008nsss(0) <='1';
          else
          cVar2S21S77N009P008nsss(0) <='0';
          end if;
        if(cVar1S22S77N017N041P062P027(0)='1' AND  A( 5)='0' AND A(15)='0' AND A(16)='1' )then
          cVar2S22S77N009N008P006nsss(0) <='1';
          else
          cVar2S22S77N009N008P006nsss(0) <='0';
          end if;
        if(cVar1S23S77N017N041P062N027(0)='1' AND  B( 8)='1' AND E( 7)='1' AND A(15)='0' )then
          cVar2S23S77P023P042P008nsss(0) <='1';
          else
          cVar2S23S77P023P042P008nsss(0) <='0';
          end if;
        if(cVar1S24S77N017N041P062N027(0)='1' AND  B( 8)='1' AND E( 7)='0' AND B( 1)='0' )then
          cVar2S24S77P023N042P037nsss(0) <='1';
          else
          cVar2S24S77P023N042P037nsss(0) <='0';
          end if;
        if(cVar1S25S77N017N041P062N027(0)='1' AND  B( 8)='0' AND A( 3)='1' AND B( 4)='1' )then
          cVar2S25S77N023P013P031nsss(0) <='1';
          else
          cVar2S25S77N023P013P031nsss(0) <='0';
          end if;
        if(cVar1S26S77N017N041P062N027(0)='1' AND  B( 8)='0' AND A( 3)='0' AND D( 9)='1' )then
          cVar2S26S77N023N013P065nsss(0) <='1';
          else
          cVar2S26S77N023N013P065nsss(0) <='0';
          end if;
        if(cVar1S27S77N017N041P062P010(0)='1' AND  A( 8)='0' AND D( 4)='1' )then
          cVar2S27S77P003P052nsss(0) <='1';
          else
          cVar2S27S77P003P052nsss(0) <='0';
          end if;
        if(cVar1S28S77N017N041P062P010(0)='1' AND  A( 8)='0' AND D( 4)='0' AND A(11)='1' )then
          cVar2S28S77P003N052P016nsss(0) <='1';
          else
          cVar2S28S77P003N052P016nsss(0) <='0';
          end if;
        if(cVar1S29S77N017N041P062P010(0)='1' AND  A( 8)='1' AND B(12)='0' AND A( 3)='1' )then
          cVar2S29S77P003N034P013nsss(0) <='1';
          else
          cVar2S29S77P003N034P013nsss(0) <='0';
          end if;
        if(cVar1S30S77N017N041P062P010(0)='1' AND  A(15)='0' AND E( 3)='1' )then
          cVar2S30S77P008P058nsss(0) <='1';
          else
          cVar2S30S77P008P058nsss(0) <='0';
          end if;
        if(cVar1S0S78P062P063P007P025(0)='1' AND  D(13)='1' )then
          cVar2S0S78P049nsss(0) <='1';
          else
          cVar2S0S78P049nsss(0) <='0';
          end if;
        if(cVar1S1S78P062P063P007P025(0)='1' AND  D(13)='0' AND E( 1)='0' )then
          cVar2S1S78N049P066nsss(0) <='1';
          else
          cVar2S1S78N049P066nsss(0) <='0';
          end if;
        if(cVar1S2S78P062P063P007N025(0)='1' AND  A( 4)='0' AND D( 0)='0' )then
          cVar2S2S78P011P068nsss(0) <='1';
          else
          cVar2S2S78P011P068nsss(0) <='0';
          end if;
        if(cVar1S3S78P062P063P007N025(0)='1' AND  A( 4)='0' AND D( 0)='1' AND A( 0)='1' )then
          cVar2S3S78P011P068P019nsss(0) <='1';
          else
          cVar2S3S78P011P068P019nsss(0) <='0';
          end if;
        if(cVar1S4S78P062P063P007N025(0)='1' AND  A( 4)='1' AND A( 2)='1' AND A( 8)='1' )then
          cVar2S4S78P011P015P003nsss(0) <='1';
          else
          cVar2S4S78P011P015P003nsss(0) <='0';
          end if;
        if(cVar1S5S78P062P063P007N025(0)='1' AND  A( 4)='1' AND A( 2)='0' AND A(13)='1' )then
          cVar2S5S78P011N015P012nsss(0) <='1';
          else
          cVar2S5S78P011N015P012nsss(0) <='0';
          end if;
        if(cVar1S6S78P062P063N007P029(0)='1' AND  A( 4)='1' AND B( 3)='0' )then
          cVar2S6S78P011P033nsss(0) <='1';
          else
          cVar2S6S78P011P033nsss(0) <='0';
          end if;
        if(cVar1S7S78P062P063N007P029(0)='1' AND  A( 4)='0' AND A( 2)='1' AND A( 3)='0' )then
          cVar2S7S78N011P015P013nsss(0) <='1';
          else
          cVar2S7S78N011P015P013nsss(0) <='0';
          end if;
        if(cVar1S8S78P062P063N007P029(0)='1' AND  A( 4)='0' AND A( 2)='0' AND A(10)='0' )then
          cVar2S8S78N011N015P018nsss(0) <='1';
          else
          cVar2S8S78N011N015P018nsss(0) <='0';
          end if;
        if(cVar1S9S78P062P063N007N029(0)='1' AND  B(15)='1' AND D(12)='1' AND A(13)='0' )then
          cVar2S9S78P028P053P012nsss(0) <='1';
          else
          cVar2S9S78P028P053P012nsss(0) <='0';
          end if;
        if(cVar1S10S78P062P063N007N029(0)='1' AND  B(15)='1' AND D(12)='0' AND E( 4)='1' )then
          cVar2S10S78P028N053P054nsss(0) <='1';
          else
          cVar2S10S78P028N053P054nsss(0) <='0';
          end if;
        if(cVar1S11S78P062P063N007N029(0)='1' AND  B(15)='0' AND B(16)='1' )then
          cVar2S11S78N028P026nsss(0) <='1';
          else
          cVar2S11S78N028P026nsss(0) <='0';
          end if;
        if(cVar1S12S78P062P063N007N029(0)='1' AND  B(15)='0' AND B(16)='0' AND E(13)='0' )then
          cVar2S12S78N028N026P051nsss(0) <='1';
          else
          cVar2S12S78N028N026P051nsss(0) <='0';
          end if;
        if(cVar1S13S78P062P063P035P058(0)='1' AND  B(11)='0' AND B(12)='0' )then
          cVar2S13S78P036P034nsss(0) <='1';
          else
          cVar2S13S78P036P034nsss(0) <='0';
          end if;
        if(cVar1S14S78P062P063P035P058(0)='1' AND  B(11)='0' AND B(12)='1' AND A(11)='1' )then
          cVar2S14S78P036P034P016nsss(0) <='1';
          else
          cVar2S14S78P036P034P016nsss(0) <='0';
          end if;
        if(cVar1S15S78P062P063P035P058(0)='1' AND  B(11)='1' AND A(11)='1' )then
          cVar2S15S78P036P016nsss(0) <='1';
          else
          cVar2S15S78P036P016nsss(0) <='0';
          end if;
        if(cVar1S16S78P062P063N035P034(0)='1' AND  D( 1)='0' AND A(16)='0' AND B( 4)='0' )then
          cVar2S16S78P064P006P031nsss(0) <='1';
          else
          cVar2S16S78P064P006P031nsss(0) <='0';
          end if;
        if(cVar1S17S78P062P063N035P034(0)='1' AND  D( 1)='1' AND A(12)='1' )then
          cVar2S17S78P064P014nsss(0) <='1';
          else
          cVar2S17S78P064P014nsss(0) <='0';
          end if;
        if(cVar1S18S78P062P063N035N034(0)='1' AND  B(11)='1' AND A( 6)='0' AND A( 2)='0' )then
          cVar2S18S78P036P007P015nsss(0) <='1';
          else
          cVar2S18S78P036P007P015nsss(0) <='0';
          end if;
        if(cVar1S19S78P062P063N035N034(0)='1' AND  B(11)='0' AND D( 9)='0' AND E( 1)='1' )then
          cVar2S19S78N036P065P066nsss(0) <='1';
          else
          cVar2S19S78N036P065P066nsss(0) <='0';
          end if;
        if(cVar1S20S78P062P063N035N034(0)='1' AND  B(11)='0' AND D( 9)='1' AND B( 1)='1' )then
          cVar2S20S78N036P065P037nsss(0) <='1';
          else
          cVar2S20S78N036P065P037nsss(0) <='0';
          end if;
        if(cVar1S21S78P062P026P027P060(0)='1' AND  D( 1)='0' AND A(14)='0' )then
          cVar2S21S78P064P010nsss(0) <='1';
          else
          cVar2S21S78P064P010nsss(0) <='0';
          end if;
        if(cVar1S22S78P062P026P027P060(0)='1' AND  D( 1)='1' AND D( 0)='1' )then
          cVar2S22S78P064P068nsss(0) <='1';
          else
          cVar2S22S78P064P068nsss(0) <='0';
          end if;
        if(cVar1S23S78P062P026P027P060(0)='1' AND  D( 1)='1' AND D( 0)='0' AND D(10)='1' )then
          cVar2S23S78P064N068P061nsss(0) <='1';
          else
          cVar2S23S78P064N068P061nsss(0) <='0';
          end if;
        if(cVar1S24S78P062P026P027N060(0)='1' AND  D( 1)='1' AND E(11)='0' AND A(12)='1' )then
          cVar2S24S78P064P059P014nsss(0) <='1';
          else
          cVar2S24S78P064P059P014nsss(0) <='0';
          end if;
        if(cVar1S25S78P062P026P027N060(0)='1' AND  D( 1)='1' AND E(11)='1' AND E(10)='1' )then
          cVar2S25S78P064P059P063nsss(0) <='1';
          else
          cVar2S25S78P064P059P063nsss(0) <='0';
          end if;
        if(cVar1S26S78P062P026P027N060(0)='1' AND  D( 1)='0' AND D( 4)='1' )then
          cVar2S26S78N064P052nsss(0) <='1';
          else
          cVar2S26S78N064P052nsss(0) <='0';
          end if;
        if(cVar1S27S78P062P026P027N060(0)='1' AND  D( 1)='0' AND D( 4)='0' AND E(13)='1' )then
          cVar2S27S78N064N052P051nsss(0) <='1';
          else
          cVar2S27S78N064N052P051nsss(0) <='0';
          end if;
        if(cVar1S1S79P051P008P065N028(0)='1' AND  B(16)='1' AND D( 0)='0' )then
          cVar2S1S79P026P068nsss(0) <='1';
          else
          cVar2S1S79P026P068nsss(0) <='0';
          end if;
        if(cVar1S2S79P051P008P065N028(0)='1' AND  B(16)='0' AND D(12)='1' )then
          cVar2S2S79N026P053nsss(0) <='1';
          else
          cVar2S2S79N026P053nsss(0) <='0';
          end if;
        if(cVar1S4S79P051N008N042P009(0)='1' AND  D(12)='1' AND B( 5)='1' )then
          cVar2S4S79P053P029nsss(0) <='1';
          else
          cVar2S4S79P053P029nsss(0) <='0';
          end if;
        if(cVar1S5S79P051N008N042P009(0)='1' AND  D(12)='1' AND B( 5)='0' AND D( 4)='0' )then
          cVar2S5S79P053N029P052nsss(0) <='1';
          else
          cVar2S5S79P053N029P052nsss(0) <='0';
          end if;
        if(cVar1S6S79P051N008N042P009(0)='1' AND  D(12)='0' AND D(13)='1' )then
          cVar2S6S79N053P049nsss(0) <='1';
          else
          cVar2S6S79N053P049nsss(0) <='0';
          end if;
        if(cVar1S7S79P051N008N042N009(0)='1' AND  A( 4)='1' AND D(12)='1' AND A(13)='0' )then
          cVar2S7S79P011P053P012nsss(0) <='1';
          else
          cVar2S7S79P011P053P012nsss(0) <='0';
          end if;
        if(cVar1S8S79P051N008N042N009(0)='1' AND  A( 4)='0' AND A( 6)='1' )then
          cVar2S8S79N011P007nsss(0) <='1';
          else
          cVar2S8S79N011P007nsss(0) <='0';
          end if;
        if(cVar1S9S79P051N008N042N009(0)='1' AND  A( 4)='0' AND A( 6)='0' AND B(12)='1' )then
          cVar2S9S79N011N007P034nsss(0) <='1';
          else
          cVar2S9S79N011N007P034nsss(0) <='0';
          end if;
        if(cVar1S11S79N051P041P020N003(0)='1' AND  A(18)='1' )then
          cVar2S11S79P002nsss(0) <='1';
          else
          cVar2S11S79P002nsss(0) <='0';
          end if;
        if(cVar1S12S79N051P041P020N003(0)='1' AND  A(18)='0' AND A( 7)='1' )then
          cVar2S12S79N002P005nsss(0) <='1';
          else
          cVar2S12S79N002P005nsss(0) <='0';
          end if;
        if(cVar1S13S79N051P041P020N003(0)='1' AND  A(18)='0' AND A( 7)='0' AND A(17)='1' )then
          cVar2S13S79N002N005P004nsss(0) <='1';
          else
          cVar2S13S79N002N005P004nsss(0) <='0';
          end if;
        if(cVar1S15S79N051P041N020N001(0)='1' AND  B( 9)='1' AND A( 7)='1' AND D( 7)='0' )then
          cVar2S15S79P021P005P040nsss(0) <='1';
          else
          cVar2S15S79P021P005P040nsss(0) <='0';
          end if;
        if(cVar1S16S79N051P041N020N001(0)='1' AND  B( 9)='1' AND A( 7)='0' )then
          cVar2S16S79P021N005psss(0) <='1';
          else
          cVar2S16S79P021N005psss(0) <='0';
          end if;
        if(cVar1S17S79N051P041N020N001(0)='1' AND  B( 9)='0' AND B( 0)='0' AND E( 9)='1' )then
          cVar2S17S79N021P039P067nsss(0) <='1';
          else
          cVar2S17S79N021P039P067nsss(0) <='0';
          end if;
        if(cVar1S18S79N051N041P047P026(0)='1' AND  A( 5)='1' )then
          cVar2S18S79P009nsss(0) <='1';
          else
          cVar2S18S79P009nsss(0) <='0';
          end if;
        if(cVar1S19S79N051N041P047P026(0)='1' AND  A( 5)='0' AND B(17)='0' AND A(13)='0' )then
          cVar2S19S79N009P024P012nsss(0) <='1';
          else
          cVar2S19S79N009P024P012nsss(0) <='0';
          end if;
        if(cVar1S20S79N051N041P047N026(0)='1' AND  B(17)='1' AND A(16)='1' AND A(15)='0' )then
          cVar2S20S79P024P006P008nsss(0) <='1';
          else
          cVar2S20S79P024P006P008nsss(0) <='0';
          end if;
        if(cVar1S21S79N051N041P047N026(0)='1' AND  B(17)='1' AND A(16)='0' )then
          cVar2S21S79P024N006psss(0) <='1';
          else
          cVar2S21S79P024N006psss(0) <='0';
          end if;
        if(cVar1S22S79N051N041P047N026(0)='1' AND  B(17)='0' AND B( 6)='1' )then
          cVar2S22S79N024P027nsss(0) <='1';
          else
          cVar2S22S79N024P027nsss(0) <='0';
          end if;
        if(cVar1S23S79N051N041P047N026(0)='1' AND  B(17)='0' AND B( 6)='0' AND B( 7)='1' )then
          cVar2S23S79N024N027P025nsss(0) <='1';
          else
          cVar2S23S79N024N027P025nsss(0) <='0';
          end if;
        if(cVar1S24S79N051N041N047P049(0)='1' AND  B(13)='1' AND A( 4)='0' AND A( 0)='0' )then
          cVar2S24S79P032P011P019nsss(0) <='1';
          else
          cVar2S24S79P032P011P019nsss(0) <='0';
          end if;
        if(cVar1S25S79N051N041N047P049(0)='1' AND  B(13)='1' AND A( 4)='1' AND D(11)='1' )then
          cVar2S25S79P032P011P057nsss(0) <='1';
          else
          cVar2S25S79P032P011P057nsss(0) <='0';
          end if;
        if(cVar1S26S79N051N041N047P049(0)='1' AND  B(13)='0' AND B(15)='1' AND A(14)='1' )then
          cVar2S26S79N032P028P010nsss(0) <='1';
          else
          cVar2S26S79N032P028P010nsss(0) <='0';
          end if;
        if(cVar1S27S79N051N041N047P049(0)='1' AND  B(12)='1' )then
          cVar2S27S79P034nsss(0) <='1';
          else
          cVar2S27S79P034nsss(0) <='0';
          end if;
        if(cVar1S28S79N051N041N047P049(0)='1' AND  B(12)='0' AND B( 3)='1' )then
          cVar2S28S79N034P033nsss(0) <='1';
          else
          cVar2S28S79N034P033nsss(0) <='0';
          end if;
        if(cVar1S29S79N051N041N047P049(0)='1' AND  B(12)='0' AND B( 3)='0' AND B( 2)='1' )then
          cVar2S29S79N034N033P035nsss(0) <='1';
          else
          cVar2S29S79N034N033P035nsss(0) <='0';
          end if;
        if(cVar1S2S80P040P002N021N041(0)='1' AND  B(10)='1' )then
          cVar2S2S80P038nsss(0) <='1';
          else
          cVar2S2S80P038nsss(0) <='0';
          end if;
        if(cVar1S4S80P040N002N057P004(0)='1' AND  B( 8)='1' )then
          cVar2S4S80P023nsss(0) <='1';
          else
          cVar2S4S80P023nsss(0) <='0';
          end if;
        if(cVar1S5S80P040N002N057P004(0)='1' AND  B( 8)='0' AND B(18)='1' )then
          cVar2S5S80N023P022nsss(0) <='1';
          else
          cVar2S5S80N023P022nsss(0) <='0';
          end if;
        if(cVar1S6S80P040N002N057P004(0)='1' AND  B( 8)='0' AND B(18)='0' AND B(10)='1' )then
          cVar2S6S80N023N022P038nsss(0) <='1';
          else
          cVar2S6S80N023N022P038nsss(0) <='0';
          end if;
        if(cVar1S7S80P040N002N057N004(0)='1' AND  A(19)='1' )then
          cVar2S7S80P000nsss(0) <='1';
          else
          cVar2S7S80P000nsss(0) <='0';
          end if;
        if(cVar1S8S80P040N002N057N004(0)='1' AND  A(19)='0' AND E( 5)='1' )then
          cVar2S8S80N000P050nsss(0) <='1';
          else
          cVar2S8S80N000P050nsss(0) <='0';
          end if;
        if(cVar1S9S80P040N002N057N004(0)='1' AND  A(19)='0' AND E( 5)='0' AND A( 7)='1' )then
          cVar2S9S80N000N050P005nsss(0) <='1';
          else
          cVar2S9S80N000N050P005nsss(0) <='0';
          end if;
        if(cVar1S10S80N040P021P007P025(0)='1' AND  E( 1)='0' )then
          cVar2S10S80P066nsss(0) <='1';
          else
          cVar2S10S80P066nsss(0) <='0';
          end if;
        if(cVar1S11S80N040P021P007P025(0)='1' AND  E( 1)='1' AND A(10)='0' )then
          cVar2S11S80P066P018nsss(0) <='1';
          else
          cVar2S11S80P066P018nsss(0) <='0';
          end if;
        if(cVar1S12S80N040P021P007N025(0)='1' AND  E(12)='0' )then
          cVar2S12S80P055nsss(0) <='1';
          else
          cVar2S12S80P055nsss(0) <='0';
          end if;
        if(cVar1S13S80N040P021P007N025(0)='1' AND  E(12)='1' AND A(14)='1' )then
          cVar2S13S80P055P010nsss(0) <='1';
          else
          cVar2S13S80P055P010nsss(0) <='0';
          end if;
        if(cVar1S14S80N040P021N007P028(0)='1' AND  D(12)='1' AND D( 1)='0' AND A(13)='0' )then
          cVar2S14S80P053P064P012nsss(0) <='1';
          else
          cVar2S14S80P053P064P012nsss(0) <='0';
          end if;
        if(cVar1S15S80N040P021N007P028(0)='1' AND  D(12)='0' AND A(18)='0' AND A( 7)='0' )then
          cVar2S15S80N053P002P005nsss(0) <='1';
          else
          cVar2S15S80N053P002P005nsss(0) <='0';
          end if;
        if(cVar1S16S80N040P021N007N028(0)='1' AND  B( 5)='1' AND A( 4)='1' AND E( 3)='0' )then
          cVar2S16S80P029P011P058nsss(0) <='1';
          else
          cVar2S16S80P029P011P058nsss(0) <='0';
          end if;
        if(cVar1S17S80N040P021N007N028(0)='1' AND  B( 5)='1' AND A( 4)='0' AND E(10)='0' )then
          cVar2S17S80P029N011P063nsss(0) <='1';
          else
          cVar2S17S80P029N011P063nsss(0) <='0';
          end if;
        if(cVar1S18S80N040P021N007N028(0)='1' AND  B( 5)='0' AND E( 2)='1' AND B( 6)='0' )then
          cVar2S18S80N029P062P027nsss(0) <='1';
          else
          cVar2S18S80N029P062P027nsss(0) <='0';
          end if;
        if(cVar1S19S80N040P021N007N028(0)='1' AND  B( 5)='0' AND E( 2)='0' )then
          cVar2S19S80N029N062psss(0) <='1';
          else
          cVar2S19S80N029N062psss(0) <='0';
          end if;
        if(cVar1S21S80N040P021N042P003(0)='1' AND  A( 0)='1' )then
          cVar2S21S80P019nsss(0) <='1';
          else
          cVar2S21S80P019nsss(0) <='0';
          end if;
        if(cVar1S22S80N040P021N042P003(0)='1' AND  A( 0)='0' AND B( 0)='1' )then
          cVar2S22S80N019P039nsss(0) <='1';
          else
          cVar2S22S80N019P039nsss(0) <='0';
          end if;
        if(cVar1S23S80N040P021N042N003(0)='1' AND  A(15)='1' AND A( 2)='1' )then
          cVar2S23S80P008P015nsss(0) <='1';
          else
          cVar2S23S80P008P015nsss(0) <='0';
          end if;
        if(cVar1S24S80N040P021N042N003(0)='1' AND  A(15)='0' AND A( 2)='1' AND E( 1)='1' )then
          cVar2S24S80N008P015P066nsss(0) <='1';
          else
          cVar2S24S80N008P015P066nsss(0) <='0';
          end if;
        if(cVar1S2S81P040N002N057P004(0)='1' AND  B( 8)='1' )then
          cVar2S2S81P023nsss(0) <='1';
          else
          cVar2S2S81P023nsss(0) <='0';
          end if;
        if(cVar1S3S81P040N002N057P004(0)='1' AND  B( 8)='0' AND B(18)='1' )then
          cVar2S3S81N023P022nsss(0) <='1';
          else
          cVar2S3S81N023P022nsss(0) <='0';
          end if;
        if(cVar1S4S81P040N002N057P004(0)='1' AND  B( 8)='0' AND B(18)='0' AND B(10)='1' )then
          cVar2S4S81N023N022P038nsss(0) <='1';
          else
          cVar2S4S81N023N022P038nsss(0) <='0';
          end if;
        if(cVar1S5S81P040N002N057N004(0)='1' AND  B(19)='0' AND A( 2)='0' )then
          cVar2S5S81P020P015nsss(0) <='1';
          else
          cVar2S5S81P020P015nsss(0) <='0';
          end if;
        if(cVar1S6S81N040P028P029P053(0)='1' AND  A(12)='0' )then
          cVar2S6S81P014nsss(0) <='1';
          else
          cVar2S6S81P014nsss(0) <='0';
          end if;
        if(cVar1S7S81N040P028P029P053(0)='1' AND  A(12)='1' AND A(14)='1' )then
          cVar2S7S81P014P010nsss(0) <='1';
          else
          cVar2S7S81P014P010nsss(0) <='0';
          end if;
        if(cVar1S8S81N040P028P029N053(0)='1' AND  D( 0)='0' AND B( 4)='0' )then
          cVar2S8S81P068P031nsss(0) <='1';
          else
          cVar2S8S81P068P031nsss(0) <='0';
          end if;
        if(cVar1S9S81N040P028P029N053(0)='1' AND  D( 0)='1' AND A(10)='1' AND B( 1)='1' )then
          cVar2S9S81P068P018P037nsss(0) <='1';
          else
          cVar2S9S81P068P018P037nsss(0) <='0';
          end if;
        if(cVar1S10S81N040N028P029P011(0)='1' AND  E( 4)='1' AND D(11)='0' AND E( 5)='0' )then
          cVar2S10S81P054P057P050nsss(0) <='1';
          else
          cVar2S10S81P054P057P050nsss(0) <='0';
          end if;
        if(cVar1S11S81N040N028P029P011(0)='1' AND  E( 4)='0' AND D(12)='1' )then
          cVar2S11S81N054P053nsss(0) <='1';
          else
          cVar2S11S81N054P053nsss(0) <='0';
          end if;
        if(cVar1S12S81N040N028P029P011(0)='1' AND  E( 4)='0' AND D(12)='0' AND D( 4)='1' )then
          cVar2S12S81N054N053P052nsss(0) <='1';
          else
          cVar2S12S81N054N053P052nsss(0) <='0';
          end if;
        if(cVar1S13S81N040N028P029N011(0)='1' AND  A(14)='1' AND D( 4)='1' )then
          cVar2S13S81P010P052nsss(0) <='1';
          else
          cVar2S13S81P010P052nsss(0) <='0';
          end if;
        if(cVar1S14S81N040N028P029N011(0)='1' AND  A(14)='1' AND D( 4)='0' AND E( 4)='1' )then
          cVar2S14S81P010N052P054nsss(0) <='1';
          else
          cVar2S14S81P010N052P054nsss(0) <='0';
          end if;
        if(cVar1S15S81N040N028P029N011(0)='1' AND  A(14)='0' AND A( 5)='1' )then
          cVar2S15S81N010P009nsss(0) <='1';
          else
          cVar2S15S81N010P009nsss(0) <='0';
          end if;
        if(cVar1S16S81N040N028P029N011(0)='1' AND  A(14)='0' AND A( 5)='0' AND A( 3)='1' )then
          cVar2S16S81N010N009P013nsss(0) <='1';
          else
          cVar2S16S81N010N009P013nsss(0) <='0';
          end if;
        if(cVar1S17S81N040N028N029P007(0)='1' AND  B( 7)='1' AND A(15)='0' )then
          cVar2S17S81P025P008nsss(0) <='1';
          else
          cVar2S17S81P025P008nsss(0) <='0';
          end if;
        if(cVar1S18S81N040N028N029P007(0)='1' AND  B( 7)='0' AND B( 6)='1' )then
          cVar2S18S81N025P027nsss(0) <='1';
          else
          cVar2S18S81N025P027nsss(0) <='0';
          end if;
        if(cVar1S19S81N040N028N029P007(0)='1' AND  B( 7)='0' AND B( 6)='0' AND B( 8)='1' )then
          cVar2S19S81N025N027P023nsss(0) <='1';
          else
          cVar2S19S81N025N027P023nsss(0) <='0';
          end if;
        if(cVar1S20S81N040N028N029N007(0)='1' AND  E( 2)='1' AND B(16)='0' AND B( 6)='0' )then
          cVar2S20S81P062P026P027nsss(0) <='1';
          else
          cVar2S20S81P062P026P027nsss(0) <='0';
          end if;
        if(cVar1S21S81N040N028N029N007(0)='1' AND  E( 2)='1' AND B(16)='1' AND D( 0)='1' )then
          cVar2S21S81P062P026P068nsss(0) <='1';
          else
          cVar2S21S81P062P026P068nsss(0) <='0';
          end if;
        if(cVar1S22S81N040N028N029N007(0)='1' AND  E( 2)='0' AND A( 2)='1' AND E( 9)='1' )then
          cVar2S22S81N062P015P067nsss(0) <='1';
          else
          cVar2S22S81N062P015P067nsss(0) <='0';
          end if;
        if(cVar1S0S82P062P007P025P009(0)='1' AND  E( 1)='0' )then
          cVar2S0S82P066nsss(0) <='1';
          else
          cVar2S0S82P066nsss(0) <='0';
          end if;
        if(cVar1S1S82P062P007P025P009(0)='1' AND  D( 5)='1' )then
          cVar2S1S82P048nsss(0) <='1';
          else
          cVar2S1S82P048nsss(0) <='0';
          end if;
        if(cVar1S2S82P062P007N025P003(0)='1' AND  A(10)='0' AND A(12)='0' )then
          cVar2S2S82P018P014nsss(0) <='1';
          else
          cVar2S2S82P018P014nsss(0) <='0';
          end if;
        if(cVar1S3S82P062P007N025P003(0)='1' AND  A(10)='1' AND A(12)='1' )then
          cVar2S3S82P018P014nsss(0) <='1';
          else
          cVar2S3S82P018P014nsss(0) <='0';
          end if;
        if(cVar1S4S82P062P007N025N003(0)='1' AND  D(13)='1' AND B(16)='1' )then
          cVar2S4S82P049P026nsss(0) <='1';
          else
          cVar2S4S82P049P026nsss(0) <='0';
          end if;
        if(cVar1S5S82P062P007N025N003(0)='1' AND  D(13)='1' AND B(16)='0' AND A( 0)='0' )then
          cVar2S5S82P049N026P019nsss(0) <='1';
          else
          cVar2S5S82P049N026P019nsss(0) <='0';
          end if;
        if(cVar1S6S82P062P007N025N003(0)='1' AND  D(13)='0' AND B( 8)='1' AND A( 2)='0' )then
          cVar2S6S82N049P023P015nsss(0) <='1';
          else
          cVar2S6S82N049P023P015nsss(0) <='0';
          end if;
        if(cVar1S7S82P062P007N025N003(0)='1' AND  D(13)='0' AND B( 8)='0' AND A(13)='1' )then
          cVar2S7S82N049N023P012nsss(0) <='1';
          else
          cVar2S7S82N049N023P012nsss(0) <='0';
          end if;
        if(cVar1S8S82P062N007P015P032(0)='1' AND  B( 9)='1' AND A(18)='1' )then
          cVar2S8S82P021P002nsss(0) <='1';
          else
          cVar2S8S82P021P002nsss(0) <='0';
          end if;
        if(cVar1S9S82P062N007P015P032(0)='1' AND  B( 9)='1' AND A(18)='0' AND A( 8)='1' )then
          cVar2S9S82P021N002P003nsss(0) <='1';
          else
          cVar2S9S82P021N002P003nsss(0) <='0';
          end if;
        if(cVar1S10S82P062N007P015P032(0)='1' AND  B( 9)='0' AND D( 1)='0' )then
          cVar2S10S82N021P064nsss(0) <='1';
          else
          cVar2S10S82N021P064nsss(0) <='0';
          end if;
        if(cVar1S11S82P062N007P015P032(0)='1' AND  A(13)='1' AND E(11)='1' AND B(14)='0' )then
          cVar2S11S82P012P059P030nsss(0) <='1';
          else
          cVar2S11S82P012P059P030nsss(0) <='0';
          end if;
        if(cVar1S12S82P062N007P015P032(0)='1' AND  A(13)='1' AND E(11)='0' AND D( 2)='1' )then
          cVar2S12S82P012N059P060nsss(0) <='1';
          else
          cVar2S12S82P012N059P060nsss(0) <='0';
          end if;
        if(cVar1S13S82P062N007P015P032(0)='1' AND  A(13)='0' AND A(12)='1' )then
          cVar2S13S82N012P014nsss(0) <='1';
          else
          cVar2S13S82N012P014nsss(0) <='0';
          end if;
        if(cVar1S14S82P062N007P015P032(0)='1' AND  A(13)='0' AND A(12)='0' AND A( 3)='1' )then
          cVar2S14S82N012N014P013nsss(0) <='1';
          else
          cVar2S14S82N012N014P013nsss(0) <='0';
          end if;
        if(cVar1S15S82P062N007P015P029(0)='1' AND  B(11)='0' )then
          cVar2S15S82P036nsss(0) <='1';
          else
          cVar2S15S82P036nsss(0) <='0';
          end if;
        if(cVar1S16S82P062N007P015N029(0)='1' AND  E( 3)='1' AND B( 2)='0' )then
          cVar2S16S82P058P035nsss(0) <='1';
          else
          cVar2S16S82P058P035nsss(0) <='0';
          end if;
        if(cVar1S17S82P062N007P015N029(0)='1' AND  E( 3)='1' AND B( 2)='1' AND A( 1)='0' )then
          cVar2S17S82P058P035P017nsss(0) <='1';
          else
          cVar2S17S82P058P035P017nsss(0) <='0';
          end if;
        if(cVar1S18S82P062N007P015N029(0)='1' AND  E( 3)='0' AND E(11)='1' AND A(14)='0' )then
          cVar2S18S82N058P059P010nsss(0) <='1';
          else
          cVar2S18S82N058P059P010nsss(0) <='0';
          end if;
        if(cVar1S19S82P062P026P029P050(0)='1' AND  A(10)='1' )then
          cVar2S19S82P018nsss(0) <='1';
          else
          cVar2S19S82P018nsss(0) <='0';
          end if;
        if(cVar1S20S82P062P026P029P050(0)='1' AND  A(10)='0' AND A(12)='0' )then
          cVar2S20S82N018P014nsss(0) <='1';
          else
          cVar2S20S82N018P014nsss(0) <='0';
          end if;
        if(cVar1S21S82P062P026P029N050(0)='1' AND  E(12)='0' AND B( 6)='0' AND D( 9)='0' )then
          cVar2S21S82P055P027P065nsss(0) <='1';
          else
          cVar2S21S82P055P027P065nsss(0) <='0';
          end if;
        if(cVar1S22S82P062P026P029N050(0)='1' AND  E(12)='1' AND D( 0)='1' )then
          cVar2S22S82P055P068nsss(0) <='1';
          else
          cVar2S22S82P055P068nsss(0) <='0';
          end if;
        if(cVar1S23S82P062P026P029P036(0)='1' AND  A( 2)='0' AND A( 4)='1' )then
          cVar2S23S82P015P011nsss(0) <='1';
          else
          cVar2S23S82P015P011nsss(0) <='0';
          end if;
        if(cVar1S1S83P007P025N046P009(0)='1' AND  E(15)='1' )then
          cVar2S1S83P043nsss(0) <='1';
          else
          cVar2S1S83P043nsss(0) <='0';
          end if;
        if(cVar1S2S83P007P025N046P009(0)='1' AND  E(15)='0' AND E( 7)='1' )then
          cVar2S2S83N043P042nsss(0) <='1';
          else
          cVar2S2S83N043P042nsss(0) <='0';
          end if;
        if(cVar1S3S83P007P025N046P009(0)='1' AND  E(15)='0' AND E( 7)='0' AND D(13)='1' )then
          cVar2S3S83N043N042P049nsss(0) <='1';
          else
          cVar2S3S83N043N042P049nsss(0) <='0';
          end if;
        if(cVar1S4S83P007N025P034P063(0)='1' AND  E( 1)='0' AND B( 6)='1' AND A( 4)='0' )then
          cVar2S4S83P066P027P011nsss(0) <='1';
          else
          cVar2S4S83P066P027P011nsss(0) <='0';
          end if;
        if(cVar1S5S83P007N025P034P063(0)='1' AND  E( 1)='0' AND B( 6)='0' )then
          cVar2S5S83P066N027psss(0) <='1';
          else
          cVar2S5S83P066N027psss(0) <='0';
          end if;
        if(cVar1S6S83P007N025P034P063(0)='1' AND  E( 1)='1' AND A( 0)='1' AND A(12)='1' )then
          cVar2S6S83P066P019P014nsss(0) <='1';
          else
          cVar2S6S83P066P019P014nsss(0) <='0';
          end if;
        if(cVar1S7S83P007N025P034P063(0)='1' AND  E( 1)='1' )then
          cVar2S7S83P066nsss(0) <='1';
          else
          cVar2S7S83P066nsss(0) <='0';
          end if;
        if(cVar1S8S83P007N025P034P063(0)='1' AND  E( 1)='0' AND B( 2)='1' )then
          cVar2S8S83N066P035nsss(0) <='1';
          else
          cVar2S8S83N066P035nsss(0) <='0';
          end if;
        if(cVar1S9S83P007N025P034P019(0)='1' AND  E( 2)='0' AND A( 3)='0' )then
          cVar2S9S83P062P013nsss(0) <='1';
          else
          cVar2S9S83P062P013nsss(0) <='0';
          end if;
        if(cVar1S10S83P007N025P034N019(0)='1' AND  A( 5)='1' )then
          cVar2S10S83P009nsss(0) <='1';
          else
          cVar2S10S83P009nsss(0) <='0';
          end if;
        if(cVar1S13S83N007P040N002N047(0)='1' AND  B( 0)='1' )then
          cVar2S13S83P039nsss(0) <='1';
          else
          cVar2S13S83P039nsss(0) <='0';
          end if;
        if(cVar1S14S83N007P040N002N047(0)='1' AND  B( 0)='0' AND A(17)='1' )then
          cVar2S14S83N039P004nsss(0) <='1';
          else
          cVar2S14S83N039P004nsss(0) <='0';
          end if;
        if(cVar1S15S83N007P040N002N047(0)='1' AND  B( 0)='0' AND A(17)='0' AND A(19)='1' )then
          cVar2S15S83N039N004P000nsss(0) <='1';
          else
          cVar2S15S83N039N004P000nsss(0) <='0';
          end if;
        if(cVar1S16S83N007N040P015P038(0)='1' AND  E( 2)='0' AND B( 5)='1' AND B( 2)='0' )then
          cVar2S16S83P062P029P035nsss(0) <='1';
          else
          cVar2S16S83P062P029P035nsss(0) <='0';
          end if;
        if(cVar1S17S83N007N040P015P038(0)='1' AND  E( 2)='0' AND B( 5)='0' AND A(16)='0' )then
          cVar2S17S83P062N029P006nsss(0) <='1';
          else
          cVar2S17S83P062N029P006nsss(0) <='0';
          end if;
        if(cVar1S18S83N007N040N015P034(0)='1' AND  A(12)='1' AND B( 3)='0' )then
          cVar2S18S83P014P033nsss(0) <='1';
          else
          cVar2S18S83P014P033nsss(0) <='0';
          end if;
        if(cVar1S19S83N007N040N015P034(0)='1' AND  A(12)='0' AND D( 1)='0' AND E(11)='0' )then
          cVar2S19S83N014P064P059nsss(0) <='1';
          else
          cVar2S19S83N014P064P059nsss(0) <='0';
          end if;
        if(cVar1S20S83N007N040N015N034(0)='1' AND  A( 9)='0' AND A( 8)='0' AND E( 5)='1' )then
          cVar2S20S83P001P003P050nsss(0) <='1';
          else
          cVar2S20S83P001P003P050nsss(0) <='0';
          end if;
        if(cVar1S21S83N007N040N015N034(0)='1' AND  A( 9)='0' AND A( 8)='1' AND B( 0)='1' )then
          cVar2S21S83P001P003P039nsss(0) <='1';
          else
          cVar2S21S83P001P003P039nsss(0) <='0';
          end if;
        if(cVar1S22S83N007N040N015N034(0)='1' AND  A( 9)='1' AND B( 0)='1' )then
          cVar2S22S83P001P039nsss(0) <='1';
          else
          cVar2S22S83P001P039nsss(0) <='0';
          end if;
        if(cVar1S23S83N007N040N015N034(0)='1' AND  A( 9)='1' AND B( 0)='0' AND A(14)='1' )then
          cVar2S23S83P001N039P010nsss(0) <='1';
          else
          cVar2S23S83P001N039P010nsss(0) <='0';
          end if;
        if(cVar1S1S84P040P021N002P012(0)='1' AND  A( 8)='1' )then
          cVar2S1S84P003nsss(0) <='1';
          else
          cVar2S1S84P003nsss(0) <='0';
          end if;
        if(cVar1S2S84P040P021N002P012(0)='1' AND  A( 8)='0' AND A(17)='1' )then
          cVar2S2S84N003P004nsss(0) <='1';
          else
          cVar2S2S84N003P004nsss(0) <='0';
          end if;
        if(cVar1S3S84P040P021N002P012(0)='1' AND  A( 8)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S3S84N003N004P005nsss(0) <='1';
          else
          cVar2S3S84N003N004P005nsss(0) <='0';
          end if;
        if(cVar1S5S84P040N021N057P008(0)='1' AND  B( 0)='1' )then
          cVar2S5S84P039nsss(0) <='1';
          else
          cVar2S5S84P039nsss(0) <='0';
          end if;
        if(cVar1S6S84P040N021N057P008(0)='1' AND  B( 0)='0' AND D( 2)='1' )then
          cVar2S6S84N039P060nsss(0) <='1';
          else
          cVar2S6S84N039P060nsss(0) <='0';
          end if;
        if(cVar1S7S84P040N021N057P008(0)='1' AND  B( 0)='0' AND D( 2)='0' AND A( 5)='0' )then
          cVar2S7S84N039N060P009nsss(0) <='1';
          else
          cVar2S7S84N039N060P009nsss(0) <='0';
          end if;
        if(cVar1S8S84N040P007P025P046(0)='1' AND  A( 4)='0' )then
          cVar2S8S84P011nsss(0) <='1';
          else
          cVar2S8S84P011nsss(0) <='0';
          end if;
        if(cVar1S9S84N040P007P025N046(0)='1' AND  E(14)='1' )then
          cVar2S9S84P047nsss(0) <='1';
          else
          cVar2S9S84P047nsss(0) <='0';
          end if;
        if(cVar1S10S84N040P007P025N046(0)='1' AND  E(14)='0' AND E( 7)='1' )then
          cVar2S10S84N047P042nsss(0) <='1';
          else
          cVar2S10S84N047P042nsss(0) <='0';
          end if;
        if(cVar1S11S84N040P007P025N046(0)='1' AND  E(14)='0' AND E( 7)='0' AND E(15)='1' )then
          cVar2S11S84N047N042P043nsss(0) <='1';
          else
          cVar2S11S84N047N042P043nsss(0) <='0';
          end if;
        if(cVar1S12S84N040P007N025P055(0)='1' AND  A( 4)='0' )then
          cVar2S12S84P011nsss(0) <='1';
          else
          cVar2S12S84P011nsss(0) <='0';
          end if;
        if(cVar1S13S84N040P007N025P055(0)='1' AND  A( 4)='1' AND A( 2)='1' AND A(13)='0' )then
          cVar2S13S84P011P015P012nsss(0) <='1';
          else
          cVar2S13S84P011P015P012nsss(0) <='0';
          end if;
        if(cVar1S14S84N040P007N025P055(0)='1' AND  A( 4)='1' AND A( 2)='0' AND A(13)='1' )then
          cVar2S14S84P011N015P012nsss(0) <='1';
          else
          cVar2S14S84P011N015P012nsss(0) <='0';
          end if;
        if(cVar1S15S84N040P007N025P055(0)='1' AND  A(14)='1' )then
          cVar2S15S84P010nsss(0) <='1';
          else
          cVar2S15S84P010nsss(0) <='0';
          end if;
        if(cVar1S16S84N040N007P015P001(0)='1' AND  A( 8)='0' AND B(19)='0' AND B( 0)='0' )then
          cVar2S16S84P003P020P039nsss(0) <='1';
          else
          cVar2S16S84P003P020P039nsss(0) <='0';
          end if;
        if(cVar1S17S84N040N007P015P001(0)='1' AND  A( 8)='0' AND B(19)='1' AND A(18)='1' )then
          cVar2S17S84P003P020P002nsss(0) <='1';
          else
          cVar2S17S84P003P020P002nsss(0) <='0';
          end if;
        if(cVar1S18S84N040N007P015P001(0)='1' AND  A( 8)='1' AND B(19)='1' )then
          cVar2S18S84P003P020nsss(0) <='1';
          else
          cVar2S18S84P003P020nsss(0) <='0';
          end if;
        if(cVar1S19S84N040N007P015P001(0)='1' AND  B( 0)='1' )then
          cVar2S19S84P039nsss(0) <='1';
          else
          cVar2S19S84P039nsss(0) <='0';
          end if;
        if(cVar1S20S84N040N007P015P001(0)='1' AND  B( 0)='0' AND A( 8)='1' )then
          cVar2S20S84N039P003nsss(0) <='1';
          else
          cVar2S20S84N039P003nsss(0) <='0';
          end if;
        if(cVar1S21S84N040N007P015P001(0)='1' AND  B( 0)='0' AND A( 8)='0' AND E( 1)='1' )then
          cVar2S21S84N039N003P066nsss(0) <='1';
          else
          cVar2S21S84N039N003P066nsss(0) <='0';
          end if;
        if(cVar1S22S84N040N007P015P035(0)='1' AND  D( 9)='1' AND E( 3)='0' )then
          cVar2S22S84P065P058nsss(0) <='1';
          else
          cVar2S22S84P065P058nsss(0) <='0';
          end if;
        if(cVar1S23S84N040N007P015P035(0)='1' AND  D( 9)='0' AND A( 1)='0' AND D( 0)='0' )then
          cVar2S23S84N065P017P068nsss(0) <='1';
          else
          cVar2S23S84N065P017P068nsss(0) <='0';
          end if;
        if(cVar1S24S84N040N007P015P035(0)='1' AND  D( 9)='0' AND A( 1)='1' AND A(10)='1' )then
          cVar2S24S84N065P017P018nsss(0) <='1';
          else
          cVar2S24S84N065P017P018nsss(0) <='0';
          end if;
        if(cVar1S25S84N040N007P015N035(0)='1' AND  B( 5)='1' AND E(13)='1' )then
          cVar2S25S84P029P051nsss(0) <='1';
          else
          cVar2S25S84P029P051nsss(0) <='0';
          end if;
        if(cVar1S26S84N040N007P015N035(0)='1' AND  B( 5)='1' AND E(13)='0' AND B(15)='0' )then
          cVar2S26S84P029N051P028nsss(0) <='1';
          else
          cVar2S26S84P029N051P028nsss(0) <='0';
          end if;
        if(cVar1S27S84N040N007P015N035(0)='1' AND  B( 5)='0' AND E( 9)='1' )then
          cVar2S27S84N029P067nsss(0) <='1';
          else
          cVar2S27S84N029P067nsss(0) <='0';
          end if;
        if(cVar1S28S84N040N007P015N035(0)='1' AND  B( 5)='0' AND E( 9)='0' AND B(16)='1' )then
          cVar2S28S84N029N067P026nsss(0) <='1';
          else
          cVar2S28S84N029N067P026nsss(0) <='0';
          end if;
        if(cVar1S1S85P015P032N005P003(0)='1' AND  A( 4)='0' AND A(13)='0' )then
          cVar2S1S85P011P012nsss(0) <='1';
          else
          cVar2S1S85P011P012nsss(0) <='0';
          end if;
        if(cVar1S2S85P015P032N005P003(0)='1' AND  A( 4)='0' AND A(13)='1' AND E( 3)='1' )then
          cVar2S2S85P011P012P058nsss(0) <='1';
          else
          cVar2S2S85P011P012P058nsss(0) <='0';
          end if;
        if(cVar1S3S85P015N032P011P008(0)='1' AND  B( 9)='0' )then
          cVar2S3S85P021nsss(0) <='1';
          else
          cVar2S3S85P021nsss(0) <='0';
          end if;
        if(cVar1S4S85P015N032P011P008(0)='1' AND  A(10)='1' AND A( 0)='1' )then
          cVar2S4S85P018P019nsss(0) <='1';
          else
          cVar2S4S85P018P019nsss(0) <='0';
          end if;
        if(cVar1S5S85P015N032N011P000(0)='1' AND  A(14)='1' )then
          cVar2S5S85P010nsss(0) <='1';
          else
          cVar2S5S85P010nsss(0) <='0';
          end if;
        if(cVar1S6S85P015N032N011P000(0)='1' AND  A(14)='0' AND B( 1)='1' )then
          cVar2S6S85N010P037nsss(0) <='1';
          else
          cVar2S6S85N010P037nsss(0) <='0';
          end if;
        if(cVar1S7S85P015N032N011P000(0)='1' AND  A(14)='0' AND B( 1)='0' AND A( 0)='0' )then
          cVar2S7S85N010N037P019nsss(0) <='1';
          else
          cVar2S7S85N010N037P019nsss(0) <='0';
          end if;
        if(cVar1S8S85P015N032N011N000(0)='1' AND  B(10)='0' AND E( 4)='1' AND B(11)='0' )then
          cVar2S8S85P038P054P036nsss(0) <='1';
          else
          cVar2S8S85P038P054P036nsss(0) <='0';
          end if;
        if(cVar1S9S85P015N032N011N000(0)='1' AND  B(10)='1' AND A(18)='1' )then
          cVar2S9S85P038P002nsss(0) <='1';
          else
          cVar2S9S85P038P002nsss(0) <='0';
          end if;
        if(cVar1S11S85N015P021N038P014(0)='1' AND  E( 7)='1' )then
          cVar2S11S85P042nsss(0) <='1';
          else
          cVar2S11S85P042nsss(0) <='0';
          end if;
        if(cVar1S12S85N015P021N038P014(0)='1' AND  E( 7)='0' AND B( 1)='1' )then
          cVar2S12S85N042P037nsss(0) <='1';
          else
          cVar2S12S85N042P037nsss(0) <='0';
          end if;
        if(cVar1S13S85N015P021N038P014(0)='1' AND  E( 7)='0' AND B( 1)='0' AND B( 0)='1' )then
          cVar2S13S85N042N037P039nsss(0) <='1';
          else
          cVar2S13S85N042N037P039nsss(0) <='0';
          end if;
        if(cVar1S14S85N015P021N038P014(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S14S85P016P018nsss(0) <='1';
          else
          cVar2S14S85P016P018nsss(0) <='0';
          end if;
        if(cVar1S16S85N015N021P044N004(0)='1' AND  B( 7)='1' AND A( 1)='0' )then
          cVar2S16S85P025P017nsss(0) <='1';
          else
          cVar2S16S85P025P017nsss(0) <='0';
          end if;
        if(cVar1S17S85N015N021P044N004(0)='1' AND  B( 7)='0' AND A( 7)='1' )then
          cVar2S17S85N025P005nsss(0) <='1';
          else
          cVar2S17S85N025P005nsss(0) <='0';
          end if;
        if(cVar1S18S85N015N021P044N004(0)='1' AND  B( 7)='0' AND A( 7)='0' AND E(15)='1' )then
          cVar2S18S85N025N005P043nsss(0) <='1';
          else
          cVar2S18S85N025N005P043nsss(0) <='0';
          end if;
        if(cVar1S19S85N015N021N044P005(0)='1' AND  A( 3)='1' AND D( 3)='1' )then
          cVar2S19S85P013P056nsss(0) <='1';
          else
          cVar2S19S85P013P056nsss(0) <='0';
          end if;
        if(cVar1S20S85N015N021N044P005(0)='1' AND  A( 3)='1' AND D( 3)='0' AND D( 2)='1' )then
          cVar2S20S85P013N056P060nsss(0) <='1';
          else
          cVar2S20S85P013N056P060nsss(0) <='0';
          end if;
        if(cVar1S21S85N015N021N044P005(0)='1' AND  A( 3)='0' AND D(11)='1' AND A( 4)='1' )then
          cVar2S21S85N013P057P011nsss(0) <='1';
          else
          cVar2S21S85N013P057P011nsss(0) <='0';
          end if;
        if(cVar1S22S85N015N021N044P005(0)='1' AND  D(13)='1' )then
          cVar2S22S85P049nsss(0) <='1';
          else
          cVar2S22S85P049nsss(0) <='0';
          end if;
        if(cVar1S23S85N015N021N044P005(0)='1' AND  D(13)='0' AND E(15)='1' AND A( 0)='0' )then
          cVar2S23S85N049P043P019nsss(0) <='1';
          else
          cVar2S23S85N049P043P019nsss(0) <='0';
          end if;
        if(cVar1S2S86P021P038N002N004(0)='1' AND  A( 8)='1' )then
          cVar2S2S86P003nsss(0) <='1';
          else
          cVar2S2S86P003nsss(0) <='0';
          end if;
        if(cVar1S3S86P021P038N002N004(0)='1' AND  A( 8)='0' AND A( 7)='1' )then
          cVar2S3S86N003P005nsss(0) <='1';
          else
          cVar2S3S86N003P005nsss(0) <='0';
          end if;
        if(cVar1S5S86P021N038P010N042(0)='1' AND  A( 4)='0' )then
          cVar2S5S86P011nsss(0) <='1';
          else
          cVar2S5S86P011nsss(0) <='0';
          end if;
        if(cVar1S8S86N021P020P039N003(0)='1' AND  A(18)='1' )then
          cVar2S8S86P002nsss(0) <='1';
          else
          cVar2S8S86P002nsss(0) <='0';
          end if;
        if(cVar1S9S86N021P020P039N003(0)='1' AND  A(18)='0' AND A( 7)='1' )then
          cVar2S9S86N002P005nsss(0) <='1';
          else
          cVar2S9S86N002P005nsss(0) <='0';
          end if;
        if(cVar1S10S86N021P020P039N003(0)='1' AND  A(18)='0' AND A( 7)='0' AND A(17)='1' )then
          cVar2S10S86N002N005P004nsss(0) <='1';
          else
          cVar2S10S86N002N005P004nsss(0) <='0';
          end if;
        if(cVar1S11S86N021P020N039P031(0)='1' AND  A( 3)='1' AND E( 1)='1' )then
          cVar2S11S86P013P066nsss(0) <='1';
          else
          cVar2S11S86P013P066nsss(0) <='0';
          end if;
        if(cVar1S12S86N021P020N039P031(0)='1' AND  A( 3)='1' AND E( 1)='0' AND A(10)='1' )then
          cVar2S12S86P013N066P018nsss(0) <='1';
          else
          cVar2S12S86P013N066P018nsss(0) <='0';
          end if;
        if(cVar1S13S86N021P020N039P031(0)='1' AND  A( 3)='0' AND A( 8)='1' )then
          cVar2S13S86N013P003nsss(0) <='1';
          else
          cVar2S13S86N013P003nsss(0) <='0';
          end if;
        if(cVar1S14S86N021P020N039P031(0)='1' AND  A( 3)='0' AND A( 8)='0' AND D(12)='1' )then
          cVar2S14S86N013N003P053nsss(0) <='1';
          else
          cVar2S14S86N013N003P053nsss(0) <='0';
          end if;
        if(cVar1S15S86N021N020P002P015(0)='1' AND  A(12)='0' AND E(12)='1' AND A( 0)='0' )then
          cVar2S15S86P014P055P019nsss(0) <='1';
          else
          cVar2S15S86P014P055P019nsss(0) <='0';
          end if;
        if(cVar1S16S86N021N020P002P015(0)='1' AND  A(12)='0' AND E(12)='0' AND A( 4)='0' )then
          cVar2S16S86P014N055P011nsss(0) <='1';
          else
          cVar2S16S86P014N055P011nsss(0) <='0';
          end if;
        if(cVar1S17S86N021N020P002P015(0)='1' AND  A(12)='1' AND A( 7)='1' )then
          cVar2S17S86P014P005nsss(0) <='1';
          else
          cVar2S17S86P014P005nsss(0) <='0';
          end if;
        if(cVar1S18S86N021N020P002N015(0)='1' AND  A( 7)='0' )then
          cVar2S18S86P005nsss(0) <='1';
          else
          cVar2S18S86P005nsss(0) <='0';
          end if;
        if(cVar1S19S86N021N020P002N015(0)='1' AND  A( 7)='1' AND D(13)='1' )then
          cVar2S19S86P005P049nsss(0) <='1';
          else
          cVar2S19S86P005P049nsss(0) <='0';
          end if;
        if(cVar1S20S86N021N020P002N015(0)='1' AND  A( 7)='1' AND D(13)='0' AND B( 8)='1' )then
          cVar2S20S86P005N049P023nsss(0) <='1';
          else
          cVar2S20S86P005N049P023nsss(0) <='0';
          end if;
        if(cVar1S21S86N021N020P002P004(0)='1' AND  A( 0)='1' )then
          cVar2S21S86P019nsss(0) <='1';
          else
          cVar2S21S86P019nsss(0) <='0';
          end if;
        if(cVar1S22S86N021N020P002P004(0)='1' AND  A( 0)='0' AND A(14)='1' )then
          cVar2S22S86N019P010nsss(0) <='1';
          else
          cVar2S22S86N019P010nsss(0) <='0';
          end if;
        if(cVar1S23S86N021N020P002N004(0)='1' AND  A(16)='1' AND A( 2)='1' )then
          cVar2S23S86P006P015nsss(0) <='1';
          else
          cVar2S23S86P006P015nsss(0) <='0';
          end if;
        if(cVar1S24S86N021N020P002N004(0)='1' AND  A(16)='0' AND E(12)='0' AND B(17)='1' )then
          cVar2S24S86N006P055P024nsss(0) <='1';
          else
          cVar2S24S86N006P055P024nsss(0) <='0';
          end if;
        if(cVar1S1S87P015P055P061N032(0)='1' AND  E( 9)='1' )then
          cVar2S1S87P067nsss(0) <='1';
          else
          cVar2S1S87P067nsss(0) <='0';
          end if;
        if(cVar1S2S87P015P055P061N032(0)='1' AND  E( 9)='0' AND A( 0)='0' AND D( 3)='0' )then
          cVar2S2S87N067P019P056nsss(0) <='1';
          else
          cVar2S2S87N067P019P056nsss(0) <='0';
          end if;
        if(cVar1S3S87P015P055P061N032(0)='1' AND  E( 9)='0' AND A( 0)='1' AND A(14)='1' )then
          cVar2S3S87N067P019P010nsss(0) <='1';
          else
          cVar2S3S87N067P019P010nsss(0) <='0';
          end if;
        if(cVar1S4S87P015N055P021P020(0)='1' AND  B( 3)='0' AND B( 0)='1' )then
          cVar2S4S87P033P039nsss(0) <='1';
          else
          cVar2S4S87P033P039nsss(0) <='0';
          end if;
        if(cVar1S5S87P015N055P021P020(0)='1' AND  B( 3)='0' AND B( 0)='0' AND A( 0)='0' )then
          cVar2S5S87P033N039P019nsss(0) <='1';
          else
          cVar2S5S87P033N039P019nsss(0) <='0';
          end if;
        if(cVar1S6S87P015N055P021N020(0)='1' AND  B( 0)='0' AND A( 6)='1' AND D( 3)='0' )then
          cVar2S6S87P039P007P056nsss(0) <='1';
          else
          cVar2S6S87P039P007P056nsss(0) <='0';
          end if;
        if(cVar1S7S87P015N055P021N020(0)='1' AND  B( 0)='0' AND A( 6)='0' )then
          cVar2S7S87P039N007psss(0) <='1';
          else
          cVar2S7S87P039N007psss(0) <='0';
          end if;
        if(cVar1S8S87P015N055P021N020(0)='1' AND  B( 0)='1' AND A( 1)='1' )then
          cVar2S8S87P039P017nsss(0) <='1';
          else
          cVar2S8S87P039P017nsss(0) <='0';
          end if;
        if(cVar1S10S87P015N055P021N066(0)='1' AND  A(12)='1' AND A(11)='0' )then
          cVar2S10S87P014P016nsss(0) <='1';
          else
          cVar2S10S87P014P016nsss(0) <='0';
          end if;
        if(cVar1S11S87P015N055P021N066(0)='1' AND  A(12)='0' AND A(10)='1' )then
          cVar2S11S87N014P018nsss(0) <='1';
          else
          cVar2S11S87N014P018nsss(0) <='0';
          end if;
        if(cVar1S13S87N015P021N038P014(0)='1' AND  E( 7)='1' AND A(18)='1' )then
          cVar2S13S87P042P002nsss(0) <='1';
          else
          cVar2S13S87P042P002nsss(0) <='0';
          end if;
        if(cVar1S14S87N015P021N038P014(0)='1' AND  E( 7)='1' AND A(18)='0' AND D(15)='0' )then
          cVar2S14S87P042N002P041nsss(0) <='1';
          else
          cVar2S14S87P042N002P041nsss(0) <='0';
          end if;
        if(cVar1S15S87N015P021N038P014(0)='1' AND  E( 7)='0' AND A( 8)='1' )then
          cVar2S15S87N042P003nsss(0) <='1';
          else
          cVar2S15S87N042P003nsss(0) <='0';
          end if;
        if(cVar1S16S87N015P021N038P014(0)='1' AND  E( 7)='0' AND A( 8)='0' AND A( 5)='0' )then
          cVar2S16S87N042N003P009nsss(0) <='1';
          else
          cVar2S16S87N042N003P009nsss(0) <='0';
          end if;
        if(cVar1S17S87N015P021N038P014(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S17S87P016P018nsss(0) <='1';
          else
          cVar2S17S87P016P018nsss(0) <='0';
          end if;
        if(cVar1S19S87N015N021P020N039(0)='1' AND  B( 2)='0' AND A( 3)='1' )then
          cVar2S19S87P035P013nsss(0) <='1';
          else
          cVar2S19S87P035P013nsss(0) <='0';
          end if;
        if(cVar1S20S87N015N021P020N039(0)='1' AND  B( 2)='0' AND A( 3)='0' AND A( 8)='1' )then
          cVar2S20S87P035N013P003nsss(0) <='1';
          else
          cVar2S20S87P035N013P003nsss(0) <='0';
          end if;
        if(cVar1S21S87N015N021N020P057(0)='1' AND  E(12)='0' AND B(16)='1' AND D(13)='1' )then
          cVar2S21S87P055P026P049nsss(0) <='1';
          else
          cVar2S21S87P055P026P049nsss(0) <='0';
          end if;
        if(cVar1S22S87N015N021N020P057(0)='1' AND  E(12)='1' AND D( 8)='1' )then
          cVar2S22S87P055P069nsss(0) <='1';
          else
          cVar2S22S87P055P069nsss(0) <='0';
          end if;
        if(cVar1S23S87N015N021N020P057(0)='1' AND  E(12)='1' AND D( 8)='0' AND A(14)='1' )then
          cVar2S23S87P055N069P010nsss(0) <='1';
          else
          cVar2S23S87P055N069P010nsss(0) <='0';
          end if;
        if(cVar1S24S87N015N021N020P057(0)='1' AND  B(14)='1' AND A(14)='1' )then
          cVar2S24S87P030P010nsss(0) <='1';
          else
          cVar2S24S87P030P010nsss(0) <='0';
          end if;
        if(cVar1S25S87N015N021N020P057(0)='1' AND  B(14)='1' AND A(14)='0' AND E( 4)='0' )then
          cVar2S25S87P030N010P054nsss(0) <='1';
          else
          cVar2S25S87P030N010P054nsss(0) <='0';
          end if;
        if(cVar1S26S87N015N021N020P057(0)='1' AND  B(14)='0' AND A( 4)='1' AND E(12)='1' )then
          cVar2S26S87N030P011P055nsss(0) <='1';
          else
          cVar2S26S87N030P011P055nsss(0) <='0';
          end if;
        if(cVar1S27S87N015N021N020P057(0)='1' AND  B(14)='0' AND A( 4)='0' AND A( 3)='1' )then
          cVar2S27S87N030N011P013nsss(0) <='1';
          else
          cVar2S27S87N030N011P013nsss(0) <='0';
          end if;
        if(cVar1S0S88P015P057P055P039(0)='1' AND  B(12)='0' AND B(19)='1' )then
          cVar2S0S88P034P020nsss(0) <='1';
          else
          cVar2S0S88P034P020nsss(0) <='0';
          end if;
        if(cVar1S1S88P015P057P055P039(0)='1' AND  B(12)='0' AND B(19)='0' AND A( 1)='0' )then
          cVar2S1S88P034N020P017nsss(0) <='1';
          else
          cVar2S1S88P034N020P017nsss(0) <='0';
          end if;
        if(cVar1S2S88P015P057P055N039(0)='1' AND  B( 2)='0' AND A( 8)='1' AND E( 1)='0' )then
          cVar2S2S88P035P003P066nsss(0) <='1';
          else
          cVar2S2S88P035P003P066nsss(0) <='0';
          end if;
        if(cVar1S3S88P015P057P055N039(0)='1' AND  B( 2)='0' AND A( 8)='0' )then
          cVar2S3S88P035N003psss(0) <='1';
          else
          cVar2S3S88P035N003psss(0) <='0';
          end if;
        if(cVar1S4S88P015P057P055N039(0)='1' AND  B( 2)='1' AND A( 1)='1' )then
          cVar2S4S88P035P017nsss(0) <='1';
          else
          cVar2S4S88P035P017nsss(0) <='0';
          end if;
        if(cVar1S5S88P015P057P055N039(0)='1' AND  B( 2)='1' AND A( 1)='0' AND A(12)='1' )then
          cVar2S5S88P035N017P014nsss(0) <='1';
          else
          cVar2S5S88P035N017P014nsss(0) <='0';
          end if;
        if(cVar1S7S88P015P057P055N069(0)='1' AND  D(12)='1' AND A(14)='1' )then
          cVar2S7S88P053P010nsss(0) <='1';
          else
          cVar2S7S88P053P010nsss(0) <='0';
          end if;
        if(cVar1S8S88P015P057P055N069(0)='1' AND  D(12)='1' AND A(14)='0' AND E(13)='0' )then
          cVar2S8S88P053N010P051nsss(0) <='1';
          else
          cVar2S8S88P053N010P051nsss(0) <='0';
          end if;
        if(cVar1S9S88P015P057P055N069(0)='1' AND  D(12)='0' AND E(10)='1' )then
          cVar2S9S88N053P063nsss(0) <='1';
          else
          cVar2S9S88N053P063nsss(0) <='0';
          end if;
        if(cVar1S10S88P015P057P010P055(0)='1' AND  B(11)='0' AND A(13)='0' )then
          cVar2S10S88P036P012nsss(0) <='1';
          else
          cVar2S10S88P036P012nsss(0) <='0';
          end if;
        if(cVar1S11S88P015P057P010P055(0)='1' AND  B(11)='0' AND A(13)='1' AND B(14)='1' )then
          cVar2S11S88P036P012P030nsss(0) <='1';
          else
          cVar2S11S88P036P012P030nsss(0) <='0';
          end if;
        if(cVar1S12S88P015P057N010P013(0)='1' AND  B( 4)='1' AND A( 1)='0' )then
          cVar2S12S88P031P017nsss(0) <='1';
          else
          cVar2S12S88P031P017nsss(0) <='0';
          end if;
        if(cVar1S13S88P015P057N010P013(0)='1' AND  B( 4)='0' AND B(14)='1' )then
          cVar2S13S88N031P030nsss(0) <='1';
          else
          cVar2S13S88N031P030nsss(0) <='0';
          end if;
        if(cVar1S14S88P015P057N010N013(0)='1' AND  D( 0)='1' AND A( 0)='1' )then
          cVar2S14S88P068P019nsss(0) <='1';
          else
          cVar2S14S88P068P019nsss(0) <='0';
          end if;
        if(cVar1S15S88P015P057N010N013(0)='1' AND  D( 0)='1' AND A( 0)='0' AND B( 1)='0' )then
          cVar2S15S88P068N019P037nsss(0) <='1';
          else
          cVar2S15S88P068N019P037nsss(0) <='0';
          end if;
        if(cVar1S16S88P015P057N010N013(0)='1' AND  D( 0)='0' AND A(13)='1' AND D( 9)='0' )then
          cVar2S16S88N068P012P065nsss(0) <='1';
          else
          cVar2S16S88N068P012P065nsss(0) <='0';
          end if;
        if(cVar1S17S88P015P057N010N013(0)='1' AND  D( 0)='0' AND A(13)='0' AND A( 4)='1' )then
          cVar2S17S88N068N012P011nsss(0) <='1';
          else
          cVar2S17S88N068N012P011nsss(0) <='0';
          end if;
        if(cVar1S19S88P015P055P061N032(0)='1' AND  D(11)='1' )then
          cVar2S19S88P057nsss(0) <='1';
          else
          cVar2S19S88P057nsss(0) <='0';
          end if;
        if(cVar1S20S88P015P055P061N032(0)='1' AND  D(11)='0' AND A( 1)='1' )then
          cVar2S20S88N057P017nsss(0) <='1';
          else
          cVar2S20S88N057P017nsss(0) <='0';
          end if;
        if(cVar1S22S88P015N055P020N002(0)='1' AND  B( 3)='0' AND A( 6)='0' AND A( 0)='0' )then
          cVar2S22S88P033P007P019nsss(0) <='1';
          else
          cVar2S22S88P033P007P019nsss(0) <='0';
          end if;
        if(cVar1S23S88P015N055N020P009(0)='1' AND  B(17)='0' AND A( 7)='1' AND A( 3)='0' )then
          cVar2S23S88P024P005P013nsss(0) <='1';
          else
          cVar2S23S88P024P005P013nsss(0) <='0';
          end if;
        if(cVar1S24S88P015N055N020P009(0)='1' AND  B(17)='0' AND A( 7)='0' )then
          cVar2S24S88P024N005psss(0) <='1';
          else
          cVar2S24S88P024N005psss(0) <='0';
          end if;
        if(cVar1S25S88P015N055N020N009(0)='1' AND  B( 0)='0' AND A( 6)='1' )then
          cVar2S25S88P039P007nsss(0) <='1';
          else
          cVar2S25S88P039P007nsss(0) <='0';
          end if;
        if(cVar1S26S88P015N055N020N009(0)='1' AND  B( 0)='1' AND A( 1)='1' )then
          cVar2S26S88P039P017nsss(0) <='1';
          else
          cVar2S26S88P039P017nsss(0) <='0';
          end if;
        if(cVar1S0S89P015P013P008P059(0)='1' AND  B( 3)='1' )then
          cVar2S0S89P033nsss(0) <='1';
          else
          cVar2S0S89P033nsss(0) <='0';
          end if;
        if(cVar1S1S89P015P013P008P059(0)='1' AND  B( 3)='0' AND B( 1)='0' AND A( 0)='0' )then
          cVar2S1S89N033P037P019nsss(0) <='1';
          else
          cVar2S1S89N033P037P019nsss(0) <='0';
          end if;
        if(cVar1S2S89P015P013P008P059(0)='1' AND  B( 3)='0' AND B( 1)='1' AND A(10)='1' )then
          cVar2S2S89N033P037P018nsss(0) <='1';
          else
          cVar2S2S89N033P037P018nsss(0) <='0';
          end if;
        if(cVar1S3S89P015P013P008N059(0)='1' AND  A(13)='1' AND B( 3)='0' AND E( 6)='0' )then
          cVar2S3S89P012P033P046nsss(0) <='1';
          else
          cVar2S3S89P012P033P046nsss(0) <='0';
          end if;
        if(cVar1S4S89P015P013P008N059(0)='1' AND  A(13)='0' AND B(13)='1' AND B( 3)='0' )then
          cVar2S4S89N012P032P033nsss(0) <='1';
          else
          cVar2S4S89N012P032P033nsss(0) <='0';
          end if;
        if(cVar1S5S89P015P013P008N059(0)='1' AND  A(13)='0' AND B(13)='0' AND B( 2)='1' )then
          cVar2S5S89N012N032P035nsss(0) <='1';
          else
          cVar2S5S89N012N032P035nsss(0) <='0';
          end if;
        if(cVar1S6S89P015P013P008P019(0)='1' AND  E(10)='1' )then
          cVar2S6S89P063nsss(0) <='1';
          else
          cVar2S6S89P063nsss(0) <='0';
          end if;
        if(cVar1S7S89P015P013P008P019(0)='1' AND  E(10)='0' AND B( 2)='0' AND A(12)='1' )then
          cVar2S7S89N063P035P014nsss(0) <='1';
          else
          cVar2S7S89N063P035P014nsss(0) <='0';
          end if;
        if(cVar1S8S89P015P013P008N019(0)='1' AND  D( 4)='1' )then
          cVar2S8S89P052nsss(0) <='1';
          else
          cVar2S8S89P052nsss(0) <='0';
          end if;
        if(cVar1S9S89P015P013P059P055(0)='1' AND  D(11)='1' )then
          cVar2S9S89P057nsss(0) <='1';
          else
          cVar2S9S89P057nsss(0) <='0';
          end if;
        if(cVar1S10S89P015P013P059N055(0)='1' AND  A( 7)='1' AND A( 0)='0' )then
          cVar2S10S89P005P019nsss(0) <='1';
          else
          cVar2S10S89P005P019nsss(0) <='0';
          end if;
        if(cVar1S11S89P015P013P059N055(0)='1' AND  A( 7)='1' AND A( 0)='1' AND A(12)='0' )then
          cVar2S11S89P005P019P014nsss(0) <='1';
          else
          cVar2S11S89P005P019P014nsss(0) <='0';
          end if;
        if(cVar1S12S89P015P013P059N055(0)='1' AND  A( 7)='0' AND A( 0)='1' AND A(10)='0' )then
          cVar2S12S89N005P019P018nsss(0) <='1';
          else
          cVar2S12S89N005P019P018nsss(0) <='0';
          end if;
        if(cVar1S13S89P015P013P059N055(0)='1' AND  A( 7)='0' AND A( 0)='0' AND D( 0)='1' )then
          cVar2S13S89N005N019P068nsss(0) <='1';
          else
          cVar2S13S89N005N019P068nsss(0) <='0';
          end if;
        if(cVar1S14S89P015P013P059P061(0)='1' AND  E( 3)='1' )then
          cVar2S14S89P058nsss(0) <='1';
          else
          cVar2S14S89P058nsss(0) <='0';
          end if;
        if(cVar1S15S89P015P013P059P061(0)='1' AND  E( 3)='0' AND B(13)='1' )then
          cVar2S15S89N058P032nsss(0) <='1';
          else
          cVar2S15S89N058P032nsss(0) <='0';
          end if;
        if(cVar1S17S89N015P039P020N003(0)='1' AND  A(18)='1' )then
          cVar2S17S89P002nsss(0) <='1';
          else
          cVar2S17S89P002nsss(0) <='0';
          end if;
        if(cVar1S18S89N015P039P020N003(0)='1' AND  A(18)='0' AND A( 7)='1' )then
          cVar2S18S89N002P005nsss(0) <='1';
          else
          cVar2S18S89N002P005nsss(0) <='0';
          end if;
        if(cVar1S19S89N015P039N020P017(0)='1' AND  B( 9)='1' )then
          cVar2S19S89P021nsss(0) <='1';
          else
          cVar2S19S89P021nsss(0) <='0';
          end if;
        if(cVar1S20S89N015P039N020P017(0)='1' AND  B( 9)='0' AND A( 4)='0' )then
          cVar2S20S89N021P011nsss(0) <='1';
          else
          cVar2S20S89N021P011nsss(0) <='0';
          end if;
        if(cVar1S21S89N015N039P044P025(0)='1' AND  A( 1)='0' AND A(12)='0' )then
          cVar2S21S89P017P014nsss(0) <='1';
          else
          cVar2S21S89P017P014nsss(0) <='0';
          end if;
        if(cVar1S22S89N015N039P044N025(0)='1' AND  A( 7)='1' AND B( 8)='1' )then
          cVar2S22S89P005P023nsss(0) <='1';
          else
          cVar2S22S89P005P023nsss(0) <='0';
          end if;
        if(cVar1S23S89N015N039P044N025(0)='1' AND  A( 7)='0' AND A(17)='1' AND E( 7)='1' )then
          cVar2S23S89N005P004P042nsss(0) <='1';
          else
          cVar2S23S89N005P004P042nsss(0) <='0';
          end if;
        if(cVar1S24S89N015N039P044N025(0)='1' AND  A( 7)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S24S89N005N004P006nsss(0) <='1';
          else
          cVar2S24S89N005N004P006nsss(0) <='0';
          end if;
        if(cVar1S25S89N015N039N044P038(0)='1' AND  B( 9)='1' )then
          cVar2S25S89P021nsss(0) <='1';
          else
          cVar2S25S89P021nsss(0) <='0';
          end if;
        if(cVar1S26S89N015N039N044P038(0)='1' AND  B( 9)='0' AND A( 1)='0' AND A(13)='1' )then
          cVar2S26S89N021P017P012nsss(0) <='1';
          else
          cVar2S26S89N021P017P012nsss(0) <='0';
          end if;
        if(cVar1S27S89N015N039N044N038(0)='1' AND  B( 6)='1' AND A( 5)='1' )then
          cVar2S27S89P027P009nsss(0) <='1';
          else
          cVar2S27S89P027P009nsss(0) <='0';
          end if;
        if(cVar1S28S89N015N039N044N038(0)='1' AND  B( 6)='1' AND A( 5)='0' AND B( 1)='0' )then
          cVar2S28S89P027N009P037nsss(0) <='1';
          else
          cVar2S28S89P027N009P037nsss(0) <='0';
          end if;
        if(cVar1S29S89N015N039N044N038(0)='1' AND  B( 6)='0' AND E( 7)='1' AND D( 1)='1' )then
          cVar2S29S89N027P042P064nsss(0) <='1';
          else
          cVar2S29S89N027P042P064nsss(0) <='0';
          end if;
        if(cVar1S1S90P020P039P010N003(0)='1' AND  D(15)='1' )then
          cVar2S1S90P041nsss(0) <='1';
          else
          cVar2S1S90P041nsss(0) <='0';
          end if;
        if(cVar1S3S90P020N039N025P031(0)='1' AND  E( 5)='0' AND B(17)='1' )then
          cVar2S3S90P050P024nsss(0) <='1';
          else
          cVar2S3S90P050P024nsss(0) <='0';
          end if;
        if(cVar1S4S90P020N039N025P031(0)='1' AND  E( 5)='0' AND B(17)='0' AND E(13)='0' )then
          cVar2S4S90P050N024P051nsss(0) <='1';
          else
          cVar2S4S90P050N024P051nsss(0) <='0';
          end if;
        if(cVar1S6S90N020P040P021N002(0)='1' AND  A(10)='1' )then
          cVar2S6S90P018nsss(0) <='1';
          else
          cVar2S6S90P018nsss(0) <='0';
          end if;
        if(cVar1S7S90N020P040P021N002(0)='1' AND  A(10)='0' AND A(17)='1' )then
          cVar2S7S90N018P004nsss(0) <='1';
          else
          cVar2S7S90N018P004nsss(0) <='0';
          end if;
        if(cVar1S8S90N020P040P021N002(0)='1' AND  A(10)='0' AND A(17)='0' AND A( 8)='1' )then
          cVar2S8S90N018N004P003nsss(0) <='1';
          else
          cVar2S8S90N018N004P003nsss(0) <='0';
          end if;
        if(cVar1S10S90N020P040N021N057(0)='1' AND  A( 8)='0' AND A( 5)='0' AND E( 7)='0' )then
          cVar2S10S90P003P009P042nsss(0) <='1';
          else
          cVar2S10S90P003P009P042nsss(0) <='0';
          end if;
        if(cVar1S11S90N020N040P039P045(0)='1' AND  E(15)='1' AND D( 9)='0' )then
          cVar2S11S90P043P065nsss(0) <='1';
          else
          cVar2S11S90P043P065nsss(0) <='0';
          end if;
        if(cVar1S12S90N020N040P039P045(0)='1' AND  E(15)='0' AND D( 5)='1' )then
          cVar2S12S90N043P048nsss(0) <='1';
          else
          cVar2S12S90N043P048nsss(0) <='0';
          end if;
        if(cVar1S13S90N020N040P039P045(0)='1' AND  E(15)='0' AND D( 5)='0' AND D( 2)='1' )then
          cVar2S13S90N043N048P060nsss(0) <='1';
          else
          cVar2S13S90N043N048P060nsss(0) <='0';
          end if;
        if(cVar1S14S90N020N040P039N045(0)='1' AND  A( 2)='1' AND A( 3)='0' AND B( 7)='0' )then
          cVar2S14S90P015P013P025nsss(0) <='1';
          else
          cVar2S14S90P015P013P025nsss(0) <='0';
          end if;
        if(cVar1S15S90N020N040P039N045(0)='1' AND  A( 2)='1' AND A( 3)='1' AND E(11)='0' )then
          cVar2S15S90P015P013P059nsss(0) <='1';
          else
          cVar2S15S90P015P013P059nsss(0) <='0';
          end if;
        if(cVar1S16S90N020N040P039N045(0)='1' AND  A( 2)='0' AND D(11)='0' AND E(12)='0' )then
          cVar2S16S90N015P057P055nsss(0) <='1';
          else
          cVar2S16S90N015P057P055nsss(0) <='0';
          end if;
        if(cVar1S17S90N020N040P039N045(0)='1' AND  A( 2)='0' AND D(11)='1' AND A(14)='1' )then
          cVar2S17S90N015P057P010nsss(0) <='1';
          else
          cVar2S17S90N015P057P010nsss(0) <='0';
          end if;
        if(cVar1S1S91P020P039P010N003(0)='1' AND  D(15)='1' )then
          cVar2S1S91P041nsss(0) <='1';
          else
          cVar2S1S91P041nsss(0) <='0';
          end if;
        if(cVar1S4S91P020N039N025N024(0)='1' AND  D(12)='1' )then
          cVar2S4S91P053nsss(0) <='1';
          else
          cVar2S4S91P053nsss(0) <='0';
          end if;
        if(cVar1S5S91P020N039N025N024(0)='1' AND  D(12)='0' AND D( 8)='0' AND B(13)='1' )then
          cVar2S5S91N053P069P032nsss(0) <='1';
          else
          cVar2S5S91N053P069P032nsss(0) <='0';
          end if;
        if(cVar1S7S91N020P045P004P018(0)='1' AND  B(18)='1' )then
          cVar2S7S91P022nsss(0) <='1';
          else
          cVar2S7S91P022nsss(0) <='0';
          end if;
        if(cVar1S8S91N020P045N004P006(0)='1' AND  B(17)='1' )then
          cVar2S8S91P024nsss(0) <='1';
          else
          cVar2S8S91P024nsss(0) <='0';
          end if;
        if(cVar1S9S91N020P045N004P006(0)='1' AND  B(17)='0' AND B(18)='1' )then
          cVar2S9S91N024P022nsss(0) <='1';
          else
          cVar2S9S91N024P022nsss(0) <='0';
          end if;
        if(cVar1S10S91N020P045N004N006(0)='1' AND  A( 6)='1' )then
          cVar2S10S91P007nsss(0) <='1';
          else
          cVar2S10S91P007nsss(0) <='0';
          end if;
        if(cVar1S11S91N020P045N004N006(0)='1' AND  A( 6)='0' AND E(13)='1' )then
          cVar2S11S91N007P051nsss(0) <='1';
          else
          cVar2S11S91N007P051nsss(0) <='0';
          end if;
        if(cVar1S12S91N020P045N004N006(0)='1' AND  A( 6)='0' AND E(13)='0' AND A(12)='1' )then
          cVar2S12S91N007N051P014nsss(0) <='1';
          else
          cVar2S12S91N007N051P014nsss(0) <='0';
          end if;
        if(cVar1S14S91N020N045P040N021(0)='1' AND  E( 4)='1' )then
          cVar2S14S91P054nsss(0) <='1';
          else
          cVar2S14S91P054nsss(0) <='0';
          end if;
        if(cVar1S15S91N020N045P040N021(0)='1' AND  E( 4)='0' AND A( 8)='0' AND A(12)='1' )then
          cVar2S15S91N054P003P014nsss(0) <='1';
          else
          cVar2S15S91N054P003P014nsss(0) <='0';
          end if;
        if(cVar1S16S91N020N045N040P055(0)='1' AND  A(14)='1' AND B(15)='1' AND A(13)='0' )then
          cVar2S16S91P010P028P012nsss(0) <='1';
          else
          cVar2S16S91P010P028P012nsss(0) <='0';
          end if;
        if(cVar1S17S91N020N045N040P055(0)='1' AND  A(14)='1' AND B(15)='0' AND B(14)='1' )then
          cVar2S17S91P010N028P030nsss(0) <='1';
          else
          cVar2S17S91P010N028P030nsss(0) <='0';
          end if;
        if(cVar1S18S91N020N045N040P055(0)='1' AND  A(14)='0' AND E( 9)='1' )then
          cVar2S18S91N010P067nsss(0) <='1';
          else
          cVar2S18S91N010P067nsss(0) <='0';
          end if;
        if(cVar1S19S91N020N045N040N055(0)='1' AND  D(11)='0' AND E(15)='1' AND D( 9)='1' )then
          cVar2S19S91P057P043P065nsss(0) <='1';
          else
          cVar2S19S91P057P043P065nsss(0) <='0';
          end if;
        if(cVar1S20S91N020N045N040N055(0)='1' AND  D(11)='1' AND E(11)='1' )then
          cVar2S20S91P057P059nsss(0) <='1';
          else
          cVar2S20S91P057P059nsss(0) <='0';
          end if;
        if(cVar1S21S91N020N045N040N055(0)='1' AND  D(11)='1' AND E(11)='0' AND D( 0)='1' )then
          cVar2S21S91P057N059P068nsss(0) <='1';
          else
          cVar2S21S91P057N059P068nsss(0) <='0';
          end if;
        if(cVar1S1S92P020P039P010N003(0)='1' AND  A(18)='1' )then
          cVar2S1S92P002nsss(0) <='1';
          else
          cVar2S1S92P002nsss(0) <='0';
          end if;
        if(cVar1S2S92P020P039P010N003(0)='1' AND  A(18)='0' AND A( 0)='0' )then
          cVar2S2S92N002P019nsss(0) <='1';
          else
          cVar2S2S92N002P019nsss(0) <='0';
          end if;
        if(cVar1S4S92P020N039N025P031(0)='1' AND  B( 2)='0' AND B( 5)='0' )then
          cVar2S4S92P035P029nsss(0) <='1';
          else
          cVar2S4S92P035P029nsss(0) <='0';
          end if;
        if(cVar1S5S92P020N039N025P031(0)='1' AND  B( 2)='1' AND A(12)='1' )then
          cVar2S5S92P035P014nsss(0) <='1';
          else
          cVar2S5S92P035P014nsss(0) <='0';
          end if;
        if(cVar1S7S92N020P045P004P018(0)='1' AND  B(18)='1' )then
          cVar2S7S92P022nsss(0) <='1';
          else
          cVar2S7S92P022nsss(0) <='0';
          end if;
        if(cVar1S8S92N020P045N004P006(0)='1' AND  B(17)='1' )then
          cVar2S8S92P024nsss(0) <='1';
          else
          cVar2S8S92P024nsss(0) <='0';
          end if;
        if(cVar1S9S92N020P045N004P006(0)='1' AND  B(17)='0' AND B(18)='1' )then
          cVar2S9S92N024P022nsss(0) <='1';
          else
          cVar2S9S92N024P022nsss(0) <='0';
          end if;
        if(cVar1S10S92N020P045N004N006(0)='1' AND  A( 6)='1' )then
          cVar2S10S92P007nsss(0) <='1';
          else
          cVar2S10S92P007nsss(0) <='0';
          end if;
        if(cVar1S11S92N020P045N004N006(0)='1' AND  A( 6)='0' AND E(13)='1' )then
          cVar2S11S92N007P051nsss(0) <='1';
          else
          cVar2S11S92N007P051nsss(0) <='0';
          end if;
        if(cVar1S12S92N020P045N004N006(0)='1' AND  A( 6)='0' AND E(13)='0' AND A(12)='1' )then
          cVar2S12S92N007N051P014nsss(0) <='1';
          else
          cVar2S12S92N007N051P014nsss(0) <='0';
          end if;
        if(cVar1S14S92N020N045P040N021(0)='1' AND  A( 8)='0' AND D( 4)='1' )then
          cVar2S14S92P003P052nsss(0) <='1';
          else
          cVar2S14S92P003P052nsss(0) <='0';
          end if;
        if(cVar1S15S92N020N045P040N021(0)='1' AND  A( 8)='0' AND D( 4)='0' AND B( 8)='1' )then
          cVar2S15S92P003N052P023nsss(0) <='1';
          else
          cVar2S15S92P003N052P023nsss(0) <='0';
          end if;
        if(cVar1S16S92N020N045N040P044(0)='1' AND  A(16)='1' AND D( 5)='0' )then
          cVar2S16S92P006P048nsss(0) <='1';
          else
          cVar2S16S92P006P048nsss(0) <='0';
          end if;
        if(cVar1S17S92N020N045N040P044(0)='1' AND  A(16)='0' AND A(18)='1' )then
          cVar2S17S92N006P002nsss(0) <='1';
          else
          cVar2S17S92N006P002nsss(0) <='0';
          end if;
        if(cVar1S18S92N020N045N040P044(0)='1' AND  A(16)='0' AND A(18)='0' AND A( 6)='1' )then
          cVar2S18S92N006N002P007nsss(0) <='1';
          else
          cVar2S18S92N006N002P007nsss(0) <='0';
          end if;
        if(cVar1S19S92N020N045N040N044(0)='1' AND  E( 7)='0' AND B( 8)='0' AND A(18)='0' )then
          cVar2S19S92P042P023P002nsss(0) <='1';
          else
          cVar2S19S92P042P023P002nsss(0) <='0';
          end if;
        if(cVar1S20S92N020N045N040N044(0)='1' AND  E( 7)='0' AND B( 8)='1' AND D(15)='1' )then
          cVar2S20S92P042P023P041nsss(0) <='1';
          else
          cVar2S20S92P042P023P041nsss(0) <='0';
          end if;
        if(cVar1S21S92N020N045N040N044(0)='1' AND  E( 7)='1' AND D( 1)='1' )then
          cVar2S21S92P042P064nsss(0) <='1';
          else
          cVar2S21S92P042P064nsss(0) <='0';
          end if;
        if(cVar1S22S92N020N045N040N044(0)='1' AND  E( 7)='1' AND D( 1)='0' AND B( 2)='1' )then
          cVar2S22S92P042N064P035nsss(0) <='1';
          else
          cVar2S22S92P042N064P035nsss(0) <='0';
          end if;
        if(cVar1S2S93P040P002N021N041(0)='1' AND  B(10)='1' )then
          cVar2S2S93P038nsss(0) <='1';
          else
          cVar2S2S93P038nsss(0) <='0';
          end if;
        if(cVar1S4S93P040N002P004N022(0)='1' AND  B( 8)='1' )then
          cVar2S4S93P023nsss(0) <='1';
          else
          cVar2S4S93P023nsss(0) <='0';
          end if;
        if(cVar1S5S93P040N002P004N022(0)='1' AND  B( 8)='0' AND B(10)='1' )then
          cVar2S5S93N023P038nsss(0) <='1';
          else
          cVar2S5S93N023P038nsss(0) <='0';
          end if;
        if(cVar1S7S93P040N002N004N000(0)='1' AND  D(11)='1' )then
          cVar2S7S93P057nsss(0) <='1';
          else
          cVar2S7S93P057nsss(0) <='0';
          end if;
        if(cVar1S8S93P040N002N004N000(0)='1' AND  D(11)='0' AND E( 5)='1' )then
          cVar2S8S93N057P050nsss(0) <='1';
          else
          cVar2S8S93N057P050nsss(0) <='0';
          end if;
        if(cVar1S9S93P040N002N004N000(0)='1' AND  D(11)='0' AND E( 5)='0' AND A( 7)='1' )then
          cVar2S9S93N057N050P005nsss(0) <='1';
          else
          cVar2S9S93N057N050P005nsss(0) <='0';
          end if;
        if(cVar1S11S93N040P045P022N019(0)='1' AND  A(12)='1' )then
          cVar2S11S93P014nsss(0) <='1';
          else
          cVar2S11S93P014nsss(0) <='0';
          end if;
        if(cVar1S12S93N040P045P022N019(0)='1' AND  A(12)='0' AND A( 6)='1' )then
          cVar2S12S93N014P007nsss(0) <='1';
          else
          cVar2S12S93N014P007nsss(0) <='0';
          end if;
        if(cVar1S13S93N040P045P022N019(0)='1' AND  A(12)='0' AND A( 6)='0' AND A(17)='1' )then
          cVar2S13S93N014N007P004nsss(0) <='1';
          else
          cVar2S13S93N014N007P004nsss(0) <='0';
          end if;
        if(cVar1S14S93N040P045N022P023(0)='1' AND  A( 1)='0' )then
          cVar2S14S93P017nsss(0) <='1';
          else
          cVar2S14S93P017nsss(0) <='0';
          end if;
        if(cVar1S15S93N040P045N022N023(0)='1' AND  B( 6)='0' AND A(16)='1' AND B(17)='1' )then
          cVar2S15S93P027P006P024nsss(0) <='1';
          else
          cVar2S15S93P027P006P024nsss(0) <='0';
          end if;
        if(cVar1S16S93N040P045N022N023(0)='1' AND  B( 6)='0' AND A(16)='0' AND A( 8)='0' )then
          cVar2S16S93P027N006P003nsss(0) <='1';
          else
          cVar2S16S93P027N006P003nsss(0) <='0';
          end if;
        if(cVar1S17S93N040N045P020P039(0)='1' AND  A( 8)='1' )then
          cVar2S17S93P003nsss(0) <='1';
          else
          cVar2S17S93P003nsss(0) <='0';
          end if;
        if(cVar1S18S93N040N045P020P039(0)='1' AND  A( 8)='0' AND A(18)='1' )then
          cVar2S18S93N003P002nsss(0) <='1';
          else
          cVar2S18S93N003P002nsss(0) <='0';
          end if;
        if(cVar1S19S93N040N045P020P039(0)='1' AND  A( 8)='0' AND A(18)='0' AND A( 7)='1' )then
          cVar2S19S93N003N002P005nsss(0) <='1';
          else
          cVar2S19S93N003N002P005nsss(0) <='0';
          end if;
        if(cVar1S20S93N040N045P020N039(0)='1' AND  A(17)='0' AND A(14)='1' )then
          cVar2S20S93P004P010nsss(0) <='1';
          else
          cVar2S20S93P004P010nsss(0) <='0';
          end if;
        if(cVar1S21S93N040N045P020N039(0)='1' AND  A(17)='0' AND A(14)='0' AND D( 5)='1' )then
          cVar2S21S93P004N010P048nsss(0) <='1';
          else
          cVar2S21S93P004N010P048nsss(0) <='0';
          end if;
        if(cVar1S22S93N040N045N020P044(0)='1' AND  A(16)='1' AND D( 5)='0' )then
          cVar2S22S93P006P048nsss(0) <='1';
          else
          cVar2S22S93P006P048nsss(0) <='0';
          end if;
        if(cVar1S23S93N040N045N020P044(0)='1' AND  A(16)='0' AND A(17)='1' AND E( 7)='1' )then
          cVar2S23S93N006P004P042nsss(0) <='1';
          else
          cVar2S23S93N006P004P042nsss(0) <='0';
          end if;
        if(cVar1S24S93N040N045N020P044(0)='1' AND  A(16)='0' AND A(17)='0' AND A( 7)='1' )then
          cVar2S24S93N006N004P005nsss(0) <='1';
          else
          cVar2S24S93N006N004P005nsss(0) <='0';
          end if;
        if(cVar1S25S93N040N045N020N044(0)='1' AND  E( 7)='0' AND A(17)='0' AND B(15)='1' )then
          cVar2S25S93P042P004P028nsss(0) <='1';
          else
          cVar2S25S93P042P004P028nsss(0) <='0';
          end if;
        if(cVar1S26S93N040N045N020N044(0)='1' AND  E( 7)='0' AND A(17)='1' AND A( 7)='1' )then
          cVar2S26S93P042P004P005nsss(0) <='1';
          else
          cVar2S26S93P042P004P005nsss(0) <='0';
          end if;
        if(cVar1S27S93N040N045N020N044(0)='1' AND  E( 7)='1' AND D( 1)='1' )then
          cVar2S27S93P042P064nsss(0) <='1';
          else
          cVar2S27S93P042P064nsss(0) <='0';
          end if;
        if(cVar1S28S93N040N045N020N044(0)='1' AND  E( 7)='1' AND D( 1)='0' AND B( 2)='1' )then
          cVar2S28S93P042N064P035nsss(0) <='1';
          else
          cVar2S28S93P042N064P035nsss(0) <='0';
          end if;
        if(cVar1S2S94P040P002N021N041(0)='1' AND  B(10)='1' )then
          cVar2S2S94P038nsss(0) <='1';
          else
          cVar2S2S94P038nsss(0) <='0';
          end if;
        if(cVar1S4S94P040N002P004N022(0)='1' AND  B( 8)='1' )then
          cVar2S4S94P023nsss(0) <='1';
          else
          cVar2S4S94P023nsss(0) <='0';
          end if;
        if(cVar1S5S94P040N002P004N022(0)='1' AND  B( 8)='0' AND B(10)='1' )then
          cVar2S5S94N023P038nsss(0) <='1';
          else
          cVar2S5S94N023P038nsss(0) <='0';
          end if;
        if(cVar1S7S94N040P044P006P048(0)='1' AND  E( 7)='1' )then
          cVar2S7S94P042nsss(0) <='1';
          else
          cVar2S7S94P042nsss(0) <='0';
          end if;
        if(cVar1S8S94N040P044P006P048(0)='1' AND  E( 7)='0' AND B( 7)='1' )then
          cVar2S8S94N042P025nsss(0) <='1';
          else
          cVar2S8S94N042P025nsss(0) <='0';
          end if;
        if(cVar1S9S94N040P044N006P023(0)='1' AND  A( 7)='1' )then
          cVar2S9S94P005nsss(0) <='1';
          else
          cVar2S9S94P005nsss(0) <='0';
          end if;
        if(cVar1S10S94N040P044N006P023(0)='1' AND  A( 7)='0' AND A(17)='1' )then
          cVar2S10S94N005P004nsss(0) <='1';
          else
          cVar2S10S94N005P004nsss(0) <='0';
          end if;
        if(cVar1S11S94N040P044N006P023(0)='1' AND  A( 7)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S11S94N005N004P007nsss(0) <='1';
          else
          cVar2S11S94N005N004P007nsss(0) <='0';
          end if;
        if(cVar1S12S94N040P044N006N023(0)='1' AND  E(13)='1' )then
          cVar2S12S94P051nsss(0) <='1';
          else
          cVar2S12S94P051nsss(0) <='0';
          end if;
        if(cVar1S13S94N040P044N006N023(0)='1' AND  E(13)='0' AND A(18)='1' )then
          cVar2S13S94N051P002nsss(0) <='1';
          else
          cVar2S13S94N051P002nsss(0) <='0';
          end if;
        if(cVar1S14S94N040P044N006N023(0)='1' AND  E(13)='0' AND A(18)='0' AND E(15)='1' )then
          cVar2S14S94N051N002P043nsss(0) <='1';
          else
          cVar2S14S94N051N002P043nsss(0) <='0';
          end if;
        if(cVar1S15S94N040N044P042P020(0)='1' AND  B( 0)='1' )then
          cVar2S15S94P039nsss(0) <='1';
          else
          cVar2S15S94P039nsss(0) <='0';
          end if;
        if(cVar1S16S94N040N044P042P020(0)='1' AND  B( 0)='0' AND A(17)='0' )then
          cVar2S16S94N039P004nsss(0) <='1';
          else
          cVar2S16S94N039P004nsss(0) <='0';
          end if;
        if(cVar1S17S94N040N044P042N020(0)='1' AND  D(14)='1' AND A(16)='1' )then
          cVar2S17S94P045P006nsss(0) <='1';
          else
          cVar2S17S94P045P006nsss(0) <='0';
          end if;
        if(cVar1S18S94N040N044P042N020(0)='1' AND  D(14)='1' AND A(16)='0' AND B(18)='1' )then
          cVar2S18S94P045N006P022nsss(0) <='1';
          else
          cVar2S18S94P045N006P022nsss(0) <='0';
          end if;
        if(cVar1S19S94N040N044P042N020(0)='1' AND  D(14)='0' AND A(17)='0' )then
          cVar2S19S94N045P004nsss(0) <='1';
          else
          cVar2S19S94N045P004nsss(0) <='0';
          end if;
        if(cVar1S20S94N040N044P042N020(0)='1' AND  D(14)='0' AND A(17)='1' AND A( 0)='1' )then
          cVar2S20S94N045P004P019nsss(0) <='1';
          else
          cVar2S20S94N045P004P019nsss(0) <='0';
          end if;
        if(cVar1S22S94N040N044P042N058(0)='1' AND  D( 8)='1' )then
          cVar2S22S94P069nsss(0) <='1';
          else
          cVar2S22S94P069nsss(0) <='0';
          end if;
        if(cVar1S23S94N040N044P042N058(0)='1' AND  D( 8)='0' AND E(15)='1' )then
          cVar2S23S94N069P043nsss(0) <='1';
          else
          cVar2S23S94N069P043nsss(0) <='0';
          end if;
        if(cVar1S2S95P044P023N005N004(0)='1' AND  A( 6)='1' )then
          cVar2S2S95P007nsss(0) <='1';
          else
          cVar2S2S95P007nsss(0) <='0';
          end if;
        if(cVar1S3S95P044P023N005N004(0)='1' AND  A( 6)='0' AND A(16)='1' )then
          cVar2S3S95N007P006nsss(0) <='1';
          else
          cVar2S3S95N007P006nsss(0) <='0';
          end if;
        if(cVar1S6S95P044N023N051N057(0)='1' AND  A(16)='1' AND B(18)='1' )then
          cVar2S6S95P006P022nsss(0) <='1';
          else
          cVar2S6S95P006P022nsss(0) <='0';
          end if;
        if(cVar1S7S95P044N023N051N057(0)='1' AND  A(16)='1' AND B(18)='0' AND B(17)='1' )then
          cVar2S7S95P006N022P024nsss(0) <='1';
          else
          cVar2S7S95P006N022P024nsss(0) <='0';
          end if;
        if(cVar1S8S95P044N023N051N057(0)='1' AND  A(16)='0' AND D( 2)='1' )then
          cVar2S8S95N006P060nsss(0) <='1';
          else
          cVar2S8S95N006P060nsss(0) <='0';
          end if;
        if(cVar1S9S95P044N023N051N057(0)='1' AND  A(16)='0' AND D( 2)='0' AND E( 4)='1' )then
          cVar2S9S95N006N060P054nsss(0) <='1';
          else
          cVar2S9S95N006N060P054nsss(0) <='0';
          end if;
        if(cVar1S11S95N044P040N002P004(0)='1' AND  B( 8)='1' )then
          cVar2S11S95P023nsss(0) <='1';
          else
          cVar2S11S95P023nsss(0) <='0';
          end if;
        if(cVar1S12S95N044P040N002P004(0)='1' AND  B( 8)='0' AND B(18)='1' )then
          cVar2S12S95N023P022nsss(0) <='1';
          else
          cVar2S12S95N023P022nsss(0) <='0';
          end if;
        if(cVar1S13S95N044P040N002P004(0)='1' AND  B( 8)='0' AND B(18)='0' AND B(10)='1' )then
          cVar2S13S95N023N022P038nsss(0) <='1';
          else
          cVar2S13S95N023N022P038nsss(0) <='0';
          end if;
        if(cVar1S14S95N044P040N002N004(0)='1' AND  A(19)='1' )then
          cVar2S14S95P000nsss(0) <='1';
          else
          cVar2S14S95P000nsss(0) <='0';
          end if;
        if(cVar1S15S95N044P040N002N004(0)='1' AND  A(19)='0' AND B( 0)='1' )then
          cVar2S15S95N000P039nsss(0) <='1';
          else
          cVar2S15S95N000P039nsss(0) <='0';
          end if;
        if(cVar1S16S95N044P040N002N004(0)='1' AND  A(19)='0' AND B( 0)='0' AND A(13)='0' )then
          cVar2S16S95N000N039P012nsss(0) <='1';
          else
          cVar2S16S95N000N039P012nsss(0) <='0';
          end if;
        if(cVar1S18S95N044N040P045N022(0)='1' AND  B( 8)='1' AND A( 1)='0' )then
          cVar2S18S95P023P017nsss(0) <='1';
          else
          cVar2S18S95P023P017nsss(0) <='0';
          end if;
        if(cVar1S19S95N044N040P045N022(0)='1' AND  B( 8)='0' AND A(16)='1' AND B(17)='1' )then
          cVar2S19S95N023P006P024nsss(0) <='1';
          else
          cVar2S19S95N023P006P024nsss(0) <='0';
          end if;
        if(cVar1S20S95N044N040P045N022(0)='1' AND  B( 8)='0' AND A(16)='0' AND E( 9)='1' )then
          cVar2S20S95N023N006P067nsss(0) <='1';
          else
          cVar2S20S95N023N006P067nsss(0) <='0';
          end if;
        if(cVar1S21S95N044N040N045P020(0)='1' AND  B( 0)='1' AND A( 8)='1' )then
          cVar2S21S95P039P003nsss(0) <='1';
          else
          cVar2S21S95P039P003nsss(0) <='0';
          end if;
        if(cVar1S22S95N044N040N045P020(0)='1' AND  B( 0)='1' AND A( 8)='0' AND A(18)='1' )then
          cVar2S22S95P039N003P002nsss(0) <='1';
          else
          cVar2S22S95P039N003P002nsss(0) <='0';
          end if;
        if(cVar1S23S95N044N040N045P020(0)='1' AND  B( 0)='0' AND D( 5)='1' )then
          cVar2S23S95N039P048nsss(0) <='1';
          else
          cVar2S23S95N039P048nsss(0) <='0';
          end if;
        if(cVar1S24S95N044N040N045P020(0)='1' AND  B( 0)='0' AND D( 5)='0' AND A(17)='0' )then
          cVar2S24S95N039N048P004nsss(0) <='1';
          else
          cVar2S24S95N039N048P004nsss(0) <='0';
          end if;
        if(cVar1S25S95N044N040N045N020(0)='1' AND  E( 7)='0' AND A(11)='1' AND B( 3)='0' )then
          cVar2S25S95P042P016P033nsss(0) <='1';
          else
          cVar2S25S95P042P016P033nsss(0) <='0';
          end if;
        if(cVar1S26S95N044N040N045N020(0)='1' AND  E( 7)='0' AND A(11)='0' AND B( 3)='1' )then
          cVar2S26S95P042N016P033nsss(0) <='1';
          else
          cVar2S26S95P042N016P033nsss(0) <='0';
          end if;
        if(cVar1S27S95N044N040N045N020(0)='1' AND  E( 7)='1' AND D( 1)='1' )then
          cVar2S27S95P042P064nsss(0) <='1';
          else
          cVar2S27S95P042P064nsss(0) <='0';
          end if;
        if(cVar1S28S95N044N040N045N020(0)='1' AND  E( 7)='1' AND D( 1)='0' AND B( 2)='1' )then
          cVar2S28S95P042N064P035nsss(0) <='1';
          else
          cVar2S28S95P042N064P035nsss(0) <='0';
          end if;
        if(cVar1S1S96P044P004N023P022(0)='1' AND  A( 0)='0' )then
          cVar2S1S96P019nsss(0) <='1';
          else
          cVar2S1S96P019nsss(0) <='0';
          end if;
        if(cVar1S3S96P044N004N021P005(0)='1' AND  B( 8)='1' )then
          cVar2S3S96P023nsss(0) <='1';
          else
          cVar2S3S96P023nsss(0) <='0';
          end if;
        if(cVar1S4S96P044N004N021N005(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S4S96P006P024nsss(0) <='1';
          else
          cVar2S4S96P006P024nsss(0) <='0';
          end if;
        if(cVar1S5S96P044N004N021N005(0)='1' AND  A(16)='1' AND B(17)='0' AND B( 7)='1' )then
          cVar2S5S96P006N024P025nsss(0) <='1';
          else
          cVar2S5S96P006N024P025nsss(0) <='0';
          end if;
        if(cVar1S6S96P044N004N021N005(0)='1' AND  A(16)='0' AND A( 6)='1' )then
          cVar2S6S96N006P007nsss(0) <='1';
          else
          cVar2S6S96N006P007nsss(0) <='0';
          end if;
        if(cVar1S7S96P044N004N021N005(0)='1' AND  A(16)='0' AND A( 6)='0' AND E( 5)='1' )then
          cVar2S7S96N006N007P050nsss(0) <='1';
          else
          cVar2S7S96N006N007P050nsss(0) <='0';
          end if;
        if(cVar1S8S96N044P016P012P056(0)='1' AND  B(14)='1' )then
          cVar2S8S96P030nsss(0) <='1';
          else
          cVar2S8S96P030nsss(0) <='0';
          end if;
        if(cVar1S9S96N044P016P012P056(0)='1' AND  B(14)='0' AND D( 9)='0' AND B( 4)='1' )then
          cVar2S9S96N030P065P031nsss(0) <='1';
          else
          cVar2S9S96N030P065P031nsss(0) <='0';
          end if;
        if(cVar1S10S96N044P016P012N056(0)='1' AND  E( 9)='0' AND D( 9)='0' )then
          cVar2S10S96P067P065nsss(0) <='1';
          else
          cVar2S10S96P067P065nsss(0) <='0';
          end if;
        if(cVar1S11S96N044P016P012N056(0)='1' AND  E( 9)='0' AND D( 9)='1' AND A( 5)='1' )then
          cVar2S11S96P067P065P009nsss(0) <='1';
          else
          cVar2S11S96P067P065P009nsss(0) <='0';
          end if;
        if(cVar1S12S96N044P016P012N056(0)='1' AND  E( 9)='1' AND B(12)='1' )then
          cVar2S12S96P067P034nsss(0) <='1';
          else
          cVar2S12S96P067P034nsss(0) <='0';
          end if;
        if(cVar1S13S96N044P016P012N056(0)='1' AND  E( 9)='1' AND B(12)='0' AND E( 2)='1' )then
          cVar2S13S96P067N034P062nsss(0) <='1';
          else
          cVar2S13S96P067N034P062nsss(0) <='0';
          end if;
        if(cVar1S14S96N044P016N012P053(0)='1' AND  B(15)='1' AND A( 2)='0' AND A(10)='0' )then
          cVar2S14S96P028P015P018nsss(0) <='1';
          else
          cVar2S14S96P028P015P018nsss(0) <='0';
          end if;
        if(cVar1S15S96N044P016N012P053(0)='1' AND  B(15)='0' AND E( 1)='0' )then
          cVar2S15S96N028P066nsss(0) <='1';
          else
          cVar2S15S96N028P066nsss(0) <='0';
          end if;
        if(cVar1S16S96N044P016N012N053(0)='1' AND  B(14)='0' )then
          cVar2S16S96P030nsss(0) <='1';
          else
          cVar2S16S96P030nsss(0) <='0';
          end if;
        if(cVar1S17S96N044P016N012N053(0)='1' AND  B(14)='1' AND B( 4)='0' AND A(14)='1' )then
          cVar2S17S96P030P031P010nsss(0) <='1';
          else
          cVar2S17S96P030P031P010nsss(0) <='0';
          end if;
        if(cVar1S18S96N044P016P052P059(0)='1' AND  E(14)='0' AND D(12)='0' AND A( 8)='1' )then
          cVar2S18S96P047P053P003nsss(0) <='1';
          else
          cVar2S18S96P047P053P003nsss(0) <='0';
          end if;
        if(cVar1S19S96N044P016P052P059(0)='1' AND  E(14)='1' AND E( 1)='1' )then
          cVar2S19S96P047P066nsss(0) <='1';
          else
          cVar2S19S96P047P066nsss(0) <='0';
          end if;
        if(cVar1S20S96N044P016P052P059(0)='1' AND  E(14)='1' AND E( 1)='0' AND B(16)='1' )then
          cVar2S20S96P047N066P026nsss(0) <='1';
          else
          cVar2S20S96P047N066P026nsss(0) <='0';
          end if;
        if(cVar1S21S96N044P016P052P059(0)='1' AND  E( 2)='1' AND D( 2)='1' )then
          cVar2S21S96P062P060nsss(0) <='1';
          else
          cVar2S21S96P062P060nsss(0) <='0';
          end if;
        if(cVar1S22S96N044P016P052P059(0)='1' AND  E( 2)='1' AND D( 2)='0' AND B(12)='0' )then
          cVar2S22S96P062N060P034nsss(0) <='1';
          else
          cVar2S22S96P062N060P034nsss(0) <='0';
          end if;
        if(cVar1S23S96N044P016P052P059(0)='1' AND  E( 2)='0' AND E( 3)='1' AND A(10)='1' )then
          cVar2S23S96N062P058P018nsss(0) <='1';
          else
          cVar2S23S96N062P058P018nsss(0) <='0';
          end if;
        if(cVar1S25S96N044P016P052N065(0)='1' AND  A( 6)='0' AND A(14)='1' AND E( 5)='1' )then
          cVar2S25S96P007P010P050nsss(0) <='1';
          else
          cVar2S25S96P007P010P050nsss(0) <='0';
          end if;
        if(cVar1S26S96N044P016P052N065(0)='1' AND  A( 6)='0' AND A(14)='0' AND A(15)='1' )then
          cVar2S26S96P007N010P008nsss(0) <='1';
          else
          cVar2S26S96P007N010P008nsss(0) <='0';
          end if;
        if(cVar1S1S97P044P004N023P016(0)='1' AND  A( 0)='0' )then
          cVar2S1S97P019nsss(0) <='1';
          else
          cVar2S1S97P019nsss(0) <='0';
          end if;
        if(cVar1S3S97P044N004N021P005(0)='1' AND  B( 8)='1' )then
          cVar2S3S97P023nsss(0) <='1';
          else
          cVar2S3S97P023nsss(0) <='0';
          end if;
        if(cVar1S4S97P044N004N021P005(0)='1' AND  B( 8)='0' AND B( 7)='1' )then
          cVar2S4S97N023P025nsss(0) <='1';
          else
          cVar2S4S97N023P025nsss(0) <='0';
          end if;
        if(cVar1S5S97P044N004N021N005(0)='1' AND  D(11)='1' )then
          cVar2S5S97P057nsss(0) <='1';
          else
          cVar2S5S97P057nsss(0) <='0';
          end if;
        if(cVar1S6S97P044N004N021N005(0)='1' AND  D(11)='0' AND A(16)='1' )then
          cVar2S6S97N057P006nsss(0) <='1';
          else
          cVar2S6S97N057P006nsss(0) <='0';
          end if;
        if(cVar1S7S97P044N004N021N005(0)='1' AND  D(11)='0' AND A(16)='0' AND E( 1)='1' )then
          cVar2S7S97N057N006P066nsss(0) <='1';
          else
          cVar2S7S97N057N006P066nsss(0) <='0';
          end if;
        if(cVar1S8S97N044P016P052P059(0)='1' AND  E(14)='0' AND D(12)='0' AND B(15)='0' )then
          cVar2S8S97P047P053P028nsss(0) <='1';
          else
          cVar2S8S97P047P053P028nsss(0) <='0';
          end if;
        if(cVar1S9S97N044P016P052P059(0)='1' AND  E(14)='1' AND E( 1)='1' )then
          cVar2S9S97P047P066nsss(0) <='1';
          else
          cVar2S9S97P047P066nsss(0) <='0';
          end if;
        if(cVar1S10S97N044P016P052P059(0)='1' AND  E(14)='1' AND E( 1)='0' AND B(16)='1' )then
          cVar2S10S97P047N066P026nsss(0) <='1';
          else
          cVar2S10S97P047N066P026nsss(0) <='0';
          end if;
        if(cVar1S11S97N044P016P052P059(0)='1' AND  D( 9)='0' AND E( 3)='0' AND A(12)='1' )then
          cVar2S11S97P065P058P014nsss(0) <='1';
          else
          cVar2S11S97P065P058P014nsss(0) <='0';
          end if;
        if(cVar1S12S97N044P016P052P059(0)='1' AND  D( 9)='0' AND E( 3)='1' AND A(10)='1' )then
          cVar2S12S97P065P058P018nsss(0) <='1';
          else
          cVar2S12S97P065P058P018nsss(0) <='0';
          end if;
        if(cVar1S13S97N044P016P052P059(0)='1' AND  D( 9)='1' AND E(10)='1' AND D( 1)='1' )then
          cVar2S13S97P065P063P064nsss(0) <='1';
          else
          cVar2S13S97P065P063P064nsss(0) <='0';
          end if;
        if(cVar1S15S97N044P016P052N065(0)='1' AND  A( 6)='0' AND A(14)='1' AND E( 5)='1' )then
          cVar2S15S97P007P010P050nsss(0) <='1';
          else
          cVar2S15S97P007P010P050nsss(0) <='0';
          end if;
        if(cVar1S16S97N044N016P012P056(0)='1' AND  B(14)='1' )then
          cVar2S16S97P030nsss(0) <='1';
          else
          cVar2S16S97P030nsss(0) <='0';
          end if;
        if(cVar1S17S97N044N016P012P056(0)='1' AND  B(14)='0' AND D( 9)='0' AND B( 4)='1' )then
          cVar2S17S97N030P065P031nsss(0) <='1';
          else
          cVar2S17S97N030P065P031nsss(0) <='0';
          end if;
        if(cVar1S18S97N044N016P012N056(0)='1' AND  B(13)='1' AND A(12)='0' AND E( 1)='0' )then
          cVar2S18S97P032P014P066nsss(0) <='1';
          else
          cVar2S18S97P032P014P066nsss(0) <='0';
          end if;
        if(cVar1S19S97N044N016P012N056(0)='1' AND  B(13)='1' AND A(12)='1' AND A( 0)='0' )then
          cVar2S19S97P032P014P019nsss(0) <='1';
          else
          cVar2S19S97P032P014P019nsss(0) <='0';
          end if;
        if(cVar1S20S97N044N016P012N056(0)='1' AND  B(13)='0' AND E( 4)='0' AND B(14)='1' )then
          cVar2S20S97N032P054P030nsss(0) <='1';
          else
          cVar2S20S97N032P054P030nsss(0) <='0';
          end if;
        if(cVar1S21S97N044N016N012P053(0)='1' AND  B(15)='1' AND A( 4)='1' )then
          cVar2S21S97P028P011nsss(0) <='1';
          else
          cVar2S21S97P028P011nsss(0) <='0';
          end if;
        if(cVar1S22S97N044N016N012P053(0)='1' AND  B(15)='1' AND A( 4)='0' AND A( 2)='0' )then
          cVar2S22S97P028N011P015nsss(0) <='1';
          else
          cVar2S22S97P028N011P015nsss(0) <='0';
          end if;
        if(cVar1S23S97N044N016N012P053(0)='1' AND  B(15)='0' AND E( 1)='0' )then
          cVar2S23S97N028P066nsss(0) <='1';
          else
          cVar2S23S97N028P066nsss(0) <='0';
          end if;
        if(cVar1S24S97N044N016N012N053(0)='1' AND  B(13)='0' AND D(15)='1' )then
          cVar2S24S97P032P041nsss(0) <='1';
          else
          cVar2S24S97P032P041nsss(0) <='0';
          end if;
        if(cVar1S25S97N044N016N012N053(0)='1' AND  B(13)='0' AND D(15)='0' AND D( 7)='1' )then
          cVar2S25S97P032N041P040nsss(0) <='1';
          else
          cVar2S25S97P032N041P040nsss(0) <='0';
          end if;
        if(cVar1S26S97N044N016N012N053(0)='1' AND  B(13)='1' AND A(12)='1' AND D( 2)='1' )then
          cVar2S26S97P032P014P060nsss(0) <='1';
          else
          cVar2S26S97P032P014P060nsss(0) <='0';
          end if;
        if(cVar1S1S98P016P044P004N023(0)='1' AND  A( 0)='0' )then
          cVar2S1S98P019nsss(0) <='1';
          else
          cVar2S1S98P019nsss(0) <='0';
          end if;
        if(cVar1S3S98P016P044N004N047(0)='1' AND  B( 9)='1' )then
          cVar2S3S98P021nsss(0) <='1';
          else
          cVar2S3S98P021nsss(0) <='0';
          end if;
        if(cVar1S4S98P016P044N004N047(0)='1' AND  B( 9)='0' AND B( 7)='1' )then
          cVar2S4S98N021P025nsss(0) <='1';
          else
          cVar2S4S98N021P025nsss(0) <='0';
          end if;
        if(cVar1S5S98P016P044N004N047(0)='1' AND  B( 9)='0' AND B( 7)='0' AND B( 8)='1' )then
          cVar2S5S98N021N025P023nsss(0) <='1';
          else
          cVar2S5S98N021N025P023nsss(0) <='0';
          end if;
        if(cVar1S6S98P016N044P012P056(0)='1' AND  B(14)='1' )then
          cVar2S6S98P030nsss(0) <='1';
          else
          cVar2S6S98P030nsss(0) <='0';
          end if;
        if(cVar1S7S98P016N044P012P056(0)='1' AND  B(14)='0' AND D( 9)='0' )then
          cVar2S7S98N030P065nsss(0) <='1';
          else
          cVar2S7S98N030P065nsss(0) <='0';
          end if;
        if(cVar1S8S98P016N044P012N056(0)='1' AND  D(15)='0' AND B(13)='1' AND A(12)='0' )then
          cVar2S8S98P041P032P014nsss(0) <='1';
          else
          cVar2S8S98P041P032P014nsss(0) <='0';
          end if;
        if(cVar1S9S98P016N044P012N056(0)='1' AND  D(15)='0' AND B(13)='0' )then
          cVar2S9S98P041N032psss(0) <='1';
          else
          cVar2S9S98P041N032psss(0) <='0';
          end if;
        if(cVar1S10S98P016N044P012N056(0)='1' AND  D(15)='1' AND A(10)='0' AND B(19)='1' )then
          cVar2S10S98P041P018P020nsss(0) <='1';
          else
          cVar2S10S98P041P018P020nsss(0) <='0';
          end if;
        if(cVar1S11S98P016N044N012P032(0)='1' AND  E( 5)='0' )then
          cVar2S11S98P050nsss(0) <='1';
          else
          cVar2S11S98P050nsss(0) <='0';
          end if;
        if(cVar1S12S98P016N044N012P032(0)='1' AND  E( 5)='1' AND A(12)='0' AND D( 4)='1' )then
          cVar2S12S98P050P014P052nsss(0) <='1';
          else
          cVar2S12S98P050P014P052nsss(0) <='0';
          end if;
        if(cVar1S13S98P016N044N012P032(0)='1' AND  E( 5)='1' AND A(12)='1' AND B( 6)='1' )then
          cVar2S13S98P050P014P027nsss(0) <='1';
          else
          cVar2S13S98P050P014P027nsss(0) <='0';
          end if;
        if(cVar1S14S98P016N044N012P032(0)='1' AND  A(12)='1' AND D( 2)='1' )then
          cVar2S14S98P014P060nsss(0) <='1';
          else
          cVar2S14S98P014P060nsss(0) <='0';
          end if;
        if(cVar1S15S98P016N044N012P032(0)='1' AND  A(12)='1' AND D( 2)='0' AND E(11)='1' )then
          cVar2S15S98P014N060P059nsss(0) <='1';
          else
          cVar2S15S98P014N060P059nsss(0) <='0';
          end if;
        if(cVar1S16S98P016N044N012P032(0)='1' AND  A(12)='0' AND E( 3)='0' AND A( 6)='1' )then
          cVar2S16S98N014P058P007nsss(0) <='1';
          else
          cVar2S16S98N014P058P007nsss(0) <='0';
          end if;
        if(cVar1S18S98P016P021P037N053(0)='1' AND  B(19)='0' AND A(18)='0' )then
          cVar2S18S98P020P002nsss(0) <='1';
          else
          cVar2S18S98P020P002nsss(0) <='0';
          end if;
        if(cVar1S19S98P016P021N037P047(0)='1' AND  A(18)='1' AND A( 5)='1' )then
          cVar2S19S98P002P009nsss(0) <='1';
          else
          cVar2S19S98P002P009nsss(0) <='0';
          end if;
        if(cVar1S20S98P016P021N037P047(0)='1' AND  A(18)='1' AND A( 5)='0' AND A(10)='0' )then
          cVar2S20S98P002N009P018nsss(0) <='1';
          else
          cVar2S20S98P002N009P018nsss(0) <='0';
          end if;
        if(cVar1S21S98P016P021N037P047(0)='1' AND  A(18)='0' AND D(14)='1' AND A(16)='0' )then
          cVar2S21S98N002P045P006nsss(0) <='1';
          else
          cVar2S21S98N002P045P006nsss(0) <='0';
          end if;
        if(cVar1S22S98P016P021N037P047(0)='1' AND  A(16)='1' )then
          cVar2S22S98P006nsss(0) <='1';
          else
          cVar2S22S98P006nsss(0) <='0';
          end if;
        if(cVar1S23S98P016P021N037P047(0)='1' AND  A(16)='0' AND A(10)='1' AND D(13)='1' )then
          cVar2S23S98N006P018P049nsss(0) <='1';
          else
          cVar2S23S98N006P018P049nsss(0) <='0';
          end if;
        if(cVar1S24S98P016P021N037P047(0)='1' AND  A(16)='0' AND A(10)='0' AND A( 6)='1' )then
          cVar2S24S98N006N018P007nsss(0) <='1';
          else
          cVar2S24S98N006N018P007nsss(0) <='0';
          end if;
        if(cVar1S26S98P016P021P069N038(0)='1' AND  A( 2)='0' AND A( 0)='1' )then
          cVar2S26S98P015P019nsss(0) <='1';
          else
          cVar2S26S98P015P019nsss(0) <='0';
          end if;
        if(cVar1S27S98P016P021P069N038(0)='1' AND  A( 2)='0' AND A( 0)='0' AND A(10)='1' )then
          cVar2S27S98P015N019P018nsss(0) <='1';
          else
          cVar2S27S98P015N019P018nsss(0) <='0';
          end if;
        if(cVar1S3S99P044N051N057N032(0)='1' AND  A(17)='1' AND B( 8)='1' )then
          cVar2S3S99P004P023nsss(0) <='1';
          else
          cVar2S3S99P004P023nsss(0) <='0';
          end if;
        if(cVar1S4S99P044N051N057N032(0)='1' AND  A(17)='1' AND B( 8)='0' AND B(18)='1' )then
          cVar2S4S99P004N023P022nsss(0) <='1';
          else
          cVar2S4S99P004N023P022nsss(0) <='0';
          end if;
        if(cVar1S5S99P044N051N057N032(0)='1' AND  A(17)='0' AND B( 9)='1' )then
          cVar2S5S99N004P021nsss(0) <='1';
          else
          cVar2S5S99N004P021nsss(0) <='0';
          end if;
        if(cVar1S6S99P044N051N057N032(0)='1' AND  A(17)='0' AND B( 9)='0' AND B(10)='0' )then
          cVar2S6S99N004N021P038nsss(0) <='1';
          else
          cVar2S6S99N004N021P038nsss(0) <='0';
          end if;
        if(cVar1S7S99N044P062P003P039(0)='1' AND  B(19)='1' )then
          cVar2S7S99P020nsss(0) <='1';
          else
          cVar2S7S99P020nsss(0) <='0';
          end if;
        if(cVar1S8S99N044P062P003P039(0)='1' AND  B(19)='0' AND B( 9)='1' )then
          cVar2S8S99N020P021nsss(0) <='1';
          else
          cVar2S8S99N020P021nsss(0) <='0';
          end if;
        if(cVar1S9S99N044P062P003N039(0)='1' AND  E( 1)='0' AND B( 2)='0' AND D( 4)='0' )then
          cVar2S9S99P066P035P052nsss(0) <='1';
          else
          cVar2S9S99P066P035P052nsss(0) <='0';
          end if;
        if(cVar1S10S99N044P062P003N039(0)='1' AND  E( 1)='0' AND B( 2)='1' AND A(11)='1' )then
          cVar2S10S99P066P035P016nsss(0) <='1';
          else
          cVar2S10S99P066P035P016nsss(0) <='0';
          end if;
        if(cVar1S11S99N044P062P003N039(0)='1' AND  E( 1)='1' AND E( 3)='0' AND A( 4)='1' )then
          cVar2S11S99P066P058P011nsss(0) <='1';
          else
          cVar2S11S99P066P058P011nsss(0) <='0';
          end if;
        if(cVar1S12S99N044P062N003P042(0)='1' AND  A(15)='1' AND B(16)='1' )then
          cVar2S12S99P008P026nsss(0) <='1';
          else
          cVar2S12S99P008P026nsss(0) <='0';
          end if;
        if(cVar1S13S99N044P062N003P042(0)='1' AND  A(15)='1' AND B(16)='0' AND B(15)='1' )then
          cVar2S13S99P008N026P028nsss(0) <='1';
          else
          cVar2S13S99P008N026P028nsss(0) <='0';
          end if;
        if(cVar1S14S99N044P062N003P042(0)='1' AND  A(15)='0' AND E(14)='0' AND A( 2)='1' )then
          cVar2S14S99N008P047P015nsss(0) <='1';
          else
          cVar2S14S99N008P047P015nsss(0) <='0';
          end if;
        if(cVar1S15S99N044P062N003P042(0)='1' AND  A(15)='0' AND E(14)='1' AND A(16)='1' )then
          cVar2S15S99N008P047P006nsss(0) <='1';
          else
          cVar2S15S99N008P047P006nsss(0) <='0';
          end if;
        if(cVar1S16S99N044P062N003P042(0)='1' AND  B( 8)='1' )then
          cVar2S16S99P023nsss(0) <='1';
          else
          cVar2S16S99P023nsss(0) <='0';
          end if;
        if(cVar1S17S99N044P062N003P042(0)='1' AND  B( 8)='0' AND B( 0)='1' )then
          cVar2S17S99N023P039nsss(0) <='1';
          else
          cVar2S17S99N023P039nsss(0) <='0';
          end if;
        if(cVar1S18S99N044P062N003P042(0)='1' AND  B( 8)='0' AND B( 0)='0' AND A(18)='1' )then
          cVar2S18S99N023N039P002nsss(0) <='1';
          else
          cVar2S18S99N023N039P002nsss(0) <='0';
          end if;
        if(cVar1S20S99N044P062P063N053(0)='1' AND  D( 3)='0' AND D( 2)='1' )then
          cVar2S20S99P056P060nsss(0) <='1';
          else
          cVar2S20S99P056P060nsss(0) <='0';
          end if;
        if(cVar1S21S99N044P062P063N053(0)='1' AND  D( 3)='0' AND D( 2)='0' AND A( 8)='0' )then
          cVar2S21S99P056N060P003nsss(0) <='1';
          else
          cVar2S21S99P056N060P003nsss(0) <='0';
          end if;
        if(cVar1S22S99N044P062N063P009(0)='1' AND  D( 3)='1' AND B( 4)='1' )then
          cVar2S22S99P056P031nsss(0) <='1';
          else
          cVar2S22S99P056P031nsss(0) <='0';
          end if;
        if(cVar1S23S99N044P062N063P009(0)='1' AND  D( 3)='1' AND B( 4)='0' AND B( 2)='0' )then
          cVar2S23S99P056N031P035nsss(0) <='1';
          else
          cVar2S23S99P056N031P035nsss(0) <='0';
          end if;
        if(cVar1S24S99N044P062N063P009(0)='1' AND  D( 3)='0' AND A( 4)='0' AND B(12)='1' )then
          cVar2S24S99N056P011P034nsss(0) <='1';
          else
          cVar2S24S99N056P011P034nsss(0) <='0';
          end if;
        if(cVar1S25S99N044P062N063P009(0)='1' AND  D( 3)='0' AND A( 4)='1' AND A( 1)='1' )then
          cVar2S25S99N056P011P017nsss(0) <='1';
          else
          cVar2S25S99N056P011P017nsss(0) <='0';
          end if;
        if(cVar1S26S99N044P062N063P009(0)='1' AND  B( 3)='0' AND E( 1)='1' AND B( 1)='1' )then
          cVar2S26S99P033P066P037nsss(0) <='1';
          else
          cVar2S26S99P033P066P037nsss(0) <='0';
          end if;
        if(cVar1S27S99N044P062N063P009(0)='1' AND  B( 3)='0' AND E( 1)='0' AND A( 0)='1' )then
          cVar2S27S99P033N066P019nsss(0) <='1';
          else
          cVar2S27S99P033N066P019nsss(0) <='0';
          end if;
        if(cVar1S2S100P015P044N004N021(0)='1' AND  B( 7)='1' AND A( 1)='0' )then
          cVar2S2S100P025P017nsss(0) <='1';
          else
          cVar2S2S100P025P017nsss(0) <='0';
          end if;
        if(cVar1S3S100P015P044N004N021(0)='1' AND  B( 7)='0' AND A( 7)='1' )then
          cVar2S3S100N025P005nsss(0) <='1';
          else
          cVar2S3S100N025P005nsss(0) <='0';
          end if;
        if(cVar1S4S100P015P044N004N021(0)='1' AND  B( 7)='0' AND A( 7)='0' AND A( 3)='0' )then
          cVar2S4S100N025N005P013nsss(0) <='1';
          else
          cVar2S4S100N025N005P013nsss(0) <='0';
          end if;
        if(cVar1S6S100P015N044P062N045(0)='1' AND  B(12)='0' AND B( 0)='1' )then
          cVar2S6S100P034P039nsss(0) <='1';
          else
          cVar2S6S100P034P039nsss(0) <='0';
          end if;
        if(cVar1S7S100P015N044P062N045(0)='1' AND  B(12)='0' AND B( 0)='0' AND A( 7)='0' )then
          cVar2S7S100P034N039P005nsss(0) <='1';
          else
          cVar2S7S100P034N039P005nsss(0) <='0';
          end if;
        if(cVar1S8S100P015N044P062N045(0)='1' AND  B(12)='1' AND A(12)='1' AND B( 3)='0' )then
          cVar2S8S100P034P014P033nsss(0) <='1';
          else
          cVar2S8S100P034P014P033nsss(0) <='0';
          end if;
        if(cVar1S9S100P015N044P062P017(0)='1' AND  A(13)='0' AND D(10)='1' )then
          cVar2S9S100P012P061nsss(0) <='1';
          else
          cVar2S9S100P012P061nsss(0) <='0';
          end if;
        if(cVar1S10S100P015N044P062P017(0)='1' AND  A(13)='0' AND D(10)='0' AND B(11)='0' )then
          cVar2S10S100P012N061P036nsss(0) <='1';
          else
          cVar2S10S100P012N061P036nsss(0) <='0';
          end if;
        if(cVar1S11S100P015N044P062P017(0)='1' AND  A(13)='1' AND B(11)='1' )then
          cVar2S11S100P012P036nsss(0) <='1';
          else
          cVar2S11S100P012P036nsss(0) <='0';
          end if;
        if(cVar1S12S100P015N044P062P017(0)='1' AND  A(13)='1' AND B(11)='0' AND A( 3)='1' )then
          cVar2S12S100P012N036P013nsss(0) <='1';
          else
          cVar2S12S100P012N036P013nsss(0) <='0';
          end if;
        if(cVar1S13S100P015N044P062N017(0)='1' AND  A(11)='1' AND A(12)='0' AND D( 1)='1' )then
          cVar2S13S100P016P014P064nsss(0) <='1';
          else
          cVar2S13S100P016P014P064nsss(0) <='0';
          end if;
        if(cVar1S14S100P015N044P062N017(0)='1' AND  A(11)='1' AND A(12)='1' AND A(10)='1' )then
          cVar2S14S100P016P014P018nsss(0) <='1';
          else
          cVar2S14S100P016P014P018nsss(0) <='0';
          end if;
        if(cVar1S15S100P015N044P062N017(0)='1' AND  A(11)='0' AND A(12)='1' AND B(12)='1' )then
          cVar2S15S100N016P014P034nsss(0) <='1';
          else
          cVar2S15S100N016P014P034nsss(0) <='0';
          end if;
        if(cVar1S16S100P015N044P062N017(0)='1' AND  A(11)='0' AND A(12)='0' AND A( 0)='1' )then
          cVar2S16S100N016N014P019nsss(0) <='1';
          else
          cVar2S16S100N016N014P019nsss(0) <='0';
          end if;
        if(cVar1S17S100P015P013P056P032(0)='1' AND  A(13)='0' AND D(11)='1' )then
          cVar2S17S100P012P057nsss(0) <='1';
          else
          cVar2S17S100P012P057nsss(0) <='0';
          end if;
        if(cVar1S18S100P015P013P056P032(0)='1' AND  A(13)='0' AND D(11)='0' AND A(10)='0' )then
          cVar2S18S100P012N057P018nsss(0) <='1';
          else
          cVar2S18S100P012N057P018nsss(0) <='0';
          end if;
        if(cVar1S19S100P015P013P056N032(0)='1' AND  D( 0)='0' AND E( 1)='1' AND A(12)='1' )then
          cVar2S19S100P068P066P014nsss(0) <='1';
          else
          cVar2S19S100P068P066P014nsss(0) <='0';
          end if;
        if(cVar1S20S100P015P013P056N032(0)='1' AND  D( 0)='1' AND E( 1)='0' AND E( 2)='0' )then
          cVar2S20S100P068P066P062nsss(0) <='1';
          else
          cVar2S20S100P068P066P062nsss(0) <='0';
          end if;
        if(cVar1S21S100P015P013P056N032(0)='1' AND  D( 0)='1' AND E( 1)='1' AND E( 2)='1' )then
          cVar2S21S100P068P066P062nsss(0) <='1';
          else
          cVar2S21S100P068P066P062nsss(0) <='0';
          end if;
        if(cVar1S22S100P015P013P056P068(0)='1' AND  A(12)='0' )then
          cVar2S22S100P014nsss(0) <='1';
          else
          cVar2S22S100P014nsss(0) <='0';
          end if;
        if(cVar1S23S100P015P013P056N068(0)='1' AND  A( 4)='1' AND A( 0)='0' )then
          cVar2S23S100P011P019nsss(0) <='1';
          else
          cVar2S23S100P011P019nsss(0) <='0';
          end if;
        if(cVar1S25S100P015P013N025P066(0)='1' AND  B( 2)='0' AND B( 1)='1' )then
          cVar2S25S100P035P037nsss(0) <='1';
          else
          cVar2S25S100P035P037nsss(0) <='0';
          end if;
        if(cVar1S26S100P015P013N025P066(0)='1' AND  B( 2)='0' AND B( 1)='0' AND A( 5)='0' )then
          cVar2S26S100P035N037P009nsss(0) <='1';
          else
          cVar2S26S100P035N037P009nsss(0) <='0';
          end if;
        if(cVar1S27S100P015P013N025P066(0)='1' AND  B( 2)='1' AND A( 1)='1' )then
          cVar2S27S100P035P017nsss(0) <='1';
          else
          cVar2S27S100P035P017nsss(0) <='0';
          end if;
        if(cVar1S28S100P015P013N025N066(0)='1' AND  B(17)='1' AND A( 0)='1' )then
          cVar2S28S100P024P019nsss(0) <='1';
          else
          cVar2S28S100P024P019nsss(0) <='0';
          end if;
        if(cVar1S29S100P015P013N025N066(0)='1' AND  B(17)='0' AND B( 4)='1' AND A( 4)='0' )then
          cVar2S29S100N024P031P011nsss(0) <='1';
          else
          cVar2S29S100N024P031P011nsss(0) <='0';
          end if;
        if(cVar1S30S100P015P013N025N066(0)='1' AND  B(17)='0' AND B( 4)='0' AND A(14)='1' )then
          cVar2S30S100N024N031P010nsss(0) <='1';
          else
          cVar2S30S100N024N031P010nsss(0) <='0';
          end if;
        if(cVar1S0S101P015P013P056P068(0)='1' AND  B( 9)='0' AND B(10)='0' )then
          cVar2S0S101P021P038nsss(0) <='1';
          else
          cVar2S0S101P021P038nsss(0) <='0';
          end if;
        if(cVar1S1S101P015P013P056P068(0)='1' AND  B( 9)='1' AND A(12)='1' )then
          cVar2S1S101P021P014nsss(0) <='1';
          else
          cVar2S1S101P021P014nsss(0) <='0';
          end if;
        if(cVar1S2S101P015P013P056P068(0)='1' AND  E( 1)='0' AND E( 9)='1' )then
          cVar2S2S101P066P067nsss(0) <='1';
          else
          cVar2S2S101P066P067nsss(0) <='0';
          end if;
        if(cVar1S3S101P015P013P056P068(0)='1' AND  E( 1)='0' AND E( 9)='0' AND A(13)='0' )then
          cVar2S3S101P066N067P012nsss(0) <='1';
          else
          cVar2S3S101P066N067P012nsss(0) <='0';
          end if;
        if(cVar1S4S101P015P013P056P068(0)='1' AND  E( 1)='1' AND A( 1)='1' AND D( 9)='0' )then
          cVar2S4S101P066P017P065nsss(0) <='1';
          else
          cVar2S4S101P066P017P065nsss(0) <='0';
          end if;
        if(cVar1S5S101P015P013P056P068(0)='1' AND  E( 1)='1' AND A( 1)='0' AND B(11)='1' )then
          cVar2S5S101P066N017P036nsss(0) <='1';
          else
          cVar2S5S101P066N017P036nsss(0) <='0';
          end if;
        if(cVar1S7S101P015P013P056N050(0)='1' AND  A(12)='0' AND B( 5)='1' )then
          cVar2S7S101P014P029nsss(0) <='1';
          else
          cVar2S7S101P014P029nsss(0) <='0';
          end if;
        if(cVar1S8S101P015P013P056N050(0)='1' AND  A(12)='0' AND B( 5)='0' AND A(11)='0' )then
          cVar2S8S101P014N029P016nsss(0) <='1';
          else
          cVar2S8S101P014N029P016nsss(0) <='0';
          end if;
        if(cVar1S10S101P015P013N025P050(0)='1' AND  D( 4)='1' )then
          cVar2S10S101P052nsss(0) <='1';
          else
          cVar2S10S101P052nsss(0) <='0';
          end if;
        if(cVar1S11S101P015P013N025P050(0)='1' AND  D( 4)='0' AND B( 6)='1' )then
          cVar2S11S101N052P027nsss(0) <='1';
          else
          cVar2S11S101N052P027nsss(0) <='0';
          end if;
        if(cVar1S12S101P015P013N025P050(0)='1' AND  D( 4)='0' AND B( 6)='0' AND A(15)='1' )then
          cVar2S12S101N052N027P008nsss(0) <='1';
          else
          cVar2S12S101N052N027P008nsss(0) <='0';
          end if;
        if(cVar1S13S101P015P013N025P050(0)='1' AND  A(13)='1' )then
          cVar2S13S101P012nsss(0) <='1';
          else
          cVar2S13S101P012nsss(0) <='0';
          end if;
        if(cVar1S14S101N015P044P025P017(0)='1' AND  A(12)='0' )then
          cVar2S14S101P014nsss(0) <='1';
          else
          cVar2S14S101P014nsss(0) <='0';
          end if;
        if(cVar1S16S101N015P044N025P005(0)='1' AND  B( 8)='1' )then
          cVar2S16S101P023nsss(0) <='1';
          else
          cVar2S16S101P023nsss(0) <='0';
          end if;
        if(cVar1S17S101N015P044N025N005(0)='1' AND  A(17)='1' AND E( 7)='1' )then
          cVar2S17S101P004P042nsss(0) <='1';
          else
          cVar2S17S101P004P042nsss(0) <='0';
          end if;
        if(cVar1S18S101N015P044N025N005(0)='1' AND  A(17)='0' AND B( 9)='1' )then
          cVar2S18S101N004P021nsss(0) <='1';
          else
          cVar2S18S101N004P021nsss(0) <='0';
          end if;
        if(cVar1S19S101N015P044N025N005(0)='1' AND  A(17)='0' AND B( 9)='0' AND D( 9)='1' )then
          cVar2S19S101N004N021P065nsss(0) <='1';
          else
          cVar2S19S101N004N021P065nsss(0) <='0';
          end if;
        if(cVar1S20S101N015N044P016P052(0)='1' AND  A( 0)='0' AND E(14)='0' AND A( 6)='0' )then
          cVar2S20S101P019P047P007nsss(0) <='1';
          else
          cVar2S20S101P019P047P007nsss(0) <='0';
          end if;
        if(cVar1S21S101N015N044P016P052(0)='1' AND  A( 0)='0' AND E(14)='1' AND A( 6)='1' )then
          cVar2S21S101P019P047P007nsss(0) <='1';
          else
          cVar2S21S101P019P047P007nsss(0) <='0';
          end if;
        if(cVar1S22S101N015N044P016P052(0)='1' AND  A( 0)='1' AND A(14)='0' AND A(17)='1' )then
          cVar2S22S101P019P010P004nsss(0) <='1';
          else
          cVar2S22S101P019P010P004nsss(0) <='0';
          end if;
        if(cVar1S23S101N015N044P016P052(0)='1' AND  A( 0)='1' AND A(14)='1' AND B( 1)='1' )then
          cVar2S23S101P019P010P037nsss(0) <='1';
          else
          cVar2S23S101P019P010P037nsss(0) <='0';
          end if;
        if(cVar1S24S101N015N044P016P052(0)='1' AND  D( 9)='1' )then
          cVar2S24S101P065nsss(0) <='1';
          else
          cVar2S24S101P065nsss(0) <='0';
          end if;
        if(cVar1S25S101N015N044N016P012(0)='1' AND  D( 3)='1' AND B(14)='1' )then
          cVar2S25S101P056P030nsss(0) <='1';
          else
          cVar2S25S101P056P030nsss(0) <='0';
          end if;
        if(cVar1S26S101N015N044N016P012(0)='1' AND  D( 3)='1' AND B(14)='0' AND A( 0)='0' )then
          cVar2S26S101P056N030P019nsss(0) <='1';
          else
          cVar2S26S101P056N030P019nsss(0) <='0';
          end if;
        if(cVar1S27S101N015N044N016P012(0)='1' AND  D( 3)='0' AND B(13)='1' AND B( 2)='0' )then
          cVar2S27S101N056P032P035nsss(0) <='1';
          else
          cVar2S27S101N056P032P035nsss(0) <='0';
          end if;
        if(cVar1S28S101N015N044N016P012(0)='1' AND  D( 3)='0' AND B(13)='0' AND B( 3)='1' )then
          cVar2S28S101N056N032P033nsss(0) <='1';
          else
          cVar2S28S101N056N032P033nsss(0) <='0';
          end if;
        if(cVar1S29S101N015N044N016N012(0)='1' AND  A(18)='1' AND A( 5)='0' )then
          cVar2S29S101P002P009nsss(0) <='1';
          else
          cVar2S29S101P002P009nsss(0) <='0';
          end if;
        if(cVar1S30S101N015N044N016N012(0)='1' AND  A(18)='0' AND B(13)='1' AND A(12)='1' )then
          cVar2S30S101N002P032P014nsss(0) <='1';
          else
          cVar2S30S101N002P032P014nsss(0) <='0';
          end if;
        if(cVar1S1S102P016P015N044P032(0)='1' AND  B( 4)='1' AND D( 3)='1' )then
          cVar2S1S102P031P056nsss(0) <='1';
          else
          cVar2S1S102P031P056nsss(0) <='0';
          end if;
        if(cVar1S2S102P016P015N044P032(0)='1' AND  B( 4)='1' AND D( 3)='0' AND D(10)='1' )then
          cVar2S2S102P031N056P061nsss(0) <='1';
          else
          cVar2S2S102P031N056P061nsss(0) <='0';
          end if;
        if(cVar1S3S102P016P015N044P032(0)='1' AND  B( 4)='0' AND E( 4)='0' )then
          cVar2S3S102N031P054nsss(0) <='1';
          else
          cVar2S3S102N031P054nsss(0) <='0';
          end if;
        if(cVar1S4S102P016P015N044P032(0)='1' AND  B( 4)='0' AND E( 4)='1' AND B( 5)='1' )then
          cVar2S4S102N031P054P029nsss(0) <='1';
          else
          cVar2S4S102N031P054P029nsss(0) <='0';
          end if;
        if(cVar1S5S102P016P015N044P032(0)='1' AND  A(13)='1' AND A(12)='0' AND B( 2)='0' )then
          cVar2S5S102P012P014P035nsss(0) <='1';
          else
          cVar2S5S102P012P014P035nsss(0) <='0';
          end if;
        if(cVar1S6S102P016P015N044P032(0)='1' AND  A(13)='1' AND A(12)='1' AND E(11)='1' )then
          cVar2S6S102P012P014P059nsss(0) <='1';
          else
          cVar2S6S102P012P014P059nsss(0) <='0';
          end if;
        if(cVar1S7S102P016P015N044P032(0)='1' AND  A(13)='0' AND E( 5)='1' )then
          cVar2S7S102N012P050nsss(0) <='1';
          else
          cVar2S7S102N012P050nsss(0) <='0';
          end if;
        if(cVar1S8S102P016P015P043P017(0)='1' AND  B( 2)='1' AND A(18)='0' AND E( 2)='1' )then
          cVar2S8S102P035P002P062nsss(0) <='1';
          else
          cVar2S8S102P035P002P062nsss(0) <='0';
          end if;
        if(cVar1S9S102P016P015P043P017(0)='1' AND  B( 2)='0' AND E(10)='0' AND D( 5)='1' )then
          cVar2S9S102N035P063P048nsss(0) <='1';
          else
          cVar2S9S102N035P063P048nsss(0) <='0';
          end if;
        if(cVar1S10S102P016P015P043P017(0)='1' AND  B( 2)='0' AND E(10)='1' AND B(12)='1' )then
          cVar2S10S102N035P063P034nsss(0) <='1';
          else
          cVar2S10S102N035P063P034nsss(0) <='0';
          end if;
        if(cVar1S11S102P016P015P043P017(0)='1' AND  B(11)='1' AND A( 3)='0' )then
          cVar2S11S102P036P013nsss(0) <='1';
          else
          cVar2S11S102P036P013nsss(0) <='0';
          end if;
        if(cVar1S12S102P016P015P043P017(0)='1' AND  B(11)='1' AND A( 3)='1' AND A(10)='1' )then
          cVar2S12S102P036P013P018nsss(0) <='1';
          else
          cVar2S12S102P036P013P018nsss(0) <='0';
          end if;
        if(cVar1S13S102P016P015P043P017(0)='1' AND  B(11)='0' AND D( 0)='1' AND B( 2)='0' )then
          cVar2S13S102N036P068P035nsss(0) <='1';
          else
          cVar2S13S102N036P068P035nsss(0) <='0';
          end if;
        if(cVar1S14S102P016P015P043P017(0)='1' AND  B(11)='0' AND D( 0)='0' AND B(15)='1' )then
          cVar2S14S102N036N068P028nsss(0) <='1';
          else
          cVar2S14S102N036N068P028nsss(0) <='0';
          end if;
        if(cVar1S16S102P016P015P043N005(0)='1' AND  A(17)='1' )then
          cVar2S16S102P004nsss(0) <='1';
          else
          cVar2S16S102P004nsss(0) <='0';
          end if;
        if(cVar1S17S102P016P021P012P056(0)='1' AND  A( 0)='1' )then
          cVar2S17S102P019nsss(0) <='1';
          else
          cVar2S17S102P019nsss(0) <='0';
          end if;
        if(cVar1S18S102P016P021P012P056(0)='1' AND  A( 0)='0' AND A( 4)='1' AND E( 4)='0' )then
          cVar2S18S102N019P011P054nsss(0) <='1';
          else
          cVar2S18S102N019P011P054nsss(0) <='0';
          end if;
        if(cVar1S19S102P016P021P012P056(0)='1' AND  A( 7)='1' )then
          cVar2S19S102P005nsss(0) <='1';
          else
          cVar2S19S102P005nsss(0) <='0';
          end if;
        if(cVar1S20S102P016P021P012P056(0)='1' AND  A( 7)='0' AND A( 3)='1' AND E( 4)='1' )then
          cVar2S20S102N005P013P054nsss(0) <='1';
          else
          cVar2S20S102N005P013P054nsss(0) <='0';
          end if;
        if(cVar1S22S102P016P021P012N040(0)='1' AND  A(19)='1' AND A(14)='1' )then
          cVar2S22S102P000P010nsss(0) <='1';
          else
          cVar2S22S102P000P010nsss(0) <='0';
          end if;
        if(cVar1S23S102P016P021P012N040(0)='1' AND  A(19)='1' AND A(14)='0' AND A(10)='1' )then
          cVar2S23S102P000N010P018nsss(0) <='1';
          else
          cVar2S23S102P000N010P018nsss(0) <='0';
          end if;
        if(cVar1S24S102P016P021P012N040(0)='1' AND  A(19)='0' AND B(13)='1' AND A( 3)='1' )then
          cVar2S24S102N000P032P013nsss(0) <='1';
          else
          cVar2S24S102N000P032P013nsss(0) <='0';
          end if;
        if(cVar1S26S102P016P021P069N038(0)='1' AND  A(15)='1' )then
          cVar2S26S102P008nsss(0) <='1';
          else
          cVar2S26S102P008nsss(0) <='0';
          end if;
        if(cVar1S27S102P016P021P069N038(0)='1' AND  A(15)='0' AND A( 2)='0' AND A( 0)='1' )then
          cVar2S27S102N008P015P019nsss(0) <='1';
          else
          cVar2S27S102N008P015P019nsss(0) <='0';
          end if;
        if(cVar1S0S103P015P017P063P034(0)='1' AND  B(11)='0' )then
          cVar2S0S103P036nsss(0) <='1';
          else
          cVar2S0S103P036nsss(0) <='0';
          end if;
        if(cVar1S1S103P015P017P063P034(0)='1' AND  B(11)='1' AND A( 4)='1' AND A( 0)='0' )then
          cVar2S1S103P036P011P019nsss(0) <='1';
          else
          cVar2S1S103P036P011P019nsss(0) <='0';
          end if;
        if(cVar1S2S103P015P017P063P034(0)='1' AND  B(11)='1' AND A( 4)='0' AND D( 8)='1' )then
          cVar2S2S103P036N011P069nsss(0) <='1';
          else
          cVar2S2S103P036N011P069nsss(0) <='0';
          end if;
        if(cVar1S3S103P015P017P063P034(0)='1' AND  E(11)='1' AND A(11)='0' )then
          cVar2S3S103P059P016nsss(0) <='1';
          else
          cVar2S3S103P059P016nsss(0) <='0';
          end if;
        if(cVar1S4S103P015P017P063P034(0)='1' AND  E(11)='0' AND A( 0)='1' AND A(11)='0' )then
          cVar2S4S103N059P019P016nsss(0) <='1';
          else
          cVar2S4S103N059P019P016nsss(0) <='0';
          end if;
        if(cVar1S5S103P015P017P063P035(0)='1' AND  D( 9)='1' AND B(12)='0' )then
          cVar2S5S103P065P034nsss(0) <='1';
          else
          cVar2S5S103P065P034nsss(0) <='0';
          end if;
        if(cVar1S6S103P015P017P063N035(0)='1' AND  D( 8)='1' AND A(12)='1' )then
          cVar2S6S103P069P014nsss(0) <='1';
          else
          cVar2S6S103P069P014nsss(0) <='0';
          end if;
        if(cVar1S7S103P015P017P063N035(0)='1' AND  D( 8)='1' AND A(12)='0' AND A(10)='1' )then
          cVar2S7S103P069N014P018nsss(0) <='1';
          else
          cVar2S7S103P069N014P018nsss(0) <='0';
          end if;
        if(cVar1S8S103P015P017P063N035(0)='1' AND  D( 8)='0' AND B(12)='1' AND A(12)='0' )then
          cVar2S8S103N069P034P014nsss(0) <='1';
          else
          cVar2S8S103N069P034P014nsss(0) <='0';
          end if;
        if(cVar1S9S103P015P017P035P014(0)='1' AND  A( 9)='0' AND B( 6)='0' )then
          cVar2S9S103P001P027nsss(0) <='1';
          else
          cVar2S9S103P001P027nsss(0) <='0';
          end if;
        if(cVar1S10S103P015P017P035N014(0)='1' AND  D( 9)='0' AND B(12)='1' )then
          cVar2S10S103P065P034nsss(0) <='1';
          else
          cVar2S10S103P065P034nsss(0) <='0';
          end if;
        if(cVar1S11S103P015P017P035N014(0)='1' AND  D( 9)='0' AND B(12)='0' AND B(17)='1' )then
          cVar2S11S103P065N034P024nsss(0) <='1';
          else
          cVar2S11S103P065N034P024nsss(0) <='0';
          end if;
        if(cVar1S12S103P015P017P035N014(0)='1' AND  D( 9)='1' AND A( 4)='0' AND B(12)='1' )then
          cVar2S12S103P065P011P034nsss(0) <='1';
          else
          cVar2S12S103P065P011P034nsss(0) <='0';
          end if;
        if(cVar1S13S103P015P017P035P065(0)='1' AND  B( 1)='0' )then
          cVar2S13S103P037nsss(0) <='1';
          else
          cVar2S13S103P037nsss(0) <='0';
          end if;
        if(cVar1S15S103N015P044P004N023(0)='1' AND  B(18)='1' )then
          cVar2S15S103P022nsss(0) <='1';
          else
          cVar2S15S103P022nsss(0) <='0';
          end if;
        if(cVar1S16S103N015P044N004P007(0)='1' AND  B( 8)='1' )then
          cVar2S16S103P023nsss(0) <='1';
          else
          cVar2S16S103P023nsss(0) <='0';
          end if;
        if(cVar1S17S103N015P044N004P007(0)='1' AND  B( 8)='0' AND B( 7)='1' )then
          cVar2S17S103N023P025nsss(0) <='1';
          else
          cVar2S17S103N023P025nsss(0) <='0';
          end if;
        if(cVar1S18S103N015P044N004N007(0)='1' AND  E(11)='1' )then
          cVar2S18S103P059nsss(0) <='1';
          else
          cVar2S18S103P059nsss(0) <='0';
          end if;
        if(cVar1S19S103N015P044N004N007(0)='1' AND  E(11)='0' AND A(12)='0' )then
          cVar2S19S103N059P014nsss(0) <='1';
          else
          cVar2S19S103N059P014nsss(0) <='0';
          end if;
        if(cVar1S20S103N015P044N004N007(0)='1' AND  E(11)='0' AND A(12)='1' AND E( 6)='1' )then
          cVar2S20S103N059P014P046nsss(0) <='1';
          else
          cVar2S20S103N059P014P046nsss(0) <='0';
          end if;
        if(cVar1S21S103N015N044P031P013(0)='1' AND  E( 4)='1' )then
          cVar2S21S103P054nsss(0) <='1';
          else
          cVar2S21S103P054nsss(0) <='0';
          end if;
        if(cVar1S22S103N015N044P031P013(0)='1' AND  E( 4)='0' AND A( 4)='0' )then
          cVar2S22S103N054P011nsss(0) <='1';
          else
          cVar2S22S103N054P011nsss(0) <='0';
          end if;
        if(cVar1S23S103N015N044P031N013(0)='1' AND  A( 4)='1' AND D(11)='1' )then
          cVar2S23S103P011P057nsss(0) <='1';
          else
          cVar2S23S103P011P057nsss(0) <='0';
          end if;
        if(cVar1S24S103N015N044P031N013(0)='1' AND  A( 4)='1' AND D(11)='0' AND A( 1)='0' )then
          cVar2S24S103P011N057P017nsss(0) <='1';
          else
          cVar2S24S103P011N057P017nsss(0) <='0';
          end if;
        if(cVar1S25S103N015N044P031N013(0)='1' AND  A( 4)='0' AND E(12)='0' AND A(13)='1' )then
          cVar2S25S103N011P055P012nsss(0) <='1';
          else
          cVar2S25S103N011P055P012nsss(0) <='0';
          end if;
        if(cVar1S26S103N015N044N031P030(0)='1' AND  D( 2)='0' AND A(14)='1' AND B(11)='0' )then
          cVar2S26S103P060P010P036nsss(0) <='1';
          else
          cVar2S26S103P060P010P036nsss(0) <='0';
          end if;
        if(cVar1S27S103N015N044N031P030(0)='1' AND  D( 2)='0' AND A(14)='0' AND A(13)='1' )then
          cVar2S27S103P060N010P012nsss(0) <='1';
          else
          cVar2S27S103P060N010P012nsss(0) <='0';
          end if;
        if(cVar1S28S103N015N044N031P030(0)='1' AND  D( 2)='1' AND E( 1)='1' )then
          cVar2S28S103P060P066nsss(0) <='1';
          else
          cVar2S28S103P060P066nsss(0) <='0';
          end if;
        if(cVar1S29S103N015N044N031P030(0)='1' AND  D( 2)='1' AND E( 1)='0' AND A( 1)='1' )then
          cVar2S29S103P060N066P017nsss(0) <='1';
          else
          cVar2S29S103P060N066P017nsss(0) <='0';
          end if;
        if(cVar1S30S103N015N044N031N030(0)='1' AND  D(11)='0' AND A(14)='1' AND D(12)='1' )then
          cVar2S30S103P057P010P053nsss(0) <='1';
          else
          cVar2S30S103P057P010P053nsss(0) <='0';
          end if;
        if(cVar1S31S103N015N044N031N030(0)='1' AND  D(11)='1' AND D( 2)='1' )then
          cVar2S31S103P057P060nsss(0) <='1';
          else
          cVar2S31S103P057P060nsss(0) <='0';
          end if;
        if(cVar1S32S103N015N044N031N030(0)='1' AND  D(11)='1' AND D( 2)='0' AND E(15)='1' )then
          cVar2S32S103P057N060P043nsss(0) <='1';
          else
          cVar2S32S103P057N060P043nsss(0) <='0';
          end if;
        if(cVar1S0S104P015P005P060P028(0)='1' AND  D( 9)='0' )then
          cVar2S0S104P065nsss(0) <='1';
          else
          cVar2S0S104P065nsss(0) <='0';
          end if;
        if(cVar1S1S104P015P005P060P028(0)='1' AND  D( 9)='1' AND A(10)='1' )then
          cVar2S1S104P065P018nsss(0) <='1';
          else
          cVar2S1S104P065P018nsss(0) <='0';
          end if;
        if(cVar1S2S104P015P005P060P028(0)='1' AND  A(14)='0' )then
          cVar2S2S104P010nsss(0) <='1';
          else
          cVar2S2S104P010nsss(0) <='0';
          end if;
        if(cVar1S4S104P015N005P063P052(0)='1' AND  D( 9)='1' )then
          cVar2S4S104P065nsss(0) <='1';
          else
          cVar2S4S104P065nsss(0) <='0';
          end if;
        if(cVar1S5S104P015N005P063N052(0)='1' AND  B(16)='0' AND B( 2)='1' AND A( 1)='1' )then
          cVar2S5S104P026P035P017nsss(0) <='1';
          else
          cVar2S5S104P026P035P017nsss(0) <='0';
          end if;
        if(cVar1S6S104P015N005P063N052(0)='1' AND  B(16)='0' AND B( 2)='0' AND B( 6)='0' )then
          cVar2S6S104P026N035P027nsss(0) <='1';
          else
          cVar2S6S104P026N035P027nsss(0) <='0';
          end if;
        if(cVar1S7S104P015N005P063N052(0)='1' AND  B(16)='1' AND B(12)='1' )then
          cVar2S7S104P026P034nsss(0) <='1';
          else
          cVar2S7S104P026P034nsss(0) <='0';
          end if;
        if(cVar1S8S104P015N005N063P017(0)='1' AND  A( 3)='1' AND B( 4)='1' )then
          cVar2S8S104P013P031nsss(0) <='1';
          else
          cVar2S8S104P013P031nsss(0) <='0';
          end if;
        if(cVar1S9S104P015N005N063P017(0)='1' AND  A( 3)='1' AND B( 4)='0' AND A(18)='0' )then
          cVar2S9S104P013N031P002nsss(0) <='1';
          else
          cVar2S9S104P013N031P002nsss(0) <='0';
          end if;
        if(cVar1S10S104P015N005N063P017(0)='1' AND  A( 3)='0' AND D(10)='0' AND B(12)='0' )then
          cVar2S10S104N013P061P034nsss(0) <='1';
          else
          cVar2S10S104N013P061P034nsss(0) <='0';
          end if;
        if(cVar1S11S104P015N005N063P017(0)='1' AND  A(15)='1' AND E(14)='1' )then
          cVar2S11S104P008P047nsss(0) <='1';
          else
          cVar2S11S104P008P047nsss(0) <='0';
          end if;
        if(cVar1S12S104P015N005N063P017(0)='1' AND  A(15)='1' AND E(14)='0' AND D( 2)='0' )then
          cVar2S12S104P008N047P060nsss(0) <='1';
          else
          cVar2S12S104P008N047P060nsss(0) <='0';
          end if;
        if(cVar1S13S104P015N005N063P017(0)='1' AND  A(15)='0' AND E(14)='0' AND A( 4)='1' )then
          cVar2S13S104N008P047P011nsss(0) <='1';
          else
          cVar2S13S104N008P047P011nsss(0) <='0';
          end if;
        if(cVar1S14S104P015N005N063P017(0)='1' AND  A(15)='0' AND E(14)='1' AND E( 6)='1' )then
          cVar2S14S104N008P047P046nsss(0) <='1';
          else
          cVar2S14S104N008P047P046nsss(0) <='0';
          end if;
        if(cVar1S15S104P015P029P060P065(0)='1' AND  A( 0)='0' )then
          cVar2S15S104P019nsss(0) <='1';
          else
          cVar2S15S104P019nsss(0) <='0';
          end if;
        if(cVar1S16S104P015P029P060P065(0)='1' AND  A( 0)='1' AND A(13)='1' )then
          cVar2S16S104P019P012nsss(0) <='1';
          else
          cVar2S16S104P019P012nsss(0) <='0';
          end if;
        if(cVar1S17S104P015P029P060P065(0)='1' AND  A( 0)='1' AND A(13)='0' AND A( 4)='1' )then
          cVar2S17S104P019N012P011nsss(0) <='1';
          else
          cVar2S17S104P019N012P011nsss(0) <='0';
          end if;
        if(cVar1S18S104P015N029P056P009(0)='1' AND  E( 4)='1' AND E( 1)='0' )then
          cVar2S18S104P054P066nsss(0) <='1';
          else
          cVar2S18S104P054P066nsss(0) <='0';
          end if;
        if(cVar1S19S104P015N029P056P009(0)='1' AND  E( 4)='0' AND B(16)='0' )then
          cVar2S19S104N054P026nsss(0) <='1';
          else
          cVar2S19S104N054P026nsss(0) <='0';
          end if;
        if(cVar1S20S104P015N029P056P009(0)='1' AND  E( 4)='0' AND B(16)='1' AND D( 4)='1' )then
          cVar2S20S104N054P026P052nsss(0) <='1';
          else
          cVar2S20S104N054P026P052nsss(0) <='0';
          end if;
        if(cVar1S21S104P015N029P056P009(0)='1' AND  E( 4)='0' AND D(13)='1' AND A( 0)='0' )then
          cVar2S21S104P054P049P019nsss(0) <='1';
          else
          cVar2S21S104P054P049P019nsss(0) <='0';
          end if;
        if(cVar1S22S104P015N029P056P009(0)='1' AND  E( 4)='0' AND D(13)='0' AND E( 3)='1' )then
          cVar2S22S104P054N049P058nsss(0) <='1';
          else
          cVar2S22S104P054N049P058nsss(0) <='0';
          end if;
        if(cVar1S23S104P015N029P056P031(0)='1' AND  A(12)='0' )then
          cVar2S23S104P014nsss(0) <='1';
          else
          cVar2S23S104P014nsss(0) <='0';
          end if;
        if(cVar1S24S104P015N029P056N031(0)='1' AND  D( 0)='1' )then
          cVar2S24S104P068nsss(0) <='1';
          else
          cVar2S24S104P068nsss(0) <='0';
          end if;
        if(cVar1S25S104P015N029P056N031(0)='1' AND  D( 0)='0' AND A(13)='1' AND B(14)='1' )then
          cVar2S25S104N068P012P030nsss(0) <='1';
          else
          cVar2S25S104N068P012P030nsss(0) <='0';
          end if;
        if(cVar1S26S104P015N029P056N031(0)='1' AND  D( 0)='0' AND A(13)='0' AND B( 3)='1' )then
          cVar2S26S104N068N012P033nsss(0) <='1';
          else
          cVar2S26S104N068N012P033nsss(0) <='0';
          end if;
        if(cVar1S0S105P017P015P018P013(0)='1' AND  A( 7)='1' AND B( 1)='0' )then
          cVar2S0S105P005P037nsss(0) <='1';
          else
          cVar2S0S105P005P037nsss(0) <='0';
          end if;
        if(cVar1S1S105P017P015P018P013(0)='1' AND  A( 7)='0' )then
          cVar2S1S105N005psss(0) <='1';
          else
          cVar2S1S105N005psss(0) <='0';
          end if;
        if(cVar1S2S105P017P015P018P013(0)='1' AND  A(15)='1' )then
          cVar2S2S105P008nsss(0) <='1';
          else
          cVar2S2S105P008nsss(0) <='0';
          end if;
        if(cVar1S3S105P017P015P018P013(0)='1' AND  A(15)='0' AND A( 4)='1' AND A(14)='0' )then
          cVar2S3S105N008P011P010nsss(0) <='1';
          else
          cVar2S3S105N008P011P010nsss(0) <='0';
          end if;
        if(cVar1S4S105P017P015P018P013(0)='1' AND  A(15)='0' AND A( 4)='0' AND A(14)='1' )then
          cVar2S4S105N008N011P010nsss(0) <='1';
          else
          cVar2S4S105N008N011P010nsss(0) <='0';
          end if;
        if(cVar1S6S105P017P015P018N060(0)='1' AND  D(10)='1' AND B( 2)='1' )then
          cVar2S6S105P061P035nsss(0) <='1';
          else
          cVar2S6S105P061P035nsss(0) <='0';
          end if;
        if(cVar1S7S105P017P015P018N060(0)='1' AND  D(10)='1' AND B( 2)='0' AND E(11)='1' )then
          cVar2S7S105P061N035P059nsss(0) <='1';
          else
          cVar2S7S105P061N035P059nsss(0) <='0';
          end if;
        if(cVar1S8S105P017P015P058P048(0)='1' AND  B( 5)='1' AND E( 5)='1' )then
          cVar2S8S105P029P050nsss(0) <='1';
          else
          cVar2S8S105P029P050nsss(0) <='0';
          end if;
        if(cVar1S9S105P017P015P058P048(0)='1' AND  B( 5)='1' AND E( 5)='0' AND E( 4)='1' )then
          cVar2S9S105P029N050P054nsss(0) <='1';
          else
          cVar2S9S105P029N050P054nsss(0) <='0';
          end if;
        if(cVar1S10S105P017P015P058P048(0)='1' AND  B( 5)='0' AND B(17)='1' AND A( 4)='0' )then
          cVar2S10S105N029P024P011nsss(0) <='1';
          else
          cVar2S10S105N029P024P011nsss(0) <='0';
          end if;
        if(cVar1S11S105P017P015P058P048(0)='1' AND  B( 5)='0' AND B(17)='0' AND B(15)='1' )then
          cVar2S11S105N029N024P028nsss(0) <='1';
          else
          cVar2S11S105N029N024P028nsss(0) <='0';
          end if;
        if(cVar1S12S105P017P015P058P048(0)='1' AND  B( 7)='1' )then
          cVar2S12S105P025nsss(0) <='1';
          else
          cVar2S12S105P025nsss(0) <='0';
          end if;
        if(cVar1S13S105P017P015P058P048(0)='1' AND  B( 7)='0' AND E( 5)='1' )then
          cVar2S13S105N025P050nsss(0) <='1';
          else
          cVar2S13S105N025P050nsss(0) <='0';
          end if;
        if(cVar1S14S105P017P015P058P035(0)='1' AND  A( 3)='1' AND B( 3)='1' )then
          cVar2S14S105P013P033nsss(0) <='1';
          else
          cVar2S14S105P013P033nsss(0) <='0';
          end if;
        if(cVar1S15S105P017P015P058P035(0)='1' AND  A( 3)='0' AND A(13)='0' AND D( 0)='1' )then
          cVar2S15S105N013P012P068nsss(0) <='1';
          else
          cVar2S15S105N013P012P068nsss(0) <='0';
          end if;
        if(cVar1S16S105N017P015P034P014(0)='1' AND  E( 1)='0' AND E(11)='1' )then
          cVar2S16S105P066P059nsss(0) <='1';
          else
          cVar2S16S105P066P059nsss(0) <='0';
          end if;
        if(cVar1S17S105N017P015P034P014(0)='1' AND  E( 1)='0' AND E(11)='0' AND B( 2)='0' )then
          cVar2S17S105P066N059P035nsss(0) <='1';
          else
          cVar2S17S105P066N059P035nsss(0) <='0';
          end if;
        if(cVar1S18S105N017P015P034P014(0)='1' AND  E( 1)='1' AND B( 1)='1' )then
          cVar2S18S105P066P037nsss(0) <='1';
          else
          cVar2S18S105P066P037nsss(0) <='0';
          end if;
        if(cVar1S19S105N017P015P034N014(0)='1' AND  A(11)='1' AND B(11)='0' )then
          cVar2S19S105P016P036nsss(0) <='1';
          else
          cVar2S19S105P016P036nsss(0) <='0';
          end if;
        if(cVar1S20S105N017P015P034N014(0)='1' AND  A(11)='1' AND B(11)='1' AND E( 9)='1' )then
          cVar2S20S105P016P036P067nsss(0) <='1';
          else
          cVar2S20S105P016P036P067nsss(0) <='0';
          end if;
        if(cVar1S21S105N017P015P034N014(0)='1' AND  A(11)='0' AND B( 2)='1' )then
          cVar2S21S105N016P035nsss(0) <='1';
          else
          cVar2S21S105N016P035nsss(0) <='0';
          end if;
        if(cVar1S22S105N017P015P034N014(0)='1' AND  A(11)='0' AND B( 2)='0' AND A( 3)='1' )then
          cVar2S22S105N016N035P013nsss(0) <='1';
          else
          cVar2S22S105N016N035P013nsss(0) <='0';
          end if;
        if(cVar1S23S105N017P015N034P065(0)='1' AND  E( 2)='0' AND B( 0)='1' )then
          cVar2S23S105P062P039nsss(0) <='1';
          else
          cVar2S23S105P062P039nsss(0) <='0';
          end if;
        if(cVar1S24S105N017P015N034P065(0)='1' AND  E( 2)='0' AND B( 0)='0' AND D(10)='1' )then
          cVar2S24S105P062N039P061nsss(0) <='1';
          else
          cVar2S24S105P062N039P061nsss(0) <='0';
          end if;
        if(cVar1S25S105N017P015N034P065(0)='1' AND  E( 2)='1' AND D( 1)='0' AND D( 4)='1' )then
          cVar2S25S105P062N064P052nsss(0) <='1';
          else
          cVar2S25S105P062N064P052nsss(0) <='0';
          end if;
        if(cVar1S26S105N017P015N034P065(0)='1' AND  E( 9)='1' AND E(10)='0' )then
          cVar2S26S105P067P063nsss(0) <='1';
          else
          cVar2S26S105P067P063nsss(0) <='0';
          end if;
        if(cVar1S27S105N017P015N034P065(0)='1' AND  E( 9)='1' AND E(10)='1' AND D( 8)='1' )then
          cVar2S27S105P067P063P069nsss(0) <='1';
          else
          cVar2S27S105P067P063P069nsss(0) <='0';
          end if;
        if(cVar1S28S105N017P015N034P065(0)='1' AND  E( 9)='0' AND B(11)='1' AND A(14)='0' )then
          cVar2S28S105N067P036P010nsss(0) <='1';
          else
          cVar2S28S105N067P036P010nsss(0) <='0';
          end if;
        if(cVar1S30S105N017P015P005N004(0)='1' AND  A(13)='0' AND D( 8)='0' AND A(15)='0' )then
          cVar2S30S105P012P069P008nsss(0) <='1';
          else
          cVar2S30S105P012P069P008nsss(0) <='0';
          end if;
        if(cVar1S31S105N017P015P005N004(0)='1' AND  A(13)='1' AND A(12)='1' )then
          cVar2S31S105P012P014nsss(0) <='1';
          else
          cVar2S31S105P012P014nsss(0) <='0';
          end if;
        if(cVar1S32S105N017P015N005P043(0)='1' AND  A(12)='0' AND D( 5)='1' AND A(13)='0' )then
          cVar2S32S105P014P048P012nsss(0) <='1';
          else
          cVar2S32S105P014P048P012nsss(0) <='0';
          end if;
        if(cVar1S33S105N017P015N005P043(0)='1' AND  A(12)='0' AND D( 5)='0' AND D( 2)='1' )then
          cVar2S33S105P014N048P060nsss(0) <='1';
          else
          cVar2S33S105P014N048P060nsss(0) <='0';
          end if;
        if(cVar1S34S105N017P015N005P043(0)='1' AND  A(12)='1' AND A( 5)='1' AND E( 2)='0' )then
          cVar2S34S105P014P009P062nsss(0) <='1';
          else
          cVar2S34S105P014P009P062nsss(0) <='0';
          end if;
        if(cVar1S35S105N017P015N005P043(0)='1' AND  A(11)='1' )then
          cVar2S35S105P016nsss(0) <='1';
          else
          cVar2S35S105P016nsss(0) <='0';
          end if;
        if(cVar1S36S105N017P015N005P043(0)='1' AND  A(11)='0' AND A(16)='1' )then
          cVar2S36S105N016P006nsss(0) <='1';
          else
          cVar2S36S105N016P006nsss(0) <='0';
          end if;
        if(cVar1S37S105N017P015N005P043(0)='1' AND  A(11)='0' AND A(16)='0' AND A(17)='1' )then
          cVar2S37S105N016N006P004nsss(0) <='1';
          else
          cVar2S37S105N016N006P004nsss(0) <='0';
          end if;
        if(cVar1S0S106P065P015P045P022(0)='1' AND  D( 8)='0' )then
          cVar2S0S106P069nsss(0) <='1';
          else
          cVar2S0S106P069nsss(0) <='0';
          end if;
        if(cVar1S1S106P065P015P045N022(0)='1' AND  E( 2)='0' )then
          cVar2S1S106P062nsss(0) <='1';
          else
          cVar2S1S106P062nsss(0) <='0';
          end if;
        if(cVar1S2S106P065P015N045P043(0)='1' AND  D( 4)='0' )then
          cVar2S2S106P052nsss(0) <='1';
          else
          cVar2S2S106P052nsss(0) <='0';
          end if;
        if(cVar1S3S106P065P015N045P043(0)='1' AND  D( 4)='1' AND A(15)='1' AND B(15)='0' )then
          cVar2S3S106P052P008P028nsss(0) <='1';
          else
          cVar2S3S106P052P008P028nsss(0) <='0';
          end if;
        if(cVar1S4S106P065P015N045P043(0)='1' AND  D( 4)='1' AND A(15)='0' AND A( 5)='1' )then
          cVar2S4S106P052N008P009nsss(0) <='1';
          else
          cVar2S4S106P052N008P009nsss(0) <='0';
          end if;
        if(cVar1S5S106P065P015N045P043(0)='1' AND  B(18)='1' )then
          cVar2S5S106P022nsss(0) <='1';
          else
          cVar2S5S106P022nsss(0) <='0';
          end if;
        if(cVar1S6S106P065P015N045P043(0)='1' AND  B(18)='0' AND D(13)='1' )then
          cVar2S6S106N022P049nsss(0) <='1';
          else
          cVar2S6S106N022P049nsss(0) <='0';
          end if;
        if(cVar1S7S106P065P015N045P043(0)='1' AND  B(18)='0' AND D(13)='0' AND A( 8)='1' )then
          cVar2S7S106N022N049P003nsss(0) <='1';
          else
          cVar2S7S106N022N049P003nsss(0) <='0';
          end if;
        if(cVar1S8S106P065P015P029P060(0)='1' AND  B(11)='0' AND A( 6)='0' )then
          cVar2S8S106P036P007nsss(0) <='1';
          else
          cVar2S8S106P036P007nsss(0) <='0';
          end if;
        if(cVar1S9S106P065P015N029P014(0)='1' AND  E(12)='1' AND A(13)='0' AND A( 0)='0' )then
          cVar2S9S106P055P012P019nsss(0) <='1';
          else
          cVar2S9S106P055P012P019nsss(0) <='0';
          end if;
        if(cVar1S10S106P065P015N029P014(0)='1' AND  E(12)='0' AND B( 9)='0' )then
          cVar2S10S106N055P021nsss(0) <='1';
          else
          cVar2S10S106N055P021nsss(0) <='0';
          end if;
        if(cVar1S11S106P065P015N029P014(0)='1' AND  E(12)='0' AND B( 9)='1' AND A(10)='1' )then
          cVar2S11S106N055P021P018nsss(0) <='1';
          else
          cVar2S11S106N055P021P018nsss(0) <='0';
          end if;
        if(cVar1S12S106P065P015N029P014(0)='1' AND  B( 9)='1' AND A(11)='0' )then
          cVar2S12S106P021P016nsss(0) <='1';
          else
          cVar2S12S106P021P016nsss(0) <='0';
          end if;
        if(cVar1S13S106P065P015N029P014(0)='1' AND  B( 9)='0' AND A(10)='0' AND D( 3)='0' )then
          cVar2S13S106N021P018P056nsss(0) <='1';
          else
          cVar2S13S106N021P018P056nsss(0) <='0';
          end if;
        if(cVar1S14S106P065P015N029P014(0)='1' AND  B( 9)='0' AND A(10)='1' AND B(13)='1' )then
          cVar2S14S106N021P018P032nsss(0) <='1';
          else
          cVar2S14S106N021P018P032nsss(0) <='0';
          end if;
        if(cVar1S16S106P065N052P035P017(0)='1' AND  B( 1)='0' AND B(11)='0' )then
          cVar2S16S106P037P036nsss(0) <='1';
          else
          cVar2S16S106P037P036nsss(0) <='0';
          end if;
        if(cVar1S17S106P065N052P035P017(0)='1' AND  B( 1)='0' AND B(11)='1' AND A(11)='0' )then
          cVar2S17S106P037P036P016nsss(0) <='1';
          else
          cVar2S17S106P037P036P016nsss(0) <='0';
          end if;
        if(cVar1S18S106P065N052P035P017(0)='1' AND  B( 1)='1' AND A( 0)='1' )then
          cVar2S18S106P037P019nsss(0) <='1';
          else
          cVar2S18S106P037P019nsss(0) <='0';
          end if;
        if(cVar1S19S106P065N052P035N017(0)='1' AND  A( 2)='1' AND E( 9)='1' )then
          cVar2S19S106P015P067nsss(0) <='1';
          else
          cVar2S19S106P015P067nsss(0) <='0';
          end if;
        if(cVar1S20S106P065N052P035N017(0)='1' AND  A( 2)='1' AND E( 9)='0' AND B(12)='0' )then
          cVar2S20S106P015N067P034nsss(0) <='1';
          else
          cVar2S20S106P015N067P034nsss(0) <='0';
          end if;
        if(cVar1S21S106P065N052P035N017(0)='1' AND  A( 2)='0' AND E( 2)='0' AND B(12)='1' )then
          cVar2S21S106N015P062P034nsss(0) <='1';
          else
          cVar2S21S106N015P062P034nsss(0) <='0';
          end if;
        if(cVar1S22S106P065N052N035P034(0)='1' AND  E(11)='0' AND B(17)='0' AND D(12)='0' )then
          cVar2S22S106P059P024P053nsss(0) <='1';
          else
          cVar2S22S106P059P024P053nsss(0) <='0';
          end if;
        if(cVar1S23S106P065N052N035P034(0)='1' AND  E(11)='1' AND D( 0)='0' AND A(11)='1' )then
          cVar2S23S106P059P068P016nsss(0) <='1';
          else
          cVar2S23S106P059P068P016nsss(0) <='0';
          end if;
        if(cVar1S24S106P065N052N035N034(0)='1' AND  B(11)='1' AND B( 1)='0' )then
          cVar2S24S106P036P037nsss(0) <='1';
          else
          cVar2S24S106P036P037nsss(0) <='0';
          end if;
        if(cVar1S25S106P065N052N035N034(0)='1' AND  B(11)='0' AND E( 9)='1' AND E(10)='0' )then
          cVar2S25S106N036P067P063nsss(0) <='1';
          else
          cVar2S25S106N036P067P063nsss(0) <='0';
          end if;
        if(cVar1S26S106P065N052N035N034(0)='1' AND  B(11)='0' AND E( 9)='0' AND B( 1)='1' )then
          cVar2S26S106N036N067P037nsss(0) <='1';
          else
          cVar2S26S106N036N067P037nsss(0) <='0';
          end if;
        if(cVar1S1S107P052N065P010P009(0)='1' AND  D( 8)='1' )then
          cVar2S1S107P069nsss(0) <='1';
          else
          cVar2S1S107P069nsss(0) <='0';
          end if;
        if(cVar1S2S107P052N065P010P009(0)='1' AND  D( 8)='0' AND D( 1)='0' )then
          cVar2S2S107N069P064nsss(0) <='1';
          else
          cVar2S2S107N069P064nsss(0) <='0';
          end if;
        if(cVar1S3S107P052N065N010P067(0)='1' AND  A( 2)='1' )then
          cVar2S3S107P015nsss(0) <='1';
          else
          cVar2S3S107P015nsss(0) <='0';
          end if;
        if(cVar1S4S107P052N065N010P067(0)='1' AND  A( 2)='0' AND A( 4)='0' )then
          cVar2S4S107N015P011nsss(0) <='1';
          else
          cVar2S4S107N015P011nsss(0) <='0';
          end if;
        if(cVar1S5S107P052N065N010N067(0)='1' AND  A( 5)='1' AND B( 5)='1' )then
          cVar2S5S107P009P029nsss(0) <='1';
          else
          cVar2S5S107P009P029nsss(0) <='0';
          end if;
        if(cVar1S6S107P052N065N010N067(0)='1' AND  A( 5)='1' AND B( 5)='0' AND B( 6)='1' )then
          cVar2S6S107P009N029P027nsss(0) <='1';
          else
          cVar2S6S107P009N029P027nsss(0) <='0';
          end if;
        if(cVar1S7S107P052N065N010N067(0)='1' AND  A( 5)='0' AND A(15)='1' AND D( 5)='0' )then
          cVar2S7S107N009P008P048nsss(0) <='1';
          else
          cVar2S7S107N009P008P048nsss(0) <='0';
          end if;
        if(cVar1S8S107P052N065N010N067(0)='1' AND  A( 5)='0' AND A(15)='0' AND A( 4)='1' )then
          cVar2S8S107N009N008P011nsss(0) <='1';
          else
          cVar2S8S107N009N008P011nsss(0) <='0';
          end if;
        if(cVar1S10S107N052P044P025N005(0)='1' AND  A(16)='1' )then
          cVar2S10S107P006nsss(0) <='1';
          else
          cVar2S10S107P006nsss(0) <='0';
          end if;
        if(cVar1S11S107N052P044P025N005(0)='1' AND  A(16)='0' AND A( 6)='1' )then
          cVar2S11S107N006P007nsss(0) <='1';
          else
          cVar2S11S107N006P007nsss(0) <='0';
          end if;
        if(cVar1S13S107N052P044N025N067(0)='1' AND  E( 4)='1' )then
          cVar2S13S107P054nsss(0) <='1';
          else
          cVar2S13S107P054nsss(0) <='0';
          end if;
        if(cVar1S14S107N052P044N025N067(0)='1' AND  E( 4)='0' AND B( 8)='1' AND A( 7)='1' )then
          cVar2S14S107N054P023P005nsss(0) <='1';
          else
          cVar2S14S107N054P023P005nsss(0) <='0';
          end if;
        if(cVar1S15S107N052P044N025N067(0)='1' AND  E( 4)='0' AND B( 8)='0' AND E( 2)='1' )then
          cVar2S15S107N054N023P062nsss(0) <='1';
          else
          cVar2S15S107N054N023P062nsss(0) <='0';
          end if;
        if(cVar1S16S107N052N044P058P033(0)='1' AND  A(16)='1' AND E(14)='1' AND A(12)='0' )then
          cVar2S16S107P006P047P014nsss(0) <='1';
          else
          cVar2S16S107P006P047P014nsss(0) <='0';
          end if;
        if(cVar1S17S107N052N044P058P033(0)='1' AND  A(16)='1' AND E(14)='0' AND E(15)='1' )then
          cVar2S17S107P006N047P043nsss(0) <='1';
          else
          cVar2S17S107P006N047P043nsss(0) <='0';
          end if;
        if(cVar1S18S107N052N044P058P033(0)='1' AND  A(16)='0' AND D( 2)='1' AND B( 2)='1' )then
          cVar2S18S107N006P060P035nsss(0) <='1';
          else
          cVar2S18S107N006P060P035nsss(0) <='0';
          end if;
        if(cVar1S19S107N052N044P058P033(0)='1' AND  A(16)='0' AND B( 2)='1' AND B( 1)='0' )then
          cVar2S19S107P006P035P037nsss(0) <='1';
          else
          cVar2S19S107P006P035P037nsss(0) <='0';
          end if;
        if(cVar1S20S107N052N044P058P033(0)='1' AND  A( 3)='1' AND A(14)='0' AND A(12)='0' )then
          cVar2S20S107P013P010P014nsss(0) <='1';
          else
          cVar2S20S107P013P010P014nsss(0) <='0';
          end if;
        if(cVar1S21S107N052N044P058P033(0)='1' AND  A( 3)='0' AND A(13)='1' AND A( 2)='0' )then
          cVar2S21S107N013P012P015nsss(0) <='1';
          else
          cVar2S21S107N013P012P015nsss(0) <='0';
          end if;
        if(cVar1S22S107N052N044P058P033(0)='1' AND  A( 3)='0' AND A(13)='0' AND A(12)='1' )then
          cVar2S22S107N013N012P014nsss(0) <='1';
          else
          cVar2S22S107N013N012P014nsss(0) <='0';
          end if;
        if(cVar1S23S107N052N044P058N033(0)='1' AND  D( 3)='1' AND A(13)='1' )then
          cVar2S23S107P056P012nsss(0) <='1';
          else
          cVar2S23S107P056P012nsss(0) <='0';
          end if;
        if(cVar1S24S107N052N044P058N033(0)='1' AND  D( 3)='1' AND A(13)='0' AND A(14)='1' )then
          cVar2S24S107P056N012P010nsss(0) <='1';
          else
          cVar2S24S107P056N012P010nsss(0) <='0';
          end if;
        if(cVar1S25S107N052N044P058N033(0)='1' AND  D( 3)='0' AND A(12)='1' AND B( 1)='1' )then
          cVar2S25S107N056P014P037nsss(0) <='1';
          else
          cVar2S25S107N056P014P037nsss(0) <='0';
          end if;
        if(cVar1S26S107N052N044P058N033(0)='1' AND  D( 3)='0' AND A(12)='0' AND A(14)='1' )then
          cVar2S26S107N056N014P010nsss(0) <='1';
          else
          cVar2S26S107N056N014P010nsss(0) <='0';
          end if;
        if(cVar1S0S108P058P033P060P006(0)='1' AND  B(17)='1' AND A(12)='0' )then
          cVar2S0S108P024P014nsss(0) <='1';
          else
          cVar2S0S108P024P014nsss(0) <='0';
          end if;
        if(cVar1S1S108P058P033P060P006(0)='1' AND  B(17)='1' AND A(12)='1' AND A( 1)='0' )then
          cVar2S1S108P024P014P017nsss(0) <='1';
          else
          cVar2S1S108P024P014P017nsss(0) <='0';
          end if;
        if(cVar1S2S108P058P033P060P006(0)='1' AND  B(17)='0' )then
          cVar2S2S108N024psss(0) <='1';
          else
          cVar2S2S108N024psss(0) <='0';
          end if;
        if(cVar1S3S108P058P033P060N006(0)='1' AND  B( 5)='1' AND A( 4)='1' AND A(12)='0' )then
          cVar2S3S108P029P011P014nsss(0) <='1';
          else
          cVar2S3S108P029P011P014nsss(0) <='0';
          end if;
        if(cVar1S4S108P058P033P060N006(0)='1' AND  B( 5)='1' AND A( 4)='0' AND B(16)='0' )then
          cVar2S4S108P029N011P026nsss(0) <='1';
          else
          cVar2S4S108P029N011P026nsss(0) <='0';
          end if;
        if(cVar1S5S108P058P033P060N006(0)='1' AND  B( 5)='0' )then
          cVar2S5S108N029psss(0) <='1';
          else
          cVar2S5S108N029psss(0) <='0';
          end if;
        if(cVar1S6S108P058P033P060P066(0)='1' AND  E(10)='1' )then
          cVar2S6S108P063nsss(0) <='1';
          else
          cVar2S6S108P063nsss(0) <='0';
          end if;
        if(cVar1S7S108P058P033P060P066(0)='1' AND  E(10)='0' AND A(14)='0' AND A( 1)='0' )then
          cVar2S7S108N063P010P017nsss(0) <='1';
          else
          cVar2S7S108N063P010P017nsss(0) <='0';
          end if;
        if(cVar1S8S108P058P033P060N066(0)='1' AND  E( 2)='1' AND D( 1)='0' AND B( 2)='1' )then
          cVar2S8S108P062P064P035nsss(0) <='1';
          else
          cVar2S8S108P062P064P035nsss(0) <='0';
          end if;
        if(cVar1S9S108P058P033P060N066(0)='1' AND  E( 2)='1' AND D( 1)='1' AND B(12)='1' )then
          cVar2S9S108P062P064P034nsss(0) <='1';
          else
          cVar2S9S108P062P064P034nsss(0) <='0';
          end if;
        if(cVar1S10S108P058P033P060N066(0)='1' AND  E( 2)='0' AND A( 0)='1' AND A( 2)='1' )then
          cVar2S10S108N062P019P015nsss(0) <='1';
          else
          cVar2S10S108N062P019P015nsss(0) <='0';
          end if;
        if(cVar1S11S108P058P033P006P051(0)='1' AND  D( 8)='0' AND E( 1)='1' AND A( 8)='0' )then
          cVar2S11S108P069P066P003nsss(0) <='1';
          else
          cVar2S11S108P069P066P003nsss(0) <='0';
          end if;
        if(cVar1S12S108P058P033P006P051(0)='1' AND  D( 8)='0' AND E( 1)='0' AND E( 2)='1' )then
          cVar2S12S108P069N066P062nsss(0) <='1';
          else
          cVar2S12S108P069N066P062nsss(0) <='0';
          end if;
        if(cVar1S13S108P058P033P006P051(0)='1' AND  D( 8)='1' AND B(12)='1' )then
          cVar2S13S108P069P034nsss(0) <='1';
          else
          cVar2S13S108P069P034nsss(0) <='0';
          end if;
        if(cVar1S14S108P058P033P006P017(0)='1' AND  A( 0)='1' )then
          cVar2S14S108P019nsss(0) <='1';
          else
          cVar2S14S108P019nsss(0) <='0';
          end if;
        if(cVar1S15S108P058P006P013P033(0)='1' AND  A(14)='0' AND A(13)='0' AND D( 8)='0' )then
          cVar2S15S108P010P012P069nsss(0) <='1';
          else
          cVar2S15S108P010P012P069nsss(0) <='0';
          end if;
        if(cVar1S16S108P058P006P013P033(0)='1' AND  A(14)='0' AND A(13)='1' )then
          cVar2S16S108P010P012psss(0) <='1';
          else
          cVar2S16S108P010P012psss(0) <='0';
          end if;
        if(cVar1S17S108P058P006P013N033(0)='1' AND  B( 4)='1' AND A( 4)='0' )then
          cVar2S17S108P031P011nsss(0) <='1';
          else
          cVar2S17S108P031P011nsss(0) <='0';
          end if;
        if(cVar1S18S108P058P006P013N033(0)='1' AND  B( 4)='0' AND D( 1)='1' )then
          cVar2S18S108N031P064nsss(0) <='1';
          else
          cVar2S18S108N031P064nsss(0) <='0';
          end if;
        if(cVar1S19S108P058P006P013N033(0)='1' AND  B( 4)='0' AND D( 1)='0' AND E( 9)='1' )then
          cVar2S19S108N031N064P067nsss(0) <='1';
          else
          cVar2S19S108N031N064P067nsss(0) <='0';
          end if;
        if(cVar1S20S108P058P006N013P014(0)='1' AND  A( 5)='0' AND A( 2)='0' AND D( 2)='1' )then
          cVar2S20S108P009P015P060nsss(0) <='1';
          else
          cVar2S20S108P009P015P060nsss(0) <='0';
          end if;
        if(cVar1S21S108P058P006N013P014(0)='1' AND  A( 5)='0' AND A( 2)='1' AND B( 1)='1' )then
          cVar2S21S108P009P015P037nsss(0) <='1';
          else
          cVar2S21S108P009P015P037nsss(0) <='0';
          end if;
        if(cVar1S22S108P058P006N013N014(0)='1' AND  A(13)='1' AND A( 2)='0' AND D(10)='0' )then
          cVar2S22S108P012P015P061nsss(0) <='1';
          else
          cVar2S22S108P012P015P061nsss(0) <='0';
          end if;
        if(cVar1S23S108P058P006N013N014(0)='1' AND  A(13)='1' AND A( 2)='1' AND A(10)='1' )then
          cVar2S23S108P012P015P018nsss(0) <='1';
          else
          cVar2S23S108P012P015P018nsss(0) <='0';
          end if;
        if(cVar1S24S108P058P006N013N014(0)='1' AND  A(13)='0' AND A( 2)='1' AND B( 2)='0' )then
          cVar2S24S108N012P015P035nsss(0) <='1';
          else
          cVar2S24S108N012P015P035nsss(0) <='0';
          end if;
        if(cVar1S2S109P045N004P006N024(0)='1' AND  B(18)='1' )then
          cVar2S2S109P022nsss(0) <='1';
          else
          cVar2S2S109P022nsss(0) <='0';
          end if;
        if(cVar1S4S109P045N004N006N023(0)='1' AND  E( 5)='1' )then
          cVar2S4S109P050nsss(0) <='1';
          else
          cVar2S4S109P050nsss(0) <='0';
          end if;
        if(cVar1S5S109P045N004N006N023(0)='1' AND  E( 5)='0' AND A( 6)='1' )then
          cVar2S5S109N050P007nsss(0) <='1';
          else
          cVar2S5S109N050P007nsss(0) <='0';
          end if;
        if(cVar1S6S109P045N004N006N023(0)='1' AND  E( 5)='0' AND A( 6)='0' AND E(13)='1' )then
          cVar2S6S109N050N007P051nsss(0) <='1';
          else
          cVar2S6S109N050N007P051nsss(0) <='0';
          end if;
        if(cVar1S7S109N045P029P011P054(0)='1' AND  D(11)='0' AND E( 5)='0' AND A( 5)='0' )then
          cVar2S7S109P057P050P009nsss(0) <='1';
          else
          cVar2S7S109P057P050P009nsss(0) <='0';
          end if;
        if(cVar1S8S109N045P029P011P054(0)='1' AND  D(11)='0' AND E( 5)='1' AND D( 3)='1' )then
          cVar2S8S109P057P050P056nsss(0) <='1';
          else
          cVar2S8S109P057P050P056nsss(0) <='0';
          end if;
        if(cVar1S9S109N045P029P011N054(0)='1' AND  D(12)='1' )then
          cVar2S9S109P053nsss(0) <='1';
          else
          cVar2S9S109P053nsss(0) <='0';
          end if;
        if(cVar1S10S109N045P029P011N054(0)='1' AND  D(12)='0' AND E(12)='1' )then
          cVar2S10S109N053P055nsss(0) <='1';
          else
          cVar2S10S109N053P055nsss(0) <='0';
          end if;
        if(cVar1S11S109N045P029P011N054(0)='1' AND  D(12)='0' AND E(12)='0' AND D( 4)='1' )then
          cVar2S11S109N053N055P052nsss(0) <='1';
          else
          cVar2S11S109N053N055P052nsss(0) <='0';
          end if;
        if(cVar1S12S109N045P029N011P010(0)='1' AND  D( 4)='1' )then
          cVar2S12S109P052nsss(0) <='1';
          else
          cVar2S12S109P052nsss(0) <='0';
          end if;
        if(cVar1S13S109N045P029N011P010(0)='1' AND  D( 4)='0' AND E( 4)='1' )then
          cVar2S13S109N052P054nsss(0) <='1';
          else
          cVar2S13S109N052P054nsss(0) <='0';
          end if;
        if(cVar1S14S109N045P029N011N010(0)='1' AND  A( 5)='1' AND E( 5)='1' )then
          cVar2S14S109P009P050nsss(0) <='1';
          else
          cVar2S14S109P009P050nsss(0) <='0';
          end if;
        if(cVar1S15S109N045P029N011N010(0)='1' AND  A( 5)='1' AND E( 5)='0' AND E(13)='1' )then
          cVar2S15S109P009N050P051nsss(0) <='1';
          else
          cVar2S15S109P009N050P051nsss(0) <='0';
          end if;
        if(cVar1S16S109N045P029N011N010(0)='1' AND  A( 5)='0' AND A( 2)='1' AND A( 0)='0' )then
          cVar2S16S109N009P015P019nsss(0) <='1';
          else
          cVar2S16S109N009P015P019nsss(0) <='0';
          end if;
        if(cVar1S17S109N045N029P011P007(0)='1' AND  B( 7)='1' AND E( 6)='1' )then
          cVar2S17S109P025P046nsss(0) <='1';
          else
          cVar2S17S109P025P046nsss(0) <='0';
          end if;
        if(cVar1S18S109N045N029P011P007(0)='1' AND  B( 7)='1' AND E( 6)='0' AND E(14)='1' )then
          cVar2S18S109P025N046P047nsss(0) <='1';
          else
          cVar2S18S109P025N046P047nsss(0) <='0';
          end if;
        if(cVar1S19S109N045N029P011P007(0)='1' AND  B( 7)='0' AND B(15)='0' AND B( 6)='1' )then
          cVar2S19S109N025P028P027nsss(0) <='1';
          else
          cVar2S19S109N025P028P027nsss(0) <='0';
          end if;
        if(cVar1S20S109N045N029P011N007(0)='1' AND  E(14)='0' AND A( 5)='1' AND E(13)='1' )then
          cVar2S20S109P047P009P051nsss(0) <='1';
          else
          cVar2S20S109P047P009P051nsss(0) <='0';
          end if;
        if(cVar1S21S109N045N029P011N007(0)='1' AND  E(14)='1' AND A(16)='1' AND A(12)='0' )then
          cVar2S21S109P047P006P014nsss(0) <='1';
          else
          cVar2S21S109P047P006P014nsss(0) <='0';
          end if;
        if(cVar1S22S109N045N029P011N007(0)='1' AND  E(14)='1' AND A(16)='0' AND A(15)='1' )then
          cVar2S22S109P047N006P008nsss(0) <='1';
          else
          cVar2S22S109P047N006P008nsss(0) <='0';
          end if;
        if(cVar1S23S109N045N029P011P069(0)='1' AND  B( 4)='1' AND E( 4)='1' )then
          cVar2S23S109P031P054nsss(0) <='1';
          else
          cVar2S23S109P031P054nsss(0) <='0';
          end if;
        if(cVar1S24S109N045N029P011P069(0)='1' AND  B( 4)='1' AND E( 4)='0' AND A( 3)='0' )then
          cVar2S24S109P031N054P013nsss(0) <='1';
          else
          cVar2S24S109P031N054P013nsss(0) <='0';
          end if;
        if(cVar1S25S109N045N029P011P069(0)='1' AND  B( 4)='0' AND A( 3)='1' AND B( 1)='1' )then
          cVar2S25S109N031P013P037nsss(0) <='1';
          else
          cVar2S25S109N031P013P037nsss(0) <='0';
          end if;
        if(cVar1S26S109N045N029P011P069(0)='1' AND  B( 4)='0' AND A( 3)='0' AND B(15)='1' )then
          cVar2S26S109N031N013P028nsss(0) <='1';
          else
          cVar2S26S109N031N013P028nsss(0) <='0';
          end if;
        if(cVar1S27S109N045N029P011P069(0)='1' AND  B( 1)='1' AND D( 1)='0' )then
          cVar2S27S109P037P064nsss(0) <='1';
          else
          cVar2S27S109P037P064nsss(0) <='0';
          end if;
        if(cVar1S28S109N045N029P011P069(0)='1' AND  B( 1)='0' AND E(12)='1' )then
          cVar2S28S109N037P055nsss(0) <='1';
          else
          cVar2S28S109N037P055nsss(0) <='0';
          end if;
        if(cVar1S0S110P011P029P007P025(0)='1' AND  E( 6)='1' )then
          cVar2S0S110P046nsss(0) <='1';
          else
          cVar2S0S110P046nsss(0) <='0';
          end if;
        if(cVar1S1S110P011P029P007P025(0)='1' AND  E( 6)='0' AND E(14)='1' )then
          cVar2S1S110N046P047nsss(0) <='1';
          else
          cVar2S1S110N046P047nsss(0) <='0';
          end if;
        if(cVar1S2S110P011P029P007P025(0)='1' AND  E( 6)='0' AND E(14)='0' AND E( 7)='1' )then
          cVar2S2S110N046N047P042nsss(0) <='1';
          else
          cVar2S2S110N046N047P042nsss(0) <='0';
          end if;
        if(cVar1S3S110P011P029P007N025(0)='1' AND  B(15)='0' AND A( 5)='1' AND A(14)='0' )then
          cVar2S3S110P028P009P010nsss(0) <='1';
          else
          cVar2S3S110P028P009P010nsss(0) <='0';
          end if;
        if(cVar1S4S110P011P029P007N025(0)='1' AND  B(15)='0' AND A( 5)='0' )then
          cVar2S4S110P028N009psss(0) <='1';
          else
          cVar2S4S110P028N009psss(0) <='0';
          end if;
        if(cVar1S5S110P011P029N007P049(0)='1' AND  A( 5)='0' AND B( 6)='0' )then
          cVar2S5S110P009P027nsss(0) <='1';
          else
          cVar2S5S110P009P027nsss(0) <='0';
          end if;
        if(cVar1S6S110P011P029N007P049(0)='1' AND  A( 5)='0' AND B( 6)='1' AND A(15)='1' )then
          cVar2S6S110P009P027P008nsss(0) <='1';
          else
          cVar2S6S110P009P027P008nsss(0) <='0';
          end if;
        if(cVar1S7S110P011P029N007P049(0)='1' AND  A( 5)='1' AND E( 5)='1' AND B( 6)='1' )then
          cVar2S7S110P009P050P027nsss(0) <='1';
          else
          cVar2S7S110P009P050P027nsss(0) <='0';
          end if;
        if(cVar1S8S110P011P029N007P049(0)='1' AND  A( 5)='1' AND E( 5)='0' AND A( 3)='1' )then
          cVar2S8S110P009N050P013nsss(0) <='1';
          else
          cVar2S8S110P009N050P013nsss(0) <='0';
          end if;
        if(cVar1S9S110P011P029N007P049(0)='1' AND  A(16)='1' AND B(17)='1' )then
          cVar2S9S110P006P024nsss(0) <='1';
          else
          cVar2S9S110P006P024nsss(0) <='0';
          end if;
        if(cVar1S10S110P011P029N007P049(0)='1' AND  A(16)='1' AND B(17)='0' AND B(16)='1' )then
          cVar2S10S110P006N024P026nsss(0) <='1';
          else
          cVar2S10S110P006N024P026nsss(0) <='0';
          end if;
        if(cVar1S11S110P011P029N007P049(0)='1' AND  A(16)='0' AND A( 5)='1' AND E( 5)='0' )then
          cVar2S11S110N006P009P050nsss(0) <='1';
          else
          cVar2S11S110N006P009P050nsss(0) <='0';
          end if;
        if(cVar1S12S110P011P029N007P049(0)='1' AND  A(16)='0' AND A( 5)='0' AND A(15)='1' )then
          cVar2S12S110N006N009P008nsss(0) <='1';
          else
          cVar2S12S110N006N009P008nsss(0) <='0';
          end if;
        if(cVar1S13S110P011P029P005P010(0)='1' AND  D( 4)='1' )then
          cVar2S13S110P052nsss(0) <='1';
          else
          cVar2S13S110P052nsss(0) <='0';
          end if;
        if(cVar1S14S110P011P029P005P010(0)='1' AND  D( 4)='0' AND E( 4)='1' )then
          cVar2S14S110N052P054nsss(0) <='1';
          else
          cVar2S14S110N052P054nsss(0) <='0';
          end if;
        if(cVar1S15S110P011P029P005N010(0)='1' AND  A( 5)='1' )then
          cVar2S15S110P009nsss(0) <='1';
          else
          cVar2S15S110P009nsss(0) <='0';
          end if;
        if(cVar1S16S110P011P029P005N010(0)='1' AND  A( 5)='0' AND A( 3)='1' AND E( 4)='1' )then
          cVar2S16S110N009P013P054nsss(0) <='1';
          else
          cVar2S16S110N009P013P054nsss(0) <='0';
          end if;
        if(cVar1S17S110P011P029P005N010(0)='1' AND  A( 5)='0' AND A( 3)='0' AND A( 2)='1' )then
          cVar2S17S110N009N013P015nsss(0) <='1';
          else
          cVar2S17S110N009N013P015nsss(0) <='0';
          end if;
        if(cVar1S18S110P011P029P054P057(0)='1' AND  E( 5)='0' AND A(13)='0' )then
          cVar2S18S110P050P012nsss(0) <='1';
          else
          cVar2S18S110P050P012nsss(0) <='0';
          end if;
        if(cVar1S19S110P011P029P054P057(0)='1' AND  E( 5)='1' AND D( 3)='1' )then
          cVar2S19S110P050P056nsss(0) <='1';
          else
          cVar2S19S110P050P056nsss(0) <='0';
          end if;
        if(cVar1S21S110P011P029N054N053(0)='1' AND  E(12)='1' )then
          cVar2S21S110P055nsss(0) <='1';
          else
          cVar2S21S110P055nsss(0) <='0';
          end if;
        if(cVar1S22S110P011P029N054N053(0)='1' AND  E(12)='0' AND D( 4)='1' AND A(12)='0' )then
          cVar2S22S110N055P052P014nsss(0) <='1';
          else
          cVar2S22S110N055P052P014nsss(0) <='0';
          end if;
        if(cVar1S23S110P011N029P069P030(0)='1' AND  E(14)='1' AND B(16)='1' )then
          cVar2S23S110P047P026nsss(0) <='1';
          else
          cVar2S23S110P047P026nsss(0) <='0';
          end if;
        if(cVar1S24S110P011N029P069P030(0)='1' AND  E(14)='1' AND B(16)='0' AND A( 2)='1' )then
          cVar2S24S110P047N026P015nsss(0) <='1';
          else
          cVar2S24S110P047N026P015nsss(0) <='0';
          end if;
        if(cVar1S25S110P011N029P069P030(0)='1' AND  E(14)='0' AND B(19)='1' AND A(10)='0' )then
          cVar2S25S110N047P020P018nsss(0) <='1';
          else
          cVar2S25S110N047P020P018nsss(0) <='0';
          end if;
        if(cVar1S26S110P011N029P069P030(0)='1' AND  E(14)='0' AND B(19)='0' AND A(14)='0' )then
          cVar2S26S110N047N020P010nsss(0) <='1';
          else
          cVar2S26S110N047N020P010nsss(0) <='0';
          end if;
        if(cVar1S27S110P011N029P069P030(0)='1' AND  D( 3)='1' )then
          cVar2S27S110P056nsss(0) <='1';
          else
          cVar2S27S110P056nsss(0) <='0';
          end if;
        if(cVar1S28S110P011N029P069P030(0)='1' AND  D( 3)='0' AND D(11)='1' AND A(13)='0' )then
          cVar2S28S110N056P057P012nsss(0) <='1';
          else
          cVar2S28S110N056P057P012nsss(0) <='0';
          end if;
        if(cVar1S29S110P011N029P069P068(0)='1' AND  A(13)='1' )then
          cVar2S29S110P012nsss(0) <='1';
          else
          cVar2S29S110P012nsss(0) <='0';
          end if;
        if(cVar1S30S110P011N029P069P068(0)='1' AND  A(13)='0' AND A( 5)='0' AND B(11)='0' )then
          cVar2S30S110N012P009P036nsss(0) <='1';
          else
          cVar2S30S110N012P009P036nsss(0) <='0';
          end if;
        if(cVar1S31S110P011N029P069N068(0)='1' AND  A(10)='1' AND B( 2)='0' AND A( 2)='0' )then
          cVar2S31S110P018P035P015nsss(0) <='1';
          else
          cVar2S31S110P018P035P015nsss(0) <='0';
          end if;
        if(cVar1S32S110P011N029P069N068(0)='1' AND  A(10)='0' AND A(12)='0' AND A( 5)='1' )then
          cVar2S32S110N018P014P009nsss(0) <='1';
          else
          cVar2S32S110N018P014P009nsss(0) <='0';
          end if;
        if(cVar1S1S111P009P049N025P067(0)='1' AND  D( 0)='0' AND A( 0)='0' )then
          cVar2S1S111P068P019nsss(0) <='1';
          else
          cVar2S1S111P068P019nsss(0) <='0';
          end if;
        if(cVar1S3S111P009N049P053N029(0)='1' AND  A( 8)='0' AND E(10)='0' AND D( 0)='0' )then
          cVar2S3S111P003P063P068nsss(0) <='1';
          else
          cVar2S3S111P003P063P068nsss(0) <='0';
          end if;
        if(cVar1S4S111P009N049N053P050(0)='1' AND  B( 6)='1' AND A( 3)='0' )then
          cVar2S4S111P027P013nsss(0) <='1';
          else
          cVar2S4S111P027P013nsss(0) <='0';
          end if;
        if(cVar1S5S111P009N049N053P050(0)='1' AND  B( 6)='0' AND B( 5)='1' AND A( 4)='0' )then
          cVar2S5S111N027P029P011nsss(0) <='1';
          else
          cVar2S5S111N027P029P011nsss(0) <='0';
          end if;
        if(cVar1S6S111P009N049N053P050(0)='1' AND  B( 6)='0' AND B( 5)='0' AND A(11)='1' )then
          cVar2S6S111N027N029P016nsss(0) <='1';
          else
          cVar2S6S111N027N029P016nsss(0) <='0';
          end if;
        if(cVar1S7S111P009N049N053N050(0)='1' AND  A( 6)='1' AND B(11)='0' AND A(14)='0' )then
          cVar2S7S111P007P036P010nsss(0) <='1';
          else
          cVar2S7S111P007P036P010nsss(0) <='0';
          end if;
        if(cVar1S8S111P009N049N053N050(0)='1' AND  A( 6)='0' AND B( 6)='1' AND A( 3)='1' )then
          cVar2S8S111N007P027P013nsss(0) <='1';
          else
          cVar2S8S111N007P027P013nsss(0) <='0';
          end if;
        if(cVar1S11S111N009P044N004N051(0)='1' AND  B( 9)='1' )then
          cVar2S11S111P021nsss(0) <='1';
          else
          cVar2S11S111P021nsss(0) <='0';
          end if;
        if(cVar1S12S111N009P044N004N051(0)='1' AND  B( 9)='0' AND A( 4)='1' )then
          cVar2S12S111N021P011nsss(0) <='1';
          else
          cVar2S12S111N021P011nsss(0) <='0';
          end if;
        if(cVar1S13S111N009P044N004N051(0)='1' AND  B( 9)='0' AND A( 4)='0' AND A( 6)='1' )then
          cVar2S13S111N021N011P007nsss(0) <='1';
          else
          cVar2S13S111N021N011P007nsss(0) <='0';
          end if;
        if(cVar1S14S111N009N044P042P023(0)='1' AND  D( 0)='1' AND D( 8)='1' )then
          cVar2S14S111P068P069nsss(0) <='1';
          else
          cVar2S14S111P068P069nsss(0) <='0';
          end if;
        if(cVar1S15S111N009N044P042P023(0)='1' AND  D( 0)='0' AND B( 4)='1' AND A( 3)='1' )then
          cVar2S15S111N068P031P013nsss(0) <='1';
          else
          cVar2S15S111N068P031P013nsss(0) <='0';
          end if;
        if(cVar1S16S111N009N044P042P023(0)='1' AND  A(17)='0' AND E(15)='1' )then
          cVar2S16S111P004P043nsss(0) <='1';
          else
          cVar2S16S111P004P043nsss(0) <='0';
          end if;
        if(cVar1S17S111N009N044P042P023(0)='1' AND  A(17)='0' AND E(15)='0' AND D( 1)='1' )then
          cVar2S17S111P004N043P064nsss(0) <='1';
          else
          cVar2S17S111P004N043P064nsss(0) <='0';
          end if;
        if(cVar1S19S111N009N044P042N058(0)='1' AND  B( 8)='1' )then
          cVar2S19S111P023nsss(0) <='1';
          else
          cVar2S19S111P023nsss(0) <='0';
          end if;
        if(cVar1S20S111N009N044P042N058(0)='1' AND  B( 8)='0' AND B( 9)='1' AND A(18)='1' )then
          cVar2S20S111N023P021P002nsss(0) <='1';
          else
          cVar2S20S111N023P021P002nsss(0) <='0';
          end if;
        if(cVar1S1S112P009P049N025P067(0)='1' AND  D( 0)='0' AND A( 3)='0' )then
          cVar2S1S112P068P013nsss(0) <='1';
          else
          cVar2S1S112P068P013nsss(0) <='0';
          end if;
        if(cVar1S2S112P009N049P050P027(0)='1' AND  A( 4)='0' )then
          cVar2S2S112P011nsss(0) <='1';
          else
          cVar2S2S112P011nsss(0) <='0';
          end if;
        if(cVar1S3S112P009N049P050N027(0)='1' AND  B( 5)='1' AND A(11)='0' )then
          cVar2S3S112P029P016nsss(0) <='1';
          else
          cVar2S3S112P029P016nsss(0) <='0';
          end if;
        if(cVar1S4S112P009N049P050N027(0)='1' AND  B( 5)='0' AND E( 1)='1' )then
          cVar2S4S112N029P066nsss(0) <='1';
          else
          cVar2S4S112N029P066nsss(0) <='0';
          end if;
        if(cVar1S5S112P009N049P050N027(0)='1' AND  B( 5)='0' AND E( 1)='0' AND A( 2)='1' )then
          cVar2S5S112N029N066P015nsss(0) <='1';
          else
          cVar2S5S112N029N066P015nsss(0) <='0';
          end if;
        if(cVar1S6S112P009N049N050P053(0)='1' AND  B( 5)='1' )then
          cVar2S6S112P029nsss(0) <='1';
          else
          cVar2S6S112P029nsss(0) <='0';
          end if;
        if(cVar1S7S112P009N049N050P053(0)='1' AND  B( 5)='0' AND B( 2)='1' )then
          cVar2S7S112N029P035nsss(0) <='1';
          else
          cVar2S7S112N029P035nsss(0) <='0';
          end if;
        if(cVar1S8S112P009N049N050P053(0)='1' AND  B( 5)='0' AND B( 2)='0' AND A( 2)='0' )then
          cVar2S8S112N029N035P015nsss(0) <='1';
          else
          cVar2S8S112N029N035P015nsss(0) <='0';
          end if;
        if(cVar1S9S112P009N049N050N053(0)='1' AND  E(13)='0' AND A(14)='0' AND D( 0)='0' )then
          cVar2S9S112P051P010P068nsss(0) <='1';
          else
          cVar2S9S112P051P010P068nsss(0) <='0';
          end if;
        if(cVar1S10S112P009N049N050N053(0)='1' AND  E(13)='0' AND A(14)='1' AND D( 9)='1' )then
          cVar2S10S112P051P010P065nsss(0) <='1';
          else
          cVar2S10S112P051P010P065nsss(0) <='0';
          end if;
        if(cVar1S11S112N009P011P053P064(0)='1' AND  B(12)='0' AND D( 2)='0' AND E(11)='0' )then
          cVar2S11S112P034P060P059nsss(0) <='1';
          else
          cVar2S11S112P034P060P059nsss(0) <='0';
          end if;
        if(cVar1S12S112N009P011P053P064(0)='1' AND  B(12)='0' AND D( 2)='1' AND D( 0)='1' )then
          cVar2S12S112P034P060P068nsss(0) <='1';
          else
          cVar2S12S112P034P060P068nsss(0) <='0';
          end if;
        if(cVar1S13S112N009P011P053P064(0)='1' AND  B(12)='1' AND A(12)='1' AND A(11)='0' )then
          cVar2S13S112P034P014P016nsss(0) <='1';
          else
          cVar2S13S112P034P014P016nsss(0) <='0';
          end if;
        if(cVar1S14S112N009P011P053N064(0)='1' AND  B( 1)='0' AND E(11)='1' AND E( 3)='0' )then
          cVar2S14S112P037P059P058nsss(0) <='1';
          else
          cVar2S14S112P037P059P058nsss(0) <='0';
          end if;
        if(cVar1S15S112N009P011P053N064(0)='1' AND  B( 1)='0' AND E(11)='0' )then
          cVar2S15S112P037N059psss(0) <='1';
          else
          cVar2S15S112P037N059psss(0) <='0';
          end if;
        if(cVar1S16S112N009P011P053P036(0)='1' AND  E( 7)='1' )then
          cVar2S16S112P042nsss(0) <='1';
          else
          cVar2S16S112P042nsss(0) <='0';
          end if;
        if(cVar1S17S112N009P011P053P036(0)='1' AND  E( 7)='0' AND A( 7)='1' )then
          cVar2S17S112N042P005nsss(0) <='1';
          else
          cVar2S17S112N042P005nsss(0) <='0';
          end if;
        if(cVar1S18S112N009P011P053P036(0)='1' AND  E( 7)='0' AND A( 7)='0' AND B(19)='1' )then
          cVar2S18S112N042N005P020nsss(0) <='1';
          else
          cVar2S18S112N042N005P020nsss(0) <='0';
          end if;
        if(cVar1S19S112N009P011P053P036(0)='1' AND  A( 0)='0' AND A( 2)='1' )then
          cVar2S19S112P019P015nsss(0) <='1';
          else
          cVar2S19S112P019P015nsss(0) <='0';
          end if;
        if(cVar1S20S112N009P011P029P054(0)='1' AND  A( 1)='1' )then
          cVar2S20S112P017nsss(0) <='1';
          else
          cVar2S20S112P017nsss(0) <='0';
          end if;
        if(cVar1S21S112N009P011P029P054(0)='1' AND  A( 1)='0' AND A(12)='0' AND E( 5)='0' )then
          cVar2S21S112N017P014P050nsss(0) <='1';
          else
          cVar2S21S112N017P014P050nsss(0) <='0';
          end if;
        if(cVar1S22S112N009P011P029N054(0)='1' AND  D(12)='1' )then
          cVar2S22S112P053nsss(0) <='1';
          else
          cVar2S22S112P053nsss(0) <='0';
          end if;
        if(cVar1S23S112N009P011P029N054(0)='1' AND  D(12)='0' AND E(12)='1' )then
          cVar2S23S112N053P055nsss(0) <='1';
          else
          cVar2S23S112N053P055nsss(0) <='0';
          end if;
        if(cVar1S24S112N009P011P029N054(0)='1' AND  D(12)='0' AND E(12)='0' AND D( 4)='1' )then
          cVar2S24S112N053N055P052nsss(0) <='1';
          else
          cVar2S24S112N053N055P052nsss(0) <='0';
          end if;
        if(cVar1S25S112N009P011N029P047(0)='1' AND  B(16)='1' )then
          cVar2S25S112P026nsss(0) <='1';
          else
          cVar2S25S112P026nsss(0) <='0';
          end if;
        if(cVar1S26S112N009P011N029P047(0)='1' AND  B(16)='0' AND E( 1)='1' )then
          cVar2S26S112N026P066nsss(0) <='1';
          else
          cVar2S26S112N026P066nsss(0) <='0';
          end if;
        if(cVar1S27S112N009P011N029P047(0)='1' AND  B(16)='0' AND E( 1)='0' AND B(17)='0' )then
          cVar2S27S112N026N066P024nsss(0) <='1';
          else
          cVar2S27S112N026N066P024nsss(0) <='0';
          end if;
        if(cVar1S28S112N009P011N029N047(0)='1' AND  B(19)='1' AND D(15)='1' )then
          cVar2S28S112P020P041nsss(0) <='1';
          else
          cVar2S28S112P020P041nsss(0) <='0';
          end if;
        if(cVar1S29S112N009P011N029N047(0)='1' AND  B(19)='1' AND D(15)='0' AND A(10)='0' )then
          cVar2S29S112P020N041P018nsss(0) <='1';
          else
          cVar2S29S112P020N041P018nsss(0) <='0';
          end if;
        if(cVar1S30S112N009P011N029N047(0)='1' AND  B(19)='0' AND B( 0)='0' AND A( 3)='1' )then
          cVar2S30S112N020P039P013nsss(0) <='1';
          else
          cVar2S30S112N020P039P013nsss(0) <='0';
          end if;
        if(cVar1S1S113P037P066P027N047(0)='1' AND  D( 5)='0' AND E( 7)='0' AND B( 8)='0' )then
          cVar2S1S113P048P042P023nsss(0) <='1';
          else
          cVar2S1S113P048P042P023nsss(0) <='0';
          end if;
        if(cVar1S2S113P037P066P027N047(0)='1' AND  D( 5)='1' AND A( 1)='0' AND E( 6)='1' )then
          cVar2S2S113P048P017P046nsss(0) <='1';
          else
          cVar2S2S113P048P017P046nsss(0) <='0';
          end if;
        if(cVar1S3S113P037P066P027P068(0)='1' AND  A(10)='0' )then
          cVar2S3S113P018nsss(0) <='1';
          else
          cVar2S3S113P018nsss(0) <='0';
          end if;
        if(cVar1S4S113P037N066P069P068(0)='1' AND  D( 2)='0' AND D( 1)='0' AND B( 2)='0' )then
          cVar2S4S113P060P064P035nsss(0) <='1';
          else
          cVar2S4S113P060P064P035nsss(0) <='0';
          end if;
        if(cVar1S5S113P037N066P069P068(0)='1' AND  D( 2)='0' AND D( 1)='1' AND B(11)='1' )then
          cVar2S5S113P060P064P036nsss(0) <='1';
          else
          cVar2S5S113P060P064P036nsss(0) <='0';
          end if;
        if(cVar1S6S113P037N066N069P035(0)='1' AND  E( 2)='0' )then
          cVar2S6S113P062nsss(0) <='1';
          else
          cVar2S6S113P062nsss(0) <='0';
          end if;
        if(cVar1S7S113P037N066N069P035(0)='1' AND  E( 2)='1' AND D( 1)='1' AND A( 2)='0' )then
          cVar2S7S113P062P064P015nsss(0) <='1';
          else
          cVar2S7S113P062P064P015nsss(0) <='0';
          end if;
        if(cVar1S8S113P037N066N069N035(0)='1' AND  B( 9)='1' )then
          cVar2S8S113P021nsss(0) <='1';
          else
          cVar2S8S113P021nsss(0) <='0';
          end if;
        if(cVar1S9S113P037N066N069N035(0)='1' AND  B( 9)='0' AND A(10)='1' AND D(10)='0' )then
          cVar2S9S113N021P018P061nsss(0) <='1';
          else
          cVar2S9S113N021P018P061nsss(0) <='0';
          end if;
        if(cVar1S10S113P037N066N069N035(0)='1' AND  B( 9)='0' AND A(10)='0' AND E( 3)='1' )then
          cVar2S10S113N021N018P058nsss(0) <='1';
          else
          cVar2S10S113N021N018P058nsss(0) <='0';
          end if;
        if(cVar1S12S113N037P059N043P058(0)='1' AND  A(19)='0' AND E(12)='0' AND D( 9)='0' )then
          cVar2S12S113P000P055P065nsss(0) <='1';
          else
          cVar2S12S113P000P055P065nsss(0) <='0';
          end if;
        if(cVar1S13S113N037P059N043P058(0)='1' AND  E( 9)='1' )then
          cVar2S13S113P067nsss(0) <='1';
          else
          cVar2S13S113P067nsss(0) <='0';
          end if;
        if(cVar1S14S113N037P059N043P058(0)='1' AND  E( 9)='0' AND D( 2)='1' AND D(11)='1' )then
          cVar2S14S113N067P060P057nsss(0) <='1';
          else
          cVar2S14S113N067P060P057nsss(0) <='0';
          end if;
        if(cVar1S15S113N037N059P009P049(0)='1' AND  B( 7)='1' )then
          cVar2S15S113P025nsss(0) <='1';
          else
          cVar2S15S113P025nsss(0) <='0';
          end if;
        if(cVar1S16S113N037N059P009P049(0)='1' AND  B( 7)='0' AND A( 0)='0' )then
          cVar2S16S113N025P019nsss(0) <='1';
          else
          cVar2S16S113N025P019nsss(0) <='0';
          end if;
        if(cVar1S17S113N037N059P009P049(0)='1' AND  B( 7)='0' AND A( 0)='1' AND B( 6)='1' )then
          cVar2S17S113N025P019P027nsss(0) <='1';
          else
          cVar2S17S113N025P019P027nsss(0) <='0';
          end if;
        if(cVar1S18S113N037N059P009N049(0)='1' AND  D(11)='1' AND B(15)='1' )then
          cVar2S18S113P057P028nsss(0) <='1';
          else
          cVar2S18S113P057P028nsss(0) <='0';
          end if;
        if(cVar1S19S113N037N059P009N049(0)='1' AND  D(11)='1' AND B(15)='0' AND E(12)='1' )then
          cVar2S19S113P057N028P055nsss(0) <='1';
          else
          cVar2S19S113P057N028P055nsss(0) <='0';
          end if;
        if(cVar1S20S113N037N059P009N049(0)='1' AND  D(11)='0' AND B( 6)='1' AND A(10)='0' )then
          cVar2S20S113N057P027P018nsss(0) <='1';
          else
          cVar2S20S113N057P027P018nsss(0) <='0';
          end if;
        if(cVar1S21S113N037N059P009N049(0)='1' AND  D(11)='0' AND B( 6)='0' AND D( 9)='1' )then
          cVar2S21S113N057N027P065nsss(0) <='1';
          else
          cVar2S21S113N057N027P065nsss(0) <='0';
          end if;
        if(cVar1S22S113N037N059N009P054(0)='1' AND  A(14)='1' AND A( 0)='0' )then
          cVar2S22S113P010P019nsss(0) <='1';
          else
          cVar2S22S113P010P019nsss(0) <='0';
          end if;
        if(cVar1S23S113N037N059N009P054(0)='1' AND  A(14)='1' AND A( 0)='1' AND A(11)='0' )then
          cVar2S23S113P010P019P016nsss(0) <='1';
          else
          cVar2S23S113P010P019P016nsss(0) <='0';
          end if;
        if(cVar1S24S113N037N059N009P054(0)='1' AND  A(14)='0' AND A( 4)='1' AND B( 5)='1' )then
          cVar2S24S113N010P011P029nsss(0) <='1';
          else
          cVar2S24S113N010P011P029nsss(0) <='0';
          end if;
        if(cVar1S25S113N037N059N009P054(0)='1' AND  A(14)='0' AND A( 4)='0' AND A( 3)='1' )then
          cVar2S25S113N010N011P013nsss(0) <='1';
          else
          cVar2S25S113N010N011P013nsss(0) <='0';
          end if;
        if(cVar1S26S113N037N059N009N054(0)='1' AND  B( 4)='0' AND A(11)='1' AND A( 1)='1' )then
          cVar2S26S113P031P016P017nsss(0) <='1';
          else
          cVar2S26S113P031P016P017nsss(0) <='0';
          end if;
        if(cVar1S27S113N037N059N009N054(0)='1' AND  B( 4)='0' AND A(11)='0' AND D( 1)='1' )then
          cVar2S27S113P031N016P064nsss(0) <='1';
          else
          cVar2S27S113P031N016P064nsss(0) <='0';
          end if;
        if(cVar1S28S113N037N059N009N054(0)='1' AND  B( 4)='1' AND E( 3)='1' AND A( 0)='0' )then
          cVar2S28S113P031P058P019nsss(0) <='1';
          else
          cVar2S28S113P031P058P019nsss(0) <='0';
          end if;
        if(cVar1S0S114P064P037P005P043(0)='1' AND  A( 3)='0' )then
          cVar2S0S114P013nsss(0) <='1';
          else
          cVar2S0S114P013nsss(0) <='0';
          end if;
        if(cVar1S1S114P064P037P005N043(0)='1' AND  A( 6)='1' AND A( 5)='0' )then
          cVar2S1S114P007P009nsss(0) <='1';
          else
          cVar2S1S114P007P009nsss(0) <='0';
          end if;
        if(cVar1S2S114P064P037P005N043(0)='1' AND  A( 6)='0' AND D( 8)='0' AND D( 0)='0' )then
          cVar2S2S114N007P069P068nsss(0) <='1';
          else
          cVar2S2S114N007P069P068nsss(0) <='0';
          end if;
        if(cVar1S3S114P064P037P005N043(0)='1' AND  A( 6)='0' AND D( 8)='1' AND A(13)='1' )then
          cVar2S3S114N007P069P012nsss(0) <='1';
          else
          cVar2S3S114N007P069P012nsss(0) <='0';
          end if;
        if(cVar1S4S114P064P037N005P028(0)='1' AND  D(12)='1' AND A(13)='0' )then
          cVar2S4S114P053P012nsss(0) <='1';
          else
          cVar2S4S114P053P012nsss(0) <='0';
          end if;
        if(cVar1S5S114P064P037N005P028(0)='1' AND  D(12)='1' AND A(13)='1' AND A(14)='1' )then
          cVar2S5S114P053P012P010nsss(0) <='1';
          else
          cVar2S5S114P053P012P010nsss(0) <='0';
          end if;
        if(cVar1S6S114P064P037N005P028(0)='1' AND  D(12)='0' AND A(13)='1' AND E(12)='0' )then
          cVar2S6S114N053P012P055nsss(0) <='1';
          else
          cVar2S6S114N053P012P055nsss(0) <='0';
          end if;
        if(cVar1S7S114P064P037N005P028(0)='1' AND  D(12)='0' AND A(13)='0' AND D(11)='1' )then
          cVar2S7S114N053N012P057nsss(0) <='1';
          else
          cVar2S7S114N053N012P057nsss(0) <='0';
          end if;
        if(cVar1S8S114P064P037N005N028(0)='1' AND  B( 5)='1' AND E( 4)='1' AND D(11)='0' )then
          cVar2S8S114P029P054P057nsss(0) <='1';
          else
          cVar2S8S114P029P054P057nsss(0) <='0';
          end if;
        if(cVar1S9S114P064P037N005N028(0)='1' AND  B( 5)='1' AND E( 4)='0' AND B( 3)='0' )then
          cVar2S9S114P029N054P033nsss(0) <='1';
          else
          cVar2S9S114P029N054P033nsss(0) <='0';
          end if;
        if(cVar1S10S114P064P037N005N028(0)='1' AND  B( 5)='0' AND B(16)='1' AND D( 8)='0' )then
          cVar2S10S114N029P026P069nsss(0) <='1';
          else
          cVar2S10S114N029P026P069nsss(0) <='0';
          end if;
        if(cVar1S11S114P064P037N005N028(0)='1' AND  B( 5)='0' AND B(16)='0' AND D(13)='0' )then
          cVar2S11S114N029N026P049nsss(0) <='1';
          else
          cVar2S11S114N029N026P049nsss(0) <='0';
          end if;
        if(cVar1S12S114P064P037P061P012(0)='1' AND  A( 3)='1' AND A(11)='0' )then
          cVar2S12S114P013P016nsss(0) <='1';
          else
          cVar2S12S114P013P016nsss(0) <='0';
          end if;
        if(cVar1S13S114P064P037P061P012(0)='1' AND  A( 3)='1' AND A(11)='1' AND E( 1)='0' )then
          cVar2S13S114P013P016P066nsss(0) <='1';
          else
          cVar2S13S114P013P016P066nsss(0) <='0';
          end if;
        if(cVar1S14S114P064P037P061P012(0)='1' AND  A( 3)='0' AND D( 3)='1' )then
          cVar2S14S114N013P056nsss(0) <='1';
          else
          cVar2S14S114N013P056nsss(0) <='0';
          end if;
        if(cVar1S15S114P064P037P061P012(0)='1' AND  A( 3)='0' AND D( 3)='0' AND A(16)='1' )then
          cVar2S15S114N013N056P006nsss(0) <='1';
          else
          cVar2S15S114N013N056P006nsss(0) <='0';
          end if;
        if(cVar1S16S114P064P037P061N012(0)='1' AND  D( 0)='1' AND A(19)='0' AND E( 4)='0' )then
          cVar2S16S114P068P000P054nsss(0) <='1';
          else
          cVar2S16S114P068P000P054nsss(0) <='0';
          end if;
        if(cVar1S17S114P064P037P061N012(0)='1' AND  D( 0)='0' AND D( 8)='1' AND B(11)='0' )then
          cVar2S17S114N068P069P036nsss(0) <='1';
          else
          cVar2S17S114N068P069P036nsss(0) <='0';
          end if;
        if(cVar1S19S114P064P037P061N062(0)='1' AND  D( 8)='1' )then
          cVar2S19S114P069nsss(0) <='1';
          else
          cVar2S19S114P069nsss(0) <='0';
          end if;
        if(cVar1S20S114P064P037P061N062(0)='1' AND  D( 8)='0' AND A(11)='1' AND E(11)='0' )then
          cVar2S20S114N069P016P059nsss(0) <='1';
          else
          cVar2S20S114N069P016P059nsss(0) <='0';
          end if;
        if(cVar1S23S114P064N046N042P003(0)='1' AND  B(11)='1' AND E( 1)='1' )then
          cVar2S23S114P036P066nsss(0) <='1';
          else
          cVar2S23S114P036P066nsss(0) <='0';
          end if;
        if(cVar1S24S114P064N046N042P003(0)='1' AND  B(11)='0' AND A( 4)='1' AND E( 4)='1' )then
          cVar2S24S114N036P011P054nsss(0) <='1';
          else
          cVar2S24S114N036P011P054nsss(0) <='0';
          end if;
        if(cVar1S25S114P064N046N042P003(0)='1' AND  A( 6)='0' AND B(11)='1' AND A( 1)='1' )then
          cVar2S25S114P007P036P017nsss(0) <='1';
          else
          cVar2S25S114P007P036P017nsss(0) <='0';
          end if;
        if(cVar1S26S114P064N046N042P003(0)='1' AND  A( 6)='0' AND B(11)='0' AND A(14)='1' )then
          cVar2S26S114P007N036P010nsss(0) <='1';
          else
          cVar2S26S114P007N036P010nsss(0) <='0';
          end if;
        if(cVar1S1S115P049P026P033N007(0)='1' AND  A( 4)='1' )then
          cVar2S1S115P011nsss(0) <='1';
          else
          cVar2S1S115P011nsss(0) <='0';
          end if;
        if(cVar1S2S115P049P026P033N007(0)='1' AND  A( 4)='0' AND B(17)='0' )then
          cVar2S2S115N011P024nsss(0) <='1';
          else
          cVar2S2S115N011P024nsss(0) <='0';
          end if;
        if(cVar1S4S115P049N026P024N004(0)='1' AND  A(16)='1' AND A(12)='0' )then
          cVar2S4S115P006P014nsss(0) <='1';
          else
          cVar2S4S115P006P014nsss(0) <='0';
          end if;
        if(cVar1S5S115P049N026P024N004(0)='1' AND  A(16)='0' AND A( 7)='1' )then
          cVar2S5S115N006P005nsss(0) <='1';
          else
          cVar2S5S115N006P005nsss(0) <='0';
          end if;
        if(cVar1S6S115P049N026P024N004(0)='1' AND  A(16)='0' AND A( 7)='0' AND A( 6)='1' )then
          cVar2S6S115N006N005P007nsss(0) <='1';
          else
          cVar2S6S115N006N005P007nsss(0) <='0';
          end if;
        if(cVar1S7S115P049N026N024P027(0)='1' AND  D( 5)='0' )then
          cVar2S7S115P048nsss(0) <='1';
          else
          cVar2S7S115P048nsss(0) <='0';
          end if;
        if(cVar1S8S115P049N026N024P027(0)='1' AND  D( 5)='1' AND E(14)='0' )then
          cVar2S8S115P048P047nsss(0) <='1';
          else
          cVar2S8S115P048P047nsss(0) <='0';
          end if;
        if(cVar1S9S115P049N026N024P027(0)='1' AND  D( 5)='1' AND E(14)='1' AND E( 5)='1' )then
          cVar2S9S115P048P047P050nsss(0) <='1';
          else
          cVar2S9S115P048P047P050nsss(0) <='0';
          end if;
        if(cVar1S10S115P049N026N024N027(0)='1' AND  E(14)='0' AND B( 3)='1' )then
          cVar2S10S115P047P033nsss(0) <='1';
          else
          cVar2S10S115P047P033nsss(0) <='0';
          end if;
        if(cVar1S11S115P049N026N024N027(0)='1' AND  E(14)='0' AND B( 3)='0' AND B(12)='1' )then
          cVar2S11S115P047N033P034nsss(0) <='1';
          else
          cVar2S11S115P047N033P034nsss(0) <='0';
          end if;
        if(cVar1S12S115P049N026N024N027(0)='1' AND  E(14)='1' AND B( 7)='1' )then
          cVar2S12S115P047P025nsss(0) <='1';
          else
          cVar2S12S115P047P025nsss(0) <='0';
          end if;
        if(cVar1S14S115N049P064P050N065(0)='1' AND  A(10)='1' )then
          cVar2S14S115P018nsss(0) <='1';
          else
          cVar2S14S115P018nsss(0) <='0';
          end if;
        if(cVar1S15S115N049P064P050N065(0)='1' AND  A(10)='0' AND A(11)='0' AND A( 1)='1' )then
          cVar2S15S115N018P016P017nsss(0) <='1';
          else
          cVar2S15S115N018P016P017nsss(0) <='0';
          end if;
        if(cVar1S16S115N049P064N050P008(0)='1' AND  A( 7)='0' AND E(11)='0' )then
          cVar2S16S115P005P059nsss(0) <='1';
          else
          cVar2S16S115P005P059nsss(0) <='0';
          end if;
        if(cVar1S17S115N049P064N050P008(0)='1' AND  A( 7)='0' AND E(11)='1' AND E( 3)='1' )then
          cVar2S17S115P005P059P058nsss(0) <='1';
          else
          cVar2S17S115P005P059P058nsss(0) <='0';
          end if;
        if(cVar1S18S115N049P064N050P008(0)='1' AND  A( 7)='1' AND A( 0)='1' AND B( 1)='1' )then
          cVar2S18S115P005P019P037nsss(0) <='1';
          else
          cVar2S18S115P005P019P037nsss(0) <='0';
          end if;
        if(cVar1S19S115N049P064N050P008(0)='1' AND  A(14)='0' AND A( 0)='1' AND B( 1)='0' )then
          cVar2S19S115P010P019P037nsss(0) <='1';
          else
          cVar2S19S115P010P019P037nsss(0) <='0';
          end if;
        if(cVar1S20S115N049P064N050P008(0)='1' AND  A(14)='0' AND A( 0)='0' AND B(12)='1' )then
          cVar2S20S115P010N019P034nsss(0) <='1';
          else
          cVar2S20S115P010N019P034nsss(0) <='0';
          end if;
        if(cVar1S21S115N049N064P047P028(0)='1' AND  D(12)='1' AND E(10)='0' )then
          cVar2S21S115P053P063nsss(0) <='1';
          else
          cVar2S21S115P053P063nsss(0) <='0';
          end if;
        if(cVar1S22S115N049N064P047P028(0)='1' AND  D(12)='0' AND D(11)='1' )then
          cVar2S22S115N053P057nsss(0) <='1';
          else
          cVar2S22S115N053P057nsss(0) <='0';
          end if;
        if(cVar1S23S115N049N064P047P028(0)='1' AND  D(12)='0' AND D(11)='0' AND E( 4)='1' )then
          cVar2S23S115N053N057P054nsss(0) <='1';
          else
          cVar2S23S115N053N057P054nsss(0) <='0';
          end if;
        if(cVar1S24S115N049N064P047N028(0)='1' AND  B( 5)='1' AND E(10)='0' )then
          cVar2S24S115P029P063nsss(0) <='1';
          else
          cVar2S24S115P029P063nsss(0) <='0';
          end if;
        if(cVar1S25S115N049N064P047N028(0)='1' AND  B( 5)='0' AND A( 7)='1' AND D( 9)='0' )then
          cVar2S25S115N029P005P065nsss(0) <='1';
          else
          cVar2S25S115N029P005P065nsss(0) <='0';
          end if;
        if(cVar1S26S115N049N064P047N028(0)='1' AND  B( 5)='0' AND A( 7)='0' AND D( 2)='1' )then
          cVar2S26S115N029N005P060nsss(0) <='1';
          else
          cVar2S26S115N029N005P060nsss(0) <='0';
          end if;
        if(cVar1S28S115N049N064P047N069(0)='1' AND  D(14)='1' AND A(17)='1' )then
          cVar2S28S115P045P004nsss(0) <='1';
          else
          cVar2S28S115P045P004nsss(0) <='0';
          end if;
        if(cVar1S29S115N049N064P047N069(0)='1' AND  D(14)='1' AND A(17)='0' AND A( 0)='1' )then
          cVar2S29S115P045N004P019nsss(0) <='1';
          else
          cVar2S29S115P045N004P019nsss(0) <='0';
          end if;
        if(cVar1S30S115N049N064P047N069(0)='1' AND  D(14)='0' AND A(12)='0' AND A(15)='1' )then
          cVar2S30S115N045P014P008nsss(0) <='1';
          else
          cVar2S30S115N045P014P008nsss(0) <='0';
          end if;
        if(cVar1S0S116P060P062P049P024(0)='1' AND  A(17)='1' )then
          cVar2S0S116P004nsss(0) <='1';
          else
          cVar2S0S116P004nsss(0) <='0';
          end if;
        if(cVar1S1S116P060P062P049P024(0)='1' AND  A(17)='0' AND A(16)='1' AND A(12)='0' )then
          cVar2S1S116N004P006P014nsss(0) <='1';
          else
          cVar2S1S116N004P006P014nsss(0) <='0';
          end if;
        if(cVar1S2S116P060P062P049P024(0)='1' AND  A(17)='0' AND A(16)='0' )then
          cVar2S2S116N004N006psss(0) <='1';
          else
          cVar2S2S116N004N006psss(0) <='0';
          end if;
        if(cVar1S3S116P060P062P049N024(0)='1' AND  B(16)='1' )then
          cVar2S3S116P026nsss(0) <='1';
          else
          cVar2S3S116P026nsss(0) <='0';
          end if;
        if(cVar1S4S116P060P062P049N024(0)='1' AND  B(16)='0' AND B( 6)='1' )then
          cVar2S4S116N026P027nsss(0) <='1';
          else
          cVar2S4S116N026P027nsss(0) <='0';
          end if;
        if(cVar1S5S116P060P062N049P047(0)='1' AND  D( 1)='0' AND E( 7)='0' )then
          cVar2S5S116P064P042nsss(0) <='1';
          else
          cVar2S5S116P064P042nsss(0) <='0';
          end if;
        if(cVar1S6S116P060P062N049P047(0)='1' AND  D( 1)='0' AND E( 7)='1' AND A(18)='1' )then
          cVar2S6S116P064P042P002nsss(0) <='1';
          else
          cVar2S6S116P064P042P002nsss(0) <='0';
          end if;
        if(cVar1S7S116P060P062N049P047(0)='1' AND  D( 1)='1' AND E( 1)='1' AND B(12)='0' )then
          cVar2S7S116P064P066P034nsss(0) <='1';
          else
          cVar2S7S116P064P066P034nsss(0) <='0';
          end if;
        if(cVar1S8S116P060P062N049P047(0)='1' AND  D(14)='1' AND A(17)='1' )then
          cVar2S8S116P045P004nsss(0) <='1';
          else
          cVar2S8S116P045P004nsss(0) <='0';
          end if;
        if(cVar1S9S116P060P062N049P047(0)='1' AND  D(14)='1' AND A(17)='0' AND A( 2)='1' )then
          cVar2S9S116P045N004P015nsss(0) <='1';
          else
          cVar2S9S116P045N004P015nsss(0) <='0';
          end if;
        if(cVar1S10S116P060P062N049P047(0)='1' AND  D(14)='0' AND D( 8)='1' )then
          cVar2S10S116N045P069nsss(0) <='1';
          else
          cVar2S10S116N045P069nsss(0) <='0';
          end if;
        if(cVar1S12S116P060P062N050P068(0)='1' AND  A( 6)='0' AND B( 7)='0' AND A( 8)='0' )then
          cVar2S12S116P007P025P003nsss(0) <='1';
          else
          cVar2S12S116P007P025P003nsss(0) <='0';
          end if;
        if(cVar1S13S116P060P062N050P068(0)='1' AND  A( 6)='1' AND D( 9)='1' )then
          cVar2S13S116P007P065nsss(0) <='1';
          else
          cVar2S13S116P007P065nsss(0) <='0';
          end if;
        if(cVar1S14S116P060P062N050P068(0)='1' AND  D(11)='1' )then
          cVar2S14S116P057nsss(0) <='1';
          else
          cVar2S14S116P057nsss(0) <='0';
          end if;
        if(cVar1S15S116P060P062N050P068(0)='1' AND  D(11)='0' AND B(16)='1' )then
          cVar2S15S116N057P026nsss(0) <='1';
          else
          cVar2S15S116N057P026nsss(0) <='0';
          end if;
        if(cVar1S16S116P060P062N050P068(0)='1' AND  D(11)='0' AND B(16)='0' AND B(12)='1' )then
          cVar2S16S116N057N026P034nsss(0) <='1';
          else
          cVar2S16S116N057N026P034nsss(0) <='0';
          end if;
        if(cVar1S18S116P060P014P008N032(0)='1' AND  A( 2)='0' AND A(13)='0' AND E( 9)='0' )then
          cVar2S18S116P015P012P067nsss(0) <='1';
          else
          cVar2S18S116P015P012P067nsss(0) <='0';
          end if;
        if(cVar1S19S116P060P014P008N032(0)='1' AND  A( 2)='1' AND D( 1)='1' )then
          cVar2S19S116P015P064nsss(0) <='1';
          else
          cVar2S19S116P015P064nsss(0) <='0';
          end if;
        if(cVar1S20S116P060N014P033P013(0)='1' AND  A( 0)='0' AND E( 9)='0' )then
          cVar2S20S116P019P067nsss(0) <='1';
          else
          cVar2S20S116P019P067nsss(0) <='0';
          end if;
        if(cVar1S21S116P060N014P033P013(0)='1' AND  A( 0)='1' AND A(10)='1' )then
          cVar2S21S116P019P018nsss(0) <='1';
          else
          cVar2S21S116P019P018nsss(0) <='0';
          end if;
        if(cVar1S22S116P060N014P033P013(0)='1' AND  A( 0)='1' AND A(10)='0' AND A( 1)='0' )then
          cVar2S22S116P019N018P017nsss(0) <='1';
          else
          cVar2S22S116P019N018P017nsss(0) <='0';
          end if;
        if(cVar1S23S116P060N014P033N013(0)='1' AND  A( 2)='1' AND E( 9)='1' )then
          cVar2S23S116P015P067nsss(0) <='1';
          else
          cVar2S23S116P015P067nsss(0) <='0';
          end if;
        if(cVar1S24S116P060N014P033N013(0)='1' AND  A( 2)='1' AND E( 9)='0' AND D(10)='1' )then
          cVar2S24S116P015N067P061nsss(0) <='1';
          else
          cVar2S24S116P015N067P061nsss(0) <='0';
          end if;
        if(cVar1S25S116P060N014P033N013(0)='1' AND  A( 2)='0' AND A(13)='1' )then
          cVar2S25S116N015P012nsss(0) <='1';
          else
          cVar2S25S116N015P012nsss(0) <='0';
          end if;
        if(cVar1S26S116P060N014N033P066(0)='1' AND  A(11)='1' )then
          cVar2S26S116P016nsss(0) <='1';
          else
          cVar2S26S116P016nsss(0) <='0';
          end if;
        if(cVar1S27S116P060N014N033P066(0)='1' AND  A(11)='0' AND E( 3)='0' AND A( 2)='0' )then
          cVar2S27S116N016P058P015nsss(0) <='1';
          else
          cVar2S27S116N016P058P015nsss(0) <='0';
          end if;
        if(cVar1S28S116P060N014N033N066(0)='1' AND  B( 4)='1' AND A(14)='1' )then
          cVar2S28S116P031P010nsss(0) <='1';
          else
          cVar2S28S116P031P010nsss(0) <='0';
          end if;
        if(cVar1S29S116P060N014N033N066(0)='1' AND  B( 4)='1' AND A(14)='0' AND A( 3)='1' )then
          cVar2S29S116P031N010P013nsss(0) <='1';
          else
          cVar2S29S116P031N010P013nsss(0) <='0';
          end if;
        if(cVar1S30S116P060N014N033N066(0)='1' AND  B( 4)='0' AND B( 2)='1' AND D( 1)='0' )then
          cVar2S30S116N031P035P064nsss(0) <='1';
          else
          cVar2S30S116N031P035P064nsss(0) <='0';
          end if;
        if(cVar1S31S116P060N014N033N066(0)='1' AND  B( 4)='0' AND B( 2)='0' AND E(14)='1' )then
          cVar2S31S116N031N035P047nsss(0) <='1';
          else
          cVar2S31S116N031N035P047nsss(0) <='0';
          end if;
        if(cVar1S2S117P049N005N026P024(0)='1' AND  A(17)='1' )then
          cVar2S2S117P004nsss(0) <='1';
          else
          cVar2S2S117P004nsss(0) <='0';
          end if;
        if(cVar1S3S117P049N005N026P024(0)='1' AND  A(17)='0' AND A(16)='1' AND A(15)='0' )then
          cVar2S3S117N004P006P008nsss(0) <='1';
          else
          cVar2S3S117N004P006P008nsss(0) <='0';
          end if;
        if(cVar1S4S117P049N005N026P024(0)='1' AND  A(17)='0' AND A(16)='0' AND A( 6)='1' )then
          cVar2S4S117N004N006P007nsss(0) <='1';
          else
          cVar2S4S117N004N006P007nsss(0) <='0';
          end if;
        if(cVar1S5S117P049N005N026N024(0)='1' AND  B( 6)='1' )then
          cVar2S5S117P027nsss(0) <='1';
          else
          cVar2S5S117P027nsss(0) <='0';
          end if;
        if(cVar1S6S117P049N005N026N024(0)='1' AND  B( 6)='0' AND E(14)='0' AND B( 3)='1' )then
          cVar2S6S117N027P047P033nsss(0) <='1';
          else
          cVar2S6S117N027P047P033nsss(0) <='0';
          end if;
        if(cVar1S7S117P049N005N026N024(0)='1' AND  B( 6)='0' AND E(14)='1' AND B( 7)='1' )then
          cVar2S7S117N027P047P025nsss(0) <='1';
          else
          cVar2S7S117N027P047P025nsss(0) <='0';
          end if;
        if(cVar1S8S117N049P024P053P028(0)='1' AND  A(12)='0' )then
          cVar2S8S117P014nsss(0) <='1';
          else
          cVar2S8S117P014nsss(0) <='0';
          end if;
        if(cVar1S9S117N049P024P053P028(0)='1' AND  A(12)='1' AND A(11)='1' )then
          cVar2S9S117P014P016nsss(0) <='1';
          else
          cVar2S9S117P014P016nsss(0) <='0';
          end if;
        if(cVar1S10S117N049P024P053N028(0)='1' AND  B(16)='1' AND E( 1)='0' AND A( 4)='0' )then
          cVar2S10S117P026P066P011nsss(0) <='1';
          else
          cVar2S10S117P026P066P011nsss(0) <='0';
          end if;
        if(cVar1S11S117N049P024P053N028(0)='1' AND  B(16)='0' AND B( 5)='1' )then
          cVar2S11S117N026P029nsss(0) <='1';
          else
          cVar2S11S117N026P029nsss(0) <='0';
          end if;
        if(cVar1S12S117N049P024P053N028(0)='1' AND  B(16)='0' AND B( 5)='0' AND D( 5)='1' )then
          cVar2S12S117N026N029P048nsss(0) <='1';
          else
          cVar2S12S117N026N029P048nsss(0) <='0';
          end if;
        if(cVar1S13S117N049P024N053P051(0)='1' AND  B( 7)='1' AND D( 5)='1' AND E( 9)='0' )then
          cVar2S13S117P025P048P067nsss(0) <='1';
          else
          cVar2S13S117P025P048P067nsss(0) <='0';
          end if;
        if(cVar1S14S117N049P024N053P051(0)='1' AND  B( 7)='1' AND D( 5)='0' AND E(15)='1' )then
          cVar2S14S117P025N048P043nsss(0) <='1';
          else
          cVar2S14S117P025N048P043nsss(0) <='0';
          end if;
        if(cVar1S15S117N049P024N053P051(0)='1' AND  B( 7)='0' AND E( 6)='0' AND D( 4)='1' )then
          cVar2S15S117N025P046P052nsss(0) <='1';
          else
          cVar2S15S117N025P046P052nsss(0) <='0';
          end if;
        if(cVar1S16S117N049P024N053P051(0)='1' AND  B( 7)='0' AND E( 6)='1' AND B(14)='1' )then
          cVar2S16S117N025P046P030nsss(0) <='1';
          else
          cVar2S16S117N025P046P030nsss(0) <='0';
          end if;
        if(cVar1S17S117N049P024N053P051(0)='1' AND  D( 4)='0' AND A( 1)='1' )then
          cVar2S17S117P052P017nsss(0) <='1';
          else
          cVar2S17S117P052P017nsss(0) <='0';
          end if;
        if(cVar1S18S117N049P024N053P051(0)='1' AND  D( 4)='0' AND A( 1)='0' AND D(10)='1' )then
          cVar2S18S117P052N017P061nsss(0) <='1';
          else
          cVar2S18S117P052N017P061nsss(0) <='0';
          end if;
        if(cVar1S20S117N049P024P026N002(0)='1' AND  D( 0)='0' AND A(16)='1' )then
          cVar2S20S117P068P006nsss(0) <='1';
          else
          cVar2S20S117P068P006nsss(0) <='0';
          end if;
        if(cVar1S2S118P049N006P007P019(0)='1' AND  B(11)='0' )then
          cVar2S2S118P036nsss(0) <='1';
          else
          cVar2S2S118P036nsss(0) <='0';
          end if;
        if(cVar1S3S118P049N006P007P019(0)='1' AND  A( 1)='1' )then
          cVar2S3S118P017nsss(0) <='1';
          else
          cVar2S3S118P017nsss(0) <='0';
          end if;
        if(cVar1S4S118P049N006N007P009(0)='1' AND  B( 7)='1' )then
          cVar2S4S118P025nsss(0) <='1';
          else
          cVar2S4S118P025nsss(0) <='0';
          end if;
        if(cVar1S5S118P049N006N007P009(0)='1' AND  B( 7)='0' AND D( 0)='0' AND A( 1)='0' )then
          cVar2S5S118N025P068P017nsss(0) <='1';
          else
          cVar2S5S118N025P068P017nsss(0) <='0';
          end if;
        if(cVar1S6S118P049N006N007N009(0)='1' AND  A( 7)='1' )then
          cVar2S6S118P005nsss(0) <='1';
          else
          cVar2S6S118P005nsss(0) <='0';
          end if;
        if(cVar1S7S118P049N006N007N009(0)='1' AND  A( 7)='0' AND A(15)='1' AND A(14)='0' )then
          cVar2S7S118N005P008P010nsss(0) <='1';
          else
          cVar2S7S118N005P008P010nsss(0) <='0';
          end if;
        if(cVar1S8S118P049N006N007N009(0)='1' AND  A( 7)='0' AND A(15)='0' AND E(14)='0' )then
          cVar2S8S118N005N008P047nsss(0) <='1';
          else
          cVar2S8S118N005N008P047nsss(0) <='0';
          end if;
        if(cVar1S9S118N049P052P024P042(0)='1' AND  E( 3)='1' )then
          cVar2S9S118P058nsss(0) <='1';
          else
          cVar2S9S118P058nsss(0) <='0';
          end if;
        if(cVar1S10S118N049P052P024P042(0)='1' AND  E( 3)='0' AND B( 0)='1' )then
          cVar2S10S118N058P039nsss(0) <='1';
          else
          cVar2S10S118N058P039nsss(0) <='0';
          end if;
        if(cVar1S11S118N049P052P024P042(0)='1' AND  E( 3)='0' AND B( 0)='0' AND B( 8)='1' )then
          cVar2S11S118N058N039P023nsss(0) <='1';
          else
          cVar2S11S118N058N039P023nsss(0) <='0';
          end if;
        if(cVar1S12S118N049P052P024N042(0)='1' AND  A( 7)='0' AND A(17)='0' AND E(15)='0' )then
          cVar2S12S118P005P004P043nsss(0) <='1';
          else
          cVar2S12S118P005P004P043nsss(0) <='0';
          end if;
        if(cVar1S13S118N049P052P024N042(0)='1' AND  A( 7)='1' AND A(12)='1' )then
          cVar2S13S118P005P014nsss(0) <='1';
          else
          cVar2S13S118P005P014nsss(0) <='0';
          end if;
        if(cVar1S14S118N049P052P024N042(0)='1' AND  A( 7)='1' AND A(12)='0' AND B(10)='1' )then
          cVar2S14S118P005N014P038nsss(0) <='1';
          else
          cVar2S14S118P005N014P038nsss(0) <='0';
          end if;
        if(cVar1S15S118N049P052P024P068(0)='1' AND  D(11)='0' AND A(17)='1' )then
          cVar2S15S118P057P004nsss(0) <='1';
          else
          cVar2S15S118P057P004nsss(0) <='0';
          end if;
        if(cVar1S16S118N049P052P024P068(0)='1' AND  D(11)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S16S118P057N004P006nsss(0) <='1';
          else
          cVar2S16S118P057N004P006nsss(0) <='0';
          end if;
        if(cVar1S17S118N049P052P024P068(0)='1' AND  A(11)='0' AND A( 4)='1' )then
          cVar2S17S118P016P011nsss(0) <='1';
          else
          cVar2S17S118P016P011nsss(0) <='0';
          end if;
        if(cVar1S19S118N049P052N065P067(0)='1' AND  A( 2)='1' )then
          cVar2S19S118P015nsss(0) <='1';
          else
          cVar2S19S118P015nsss(0) <='0';
          end if;
        if(cVar1S20S118N049P052N065P067(0)='1' AND  A( 2)='0' AND A( 4)='0' )then
          cVar2S20S118N015P011nsss(0) <='1';
          else
          cVar2S20S118N015P011nsss(0) <='0';
          end if;
        if(cVar1S21S118N049P052N065N067(0)='1' AND  A(14)='1' AND A( 8)='0' AND A(12)='0' )then
          cVar2S21S118P010P003P014nsss(0) <='1';
          else
          cVar2S21S118P010P003P014nsss(0) <='0';
          end if;
        if(cVar1S22S118N049P052N065N067(0)='1' AND  A(14)='0' AND A( 5)='1' AND A( 0)='1' )then
          cVar2S22S118N010P009P019nsss(0) <='1';
          else
          cVar2S22S118N010P009P019nsss(0) <='0';
          end if;
        if(cVar1S23S118N049P052N065N067(0)='1' AND  A(14)='0' AND A( 5)='0' AND A(15)='1' )then
          cVar2S23S118N010N009P008nsss(0) <='1';
          else
          cVar2S23S118N010N009P008nsss(0) <='0';
          end if;
        if(cVar1S1S119P049P006P007P018(0)='1' AND  A( 1)='1' )then
          cVar2S1S119P017nsss(0) <='1';
          else
          cVar2S1S119P017nsss(0) <='0';
          end if;
        if(cVar1S3S119P049N006P007N025(0)='1' AND  A( 0)='0' )then
          cVar2S3S119P019nsss(0) <='1';
          else
          cVar2S3S119P019nsss(0) <='0';
          end if;
        if(cVar1S4S119P049N006N007P009(0)='1' AND  B( 7)='1' )then
          cVar2S4S119P025nsss(0) <='1';
          else
          cVar2S4S119P025nsss(0) <='0';
          end if;
        if(cVar1S5S119P049N006N007P009(0)='1' AND  B( 7)='0' AND E(13)='0' AND E(14)='1' )then
          cVar2S5S119N025P051P047nsss(0) <='1';
          else
          cVar2S5S119N025P051P047nsss(0) <='0';
          end if;
        if(cVar1S6S119P049N006N007P009(0)='1' AND  B( 7)='0' AND E(13)='1' AND E(14)='0' )then
          cVar2S6S119N025P051P047nsss(0) <='1';
          else
          cVar2S6S119N025P051P047nsss(0) <='0';
          end if;
        if(cVar1S7S119P049N006N007N009(0)='1' AND  A( 7)='1' )then
          cVar2S7S119P005nsss(0) <='1';
          else
          cVar2S7S119P005nsss(0) <='0';
          end if;
        if(cVar1S8S119P049N006N007N009(0)='1' AND  A( 7)='0' AND A(15)='1' AND B(16)='1' )then
          cVar2S8S119N005P008P026nsss(0) <='1';
          else
          cVar2S8S119N005P008P026nsss(0) <='0';
          end if;
        if(cVar1S10S119N049P042N051P050(0)='1' AND  A(17)='1' )then
          cVar2S10S119P004nsss(0) <='1';
          else
          cVar2S10S119P004nsss(0) <='0';
          end if;
        if(cVar1S11S119N049P042N051P050(0)='1' AND  A(17)='0' AND B( 0)='1' )then
          cVar2S11S119N004P039nsss(0) <='1';
          else
          cVar2S11S119N004P039nsss(0) <='0';
          end if;
        if(cVar1S12S119N049P042N051P050(0)='1' AND  A(17)='0' AND B( 0)='0' AND A( 7)='1' )then
          cVar2S12S119N004N039P005nsss(0) <='1';
          else
          cVar2S12S119N004N039P005nsss(0) <='0';
          end if;
        if(cVar1S14S119N049N042P045N022(0)='1' AND  D( 5)='1' )then
          cVar2S14S119P048nsss(0) <='1';
          else
          cVar2S14S119P048nsss(0) <='0';
          end if;
        if(cVar1S15S119N049N042P045N022(0)='1' AND  D( 5)='0' AND E(10)='1' )then
          cVar2S15S119N048P063nsss(0) <='1';
          else
          cVar2S15S119N048P063nsss(0) <='0';
          end if;
        if(cVar1S16S119N049N042P045N022(0)='1' AND  D( 5)='0' AND E(10)='0' AND D(10)='1' )then
          cVar2S16S119N048N063P061nsss(0) <='1';
          else
          cVar2S16S119N048N063P061nsss(0) <='0';
          end if;
        if(cVar1S17S119N049N042N045P047(0)='1' AND  B( 8)='0' AND B(19)='1' AND A( 8)='1' )then
          cVar2S17S119P023P020P003nsss(0) <='1';
          else
          cVar2S17S119P023P020P003nsss(0) <='0';
          end if;
        if(cVar1S18S119N049N042N045P047(0)='1' AND  B( 8)='1' AND D( 3)='1' )then
          cVar2S18S119P023P056nsss(0) <='1';
          else
          cVar2S18S119P023P056nsss(0) <='0';
          end if;
        if(cVar1S19S119N049N042N045P047(0)='1' AND  B( 8)='1' AND D( 3)='0' AND D(15)='1' )then
          cVar2S19S119P023N056P041nsss(0) <='1';
          else
          cVar2S19S119P023N056P041nsss(0) <='0';
          end if;
        if(cVar1S20S119N049N042N045P047(0)='1' AND  D( 8)='1' )then
          cVar2S20S119P069nsss(0) <='1';
          else
          cVar2S20S119P069nsss(0) <='0';
          end if;
        if(cVar1S0S120P049P024P010P006(0)='1' AND  A(10)='0' )then
          cVar2S0S120P018nsss(0) <='1';
          else
          cVar2S0S120P018nsss(0) <='0';
          end if;
        if(cVar1S1S120P049P024P010P006(0)='1' AND  A(10)='1' AND A( 0)='0' )then
          cVar2S1S120P018P019nsss(0) <='1';
          else
          cVar2S1S120P018P019nsss(0) <='0';
          end if;
        if(cVar1S2S120P049P024P010N006(0)='1' AND  A(11)='0' AND A(10)='0' )then
          cVar2S2S120P016P018nsss(0) <='1';
          else
          cVar2S2S120P016P018nsss(0) <='0';
          end if;
        if(cVar1S4S120P049N024P026N007(0)='1' AND  A(15)='1' AND A( 0)='0' )then
          cVar2S4S120P008P019nsss(0) <='1';
          else
          cVar2S4S120P008P019nsss(0) <='0';
          end if;
        if(cVar1S5S120P049N024P026N007(0)='1' AND  A(15)='0' AND A( 4)='1' )then
          cVar2S5S120N008P011nsss(0) <='1';
          else
          cVar2S5S120N008P011nsss(0) <='0';
          end if;
        if(cVar1S6S120P049N024P026N007(0)='1' AND  A(15)='0' AND A( 4)='0' AND A(16)='1' )then
          cVar2S6S120N008N011P006nsss(0) <='1';
          else
          cVar2S6S120N008N011P006nsss(0) <='0';
          end if;
        if(cVar1S8S120P049N024N026N027(0)='1' AND  E(14)='0' AND B(12)='1' )then
          cVar2S8S120P047P034nsss(0) <='1';
          else
          cVar2S8S120P047P034nsss(0) <='0';
          end if;
        if(cVar1S9S120P049N024N026N027(0)='1' AND  E(14)='0' AND B(12)='0' AND B( 3)='1' )then
          cVar2S9S120P047N034P033nsss(0) <='1';
          else
          cVar2S9S120P047N034P033nsss(0) <='0';
          end if;
        if(cVar1S10S120P049N024N026N027(0)='1' AND  E(14)='1' AND B( 7)='1' )then
          cVar2S10S120P047P025nsss(0) <='1';
          else
          cVar2S10S120P047P025nsss(0) <='0';
          end if;
        if(cVar1S11S120N049P042P050P004(0)='1' AND  B( 8)='1' )then
          cVar2S11S120P023nsss(0) <='1';
          else
          cVar2S11S120P023nsss(0) <='0';
          end if;
        if(cVar1S12S120N049P042P050P004(0)='1' AND  B( 8)='0' AND D( 7)='1' )then
          cVar2S12S120N023P040nsss(0) <='1';
          else
          cVar2S12S120N023P040nsss(0) <='0';
          end if;
        if(cVar1S13S120N049P042P050P004(0)='1' AND  B( 8)='0' AND D( 7)='0' AND B(18)='1' )then
          cVar2S13S120N023N040P022nsss(0) <='1';
          else
          cVar2S13S120N023N040P022nsss(0) <='0';
          end if;
        if(cVar1S14S120N049P042P050N004(0)='1' AND  A(18)='1' )then
          cVar2S14S120P002nsss(0) <='1';
          else
          cVar2S14S120P002nsss(0) <='0';
          end if;
        if(cVar1S15S120N049P042P050N004(0)='1' AND  A(18)='0' AND E( 3)='1' )then
          cVar2S15S120N002P058nsss(0) <='1';
          else
          cVar2S15S120N002P058nsss(0) <='0';
          end if;
        if(cVar1S16S120N049P042P050N004(0)='1' AND  A(18)='0' AND E( 3)='0' AND B( 7)='1' )then
          cVar2S16S120N002N058P025nsss(0) <='1';
          else
          cVar2S16S120N002N058P025nsss(0) <='0';
          end if;
        if(cVar1S18S120N049N042P045N022(0)='1' AND  B( 8)='1' AND A( 1)='0' )then
          cVar2S18S120P023P017nsss(0) <='1';
          else
          cVar2S18S120P023P017nsss(0) <='0';
          end if;
        if(cVar1S19S120N049N042P045N022(0)='1' AND  B( 8)='0' AND A( 8)='0' AND B(17)='1' )then
          cVar2S19S120N023P003P024nsss(0) <='1';
          else
          cVar2S19S120N023P003P024nsss(0) <='0';
          end if;
        if(cVar1S20S120N049N042N045P047(0)='1' AND  B( 8)='0' )then
          cVar2S20S120P023nsss(0) <='1';
          else
          cVar2S20S120P023nsss(0) <='0';
          end if;
        if(cVar1S21S120N049N042N045P047(0)='1' AND  B( 8)='1' AND D( 3)='1' )then
          cVar2S21S120P023P056nsss(0) <='1';
          else
          cVar2S21S120P023P056nsss(0) <='0';
          end if;
        if(cVar1S22S120N049N042N045P047(0)='1' AND  B( 8)='1' AND D( 3)='0' AND D(15)='1' )then
          cVar2S22S120P023N056P041nsss(0) <='1';
          else
          cVar2S22S120P023N056P041nsss(0) <='0';
          end if;
        if(cVar1S23S120N049N042N045P047(0)='1' AND  B(16)='0' AND E( 9)='1' )then
          cVar2S23S120P026P067nsss(0) <='1';
          else
          cVar2S23S120P026P067nsss(0) <='0';
          end if;
        if(cVar1S1S121P049P024P010N006(0)='1' AND  A(11)='0' AND A(10)='0' )then
          cVar2S1S121P016P018nsss(0) <='1';
          else
          cVar2S1S121P016P018nsss(0) <='0';
          end if;
        if(cVar1S3S121P049N024P026N007(0)='1' AND  A(15)='1' AND A( 0)='0' )then
          cVar2S3S121P008P019nsss(0) <='1';
          else
          cVar2S3S121P008P019nsss(0) <='0';
          end if;
        if(cVar1S4S121P049N024P026N007(0)='1' AND  A(15)='0' AND A( 4)='1' )then
          cVar2S4S121N008P011nsss(0) <='1';
          else
          cVar2S4S121N008P011nsss(0) <='0';
          end if;
        if(cVar1S5S121P049N024P026N007(0)='1' AND  A(15)='0' AND A( 4)='0' AND A(16)='1' )then
          cVar2S5S121N008N011P006nsss(0) <='1';
          else
          cVar2S5S121N008N011P006nsss(0) <='0';
          end if;
        if(cVar1S7S121P049N024N026N027(0)='1' AND  E(14)='0' AND A( 1)='1' )then
          cVar2S7S121P047P017nsss(0) <='1';
          else
          cVar2S7S121P047P017nsss(0) <='0';
          end if;
        if(cVar1S8S121P049N024N026N027(0)='1' AND  E(14)='0' AND A( 1)='0' AND A(12)='0' )then
          cVar2S8S121P047N017P014nsss(0) <='1';
          else
          cVar2S8S121P047N017P014nsss(0) <='0';
          end if;
        if(cVar1S9S121P049N024N026N027(0)='1' AND  E(14)='1' AND B( 7)='1' )then
          cVar2S9S121P047P025nsss(0) <='1';
          else
          cVar2S9S121P047P025nsss(0) <='0';
          end if;
        if(cVar1S12S121N049N042P045P004(0)='1' AND  A( 3)='0' AND B(18)='1' )then
          cVar2S12S121P013P022nsss(0) <='1';
          else
          cVar2S12S121P013P022nsss(0) <='0';
          end if;
        if(cVar1S13S121N049N042P045N004(0)='1' AND  A(12)='1' AND A( 3)='0' )then
          cVar2S13S121P014P013nsss(0) <='1';
          else
          cVar2S13S121P014P013nsss(0) <='0';
          end if;
        if(cVar1S14S121N049N042P045N004(0)='1' AND  A(12)='0' AND E(13)='1' )then
          cVar2S14S121N014P051nsss(0) <='1';
          else
          cVar2S14S121N014P051nsss(0) <='0';
          end if;
        if(cVar1S15S121N049N042P045N004(0)='1' AND  A(12)='0' AND E(13)='0' AND D( 2)='1' )then
          cVar2S15S121N014N051P060nsss(0) <='1';
          else
          cVar2S15S121N014N051P060nsss(0) <='0';
          end if;
        if(cVar1S16S121N049N042N045P047(0)='1' AND  A(13)='1' AND D( 3)='1' AND B(14)='1' )then
          cVar2S16S121P012P056P030nsss(0) <='1';
          else
          cVar2S16S121P012P056P030nsss(0) <='0';
          end if;
        if(cVar1S17S121N049N042N045P047(0)='1' AND  A(13)='0' AND D(15)='1' )then
          cVar2S17S121N012P041nsss(0) <='1';
          else
          cVar2S17S121N012P041nsss(0) <='0';
          end if;
        if(cVar1S18S121N049N042N045P047(0)='1' AND  B(16)='0' AND E( 9)='1' )then
          cVar2S18S121P026P067nsss(0) <='1';
          else
          cVar2S18S121P026P067nsss(0) <='0';
          end if;
        if(cVar1S1S122P045P027P024N013(0)='1' AND  A(16)='1' )then
          cVar2S1S122P006nsss(0) <='1';
          else
          cVar2S1S122P006nsss(0) <='0';
          end if;
        if(cVar1S2S122P045P027P024N013(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S2S122N006P004nsss(0) <='1';
          else
          cVar2S2S122N006P004nsss(0) <='0';
          end if;
        if(cVar1S3S122P045P027P024N013(0)='1' AND  A(16)='0' AND A(17)='0' AND E(14)='1' )then
          cVar2S3S122N006N004P047nsss(0) <='1';
          else
          cVar2S3S122N006N004P047nsss(0) <='0';
          end if;
        if(cVar1S4S122P045P027N024P025(0)='1' AND  E(15)='1' )then
          cVar2S4S122P043nsss(0) <='1';
          else
          cVar2S4S122P043nsss(0) <='0';
          end if;
        if(cVar1S5S122P045P027N024P025(0)='1' AND  E(15)='0' AND E( 6)='1' )then
          cVar2S5S122N043P046nsss(0) <='1';
          else
          cVar2S5S122N043P046nsss(0) <='0';
          end if;
        if(cVar1S6S122P045P027N024N025(0)='1' AND  B(18)='1' )then
          cVar2S6S122P022nsss(0) <='1';
          else
          cVar2S6S122P022nsss(0) <='0';
          end if;
        if(cVar1S7S122P045P027N024N025(0)='1' AND  B(18)='0' AND B( 8)='1' AND A( 1)='0' )then
          cVar2S7S122N022P023P017nsss(0) <='1';
          else
          cVar2S7S122N022P023P017nsss(0) <='0';
          end if;
        if(cVar1S8S122P045P027N024N025(0)='1' AND  B(18)='0' AND B( 8)='0' AND E(15)='0' )then
          cVar2S8S122N022N023P043nsss(0) <='1';
          else
          cVar2S8S122N022N023P043nsss(0) <='0';
          end if;
        if(cVar1S9S122N045P049P024P026(0)='1' AND  A(17)='1' )then
          cVar2S9S122P004nsss(0) <='1';
          else
          cVar2S9S122P004nsss(0) <='0';
          end if;
        if(cVar1S10S122N045P049P024P026(0)='1' AND  A(17)='0' AND A( 1)='0' )then
          cVar2S10S122N004P017nsss(0) <='1';
          else
          cVar2S10S122N004P017nsss(0) <='0';
          end if;
        if(cVar1S11S122N045P049P024P026(0)='1' AND  A(17)='0' AND A( 1)='1' AND A(10)='1' )then
          cVar2S11S122N004P017P018nsss(0) <='1';
          else
          cVar2S11S122N004P017P018nsss(0) <='0';
          end if;
        if(cVar1S12S122N045P049N024P026(0)='1' AND  A( 6)='1' )then
          cVar2S12S122P007nsss(0) <='1';
          else
          cVar2S12S122P007nsss(0) <='0';
          end if;
        if(cVar1S13S122N045P049N024P026(0)='1' AND  A( 6)='0' AND A(15)='1' AND A( 0)='0' )then
          cVar2S13S122N007P008P019nsss(0) <='1';
          else
          cVar2S13S122N007P008P019nsss(0) <='0';
          end if;
        if(cVar1S14S122N045P049N024P026(0)='1' AND  A( 6)='0' AND A(15)='0' AND A( 4)='1' )then
          cVar2S14S122N007N008P011nsss(0) <='1';
          else
          cVar2S14S122N007N008P011nsss(0) <='0';
          end if;
        if(cVar1S15S122N045P049N024N026(0)='1' AND  B( 6)='1' )then
          cVar2S15S122P027nsss(0) <='1';
          else
          cVar2S15S122P027nsss(0) <='0';
          end if;
        if(cVar1S16S122N045P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='0' )then
          cVar2S16S122N027P047nsss(0) <='1';
          else
          cVar2S16S122N027P047nsss(0) <='0';
          end if;
        if(cVar1S17S122N045P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='1' AND B( 7)='1' )then
          cVar2S17S122N027P047P025nsss(0) <='1';
          else
          cVar2S17S122N027P047P025nsss(0) <='0';
          end if;
        if(cVar1S18S122N045N049P047P042(0)='1' AND  E(13)='1' )then
          cVar2S18S122P051nsss(0) <='1';
          else
          cVar2S18S122P051nsss(0) <='0';
          end if;
        if(cVar1S19S122N045N049P047P042(0)='1' AND  E(13)='0' AND A(17)='1' )then
          cVar2S19S122N051P004nsss(0) <='1';
          else
          cVar2S19S122N051P004nsss(0) <='0';
          end if;
        if(cVar1S20S122N045N049P047P042(0)='1' AND  E(13)='0' AND A(17)='0' AND A(18)='1' )then
          cVar2S20S122N051N004P002nsss(0) <='1';
          else
          cVar2S20S122N051N004P002nsss(0) <='0';
          end if;
        if(cVar1S21S122N045N049P047N042(0)='1' AND  A(13)='1' AND D( 3)='1' )then
          cVar2S21S122P012P056nsss(0) <='1';
          else
          cVar2S21S122P012P056nsss(0) <='0';
          end if;
        if(cVar1S22S122N045N049P047N042(0)='1' AND  A(13)='1' AND D( 3)='0' AND E(15)='0' )then
          cVar2S22S122P012N056P043nsss(0) <='1';
          else
          cVar2S22S122P012N056P043nsss(0) <='0';
          end if;
        if(cVar1S23S122N045N049P047N042(0)='1' AND  A(13)='0' AND B(13)='0' AND A( 6)='0' )then
          cVar2S23S122N012P032P007nsss(0) <='1';
          else
          cVar2S23S122N012P032P007nsss(0) <='0';
          end if;
        if(cVar1S24S122N045N049P047N042(0)='1' AND  A(13)='0' AND B(13)='1' AND D(11)='1' )then
          cVar2S24S122N012P032P057nsss(0) <='1';
          else
          cVar2S24S122N012P032P057nsss(0) <='0';
          end if;
        if(cVar1S26S122N045N049P047N064(0)='1' AND  D( 8)='1' )then
          cVar2S26S122P069nsss(0) <='1';
          else
          cVar2S26S122P069nsss(0) <='0';
          end if;
        if(cVar1S27S122N045N049P047N064(0)='1' AND  D( 8)='0' AND A(12)='0' AND A(15)='1' )then
          cVar2S27S122N069P014P008nsss(0) <='1';
          else
          cVar2S27S122N069P014P008nsss(0) <='0';
          end if;
        if(cVar1S2S123P042N051P050N039(0)='1' AND  A(17)='1' )then
          cVar2S2S123P004nsss(0) <='1';
          else
          cVar2S2S123P004nsss(0) <='0';
          end if;
        if(cVar1S3S123P042N051P050N039(0)='1' AND  A(17)='0' AND B( 7)='1' )then
          cVar2S3S123N004P025nsss(0) <='1';
          else
          cVar2S3S123N004P025nsss(0) <='0';
          end if;
        if(cVar1S4S123P042N051P050N039(0)='1' AND  A(17)='0' AND B( 7)='0' AND E( 3)='1' )then
          cVar2S4S123N004N025P058nsss(0) <='1';
          else
          cVar2S4S123N004N025P058nsss(0) <='0';
          end if;
        if(cVar1S6S123N042P049P024N004(0)='1' AND  A(16)='1' AND A(15)='0' )then
          cVar2S6S123P006P008nsss(0) <='1';
          else
          cVar2S6S123P006P008nsss(0) <='0';
          end if;
        if(cVar1S7S123N042P049P024N004(0)='1' AND  A(16)='0' AND A( 7)='1' )then
          cVar2S7S123N006P005nsss(0) <='1';
          else
          cVar2S7S123N006P005nsss(0) <='0';
          end if;
        if(cVar1S8S123N042P049P024N004(0)='1' AND  A(16)='0' AND A( 7)='0' AND B(16)='0' )then
          cVar2S8S123N006N005P026nsss(0) <='1';
          else
          cVar2S8S123N006N005P026nsss(0) <='0';
          end if;
        if(cVar1S9S123N042P049N024P026(0)='1' AND  A( 6)='1' )then
          cVar2S9S123P007nsss(0) <='1';
          else
          cVar2S9S123P007nsss(0) <='0';
          end if;
        if(cVar1S10S123N042P049N024P026(0)='1' AND  A( 6)='0' AND A( 4)='1' )then
          cVar2S10S123N007P011nsss(0) <='1';
          else
          cVar2S10S123N007P011nsss(0) <='0';
          end if;
        if(cVar1S11S123N042P049N024P026(0)='1' AND  A( 6)='0' AND A( 4)='0' AND A(15)='1' )then
          cVar2S11S123N007N011P008nsss(0) <='1';
          else
          cVar2S11S123N007N011P008nsss(0) <='0';
          end if;
        if(cVar1S12S123N042P049N024N026(0)='1' AND  B( 6)='1' )then
          cVar2S12S123P027nsss(0) <='1';
          else
          cVar2S12S123P027nsss(0) <='0';
          end if;
        if(cVar1S13S123N042P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='0' AND A( 1)='1' )then
          cVar2S13S123N027P047P017nsss(0) <='1';
          else
          cVar2S13S123N027P047P017nsss(0) <='0';
          end if;
        if(cVar1S14S123N042P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='1' AND B( 7)='1' )then
          cVar2S14S123N027P047P025nsss(0) <='1';
          else
          cVar2S14S123N027P047P025nsss(0) <='0';
          end if;
        if(cVar1S15S123N042N049P045P007(0)='1' AND  B(18)='1' )then
          cVar2S15S123P022nsss(0) <='1';
          else
          cVar2S15S123P022nsss(0) <='0';
          end if;
        if(cVar1S16S123N042N049P045P007(0)='1' AND  B(18)='0' AND A( 2)='0' )then
          cVar2S16S123N022P015nsss(0) <='1';
          else
          cVar2S16S123N022P015nsss(0) <='0';
          end if;
        if(cVar1S17S123N042N049P045N007(0)='1' AND  A(17)='1' AND A( 3)='0' AND B(18)='1' )then
          cVar2S17S123P004P013P022nsss(0) <='1';
          else
          cVar2S17S123P004P013P022nsss(0) <='0';
          end if;
        if(cVar1S18S123N042N049P045N007(0)='1' AND  A(17)='0' AND A(16)='1' )then
          cVar2S18S123N004P006nsss(0) <='1';
          else
          cVar2S18S123N004P006nsss(0) <='0';
          end if;
        if(cVar1S19S123N042N049P045N007(0)='1' AND  A(17)='0' AND A(16)='0' AND D(11)='1' )then
          cVar2S19S123N004N006P057nsss(0) <='1';
          else
          cVar2S19S123N004N006P057nsss(0) <='0';
          end if;
        if(cVar1S20S123N042N049N045P047(0)='1' AND  A( 5)='1' AND E( 5)='1' AND B( 6)='1' )then
          cVar2S20S123P009P050P027nsss(0) <='1';
          else
          cVar2S20S123P009P050P027nsss(0) <='0';
          end if;
        if(cVar1S21S123N042N049N045P047(0)='1' AND  A( 5)='1' AND E( 5)='0' AND A(15)='1' )then
          cVar2S21S123P009N050P008nsss(0) <='1';
          else
          cVar2S21S123P009N050P008nsss(0) <='0';
          end if;
        if(cVar1S22S123N042N049N045P047(0)='1' AND  B(16)='0' AND A(12)='0' AND A(13)='1' )then
          cVar2S22S123P026P014P012nsss(0) <='1';
          else
          cVar2S22S123P026P014P012nsss(0) <='0';
          end if;
        if(cVar1S2S124P042P050N021N051(0)='1' AND  B( 7)='1' )then
          cVar2S2S124P025nsss(0) <='1';
          else
          cVar2S2S124P025nsss(0) <='0';
          end if;
        if(cVar1S3S124P042P050N021N051(0)='1' AND  B( 7)='0' AND E( 3)='1' )then
          cVar2S3S124N025P058nsss(0) <='1';
          else
          cVar2S3S124N025P058nsss(0) <='0';
          end if;
        if(cVar1S4S124P042P050N021N051(0)='1' AND  B( 7)='0' AND E( 3)='0' AND B( 0)='1' )then
          cVar2S4S124N025N058P039nsss(0) <='1';
          else
          cVar2S4S124N025N058P039nsss(0) <='0';
          end if;
        if(cVar1S5S124N042P045P027P024(0)='1' AND  A(16)='1' )then
          cVar2S5S124P006nsss(0) <='1';
          else
          cVar2S5S124P006nsss(0) <='0';
          end if;
        if(cVar1S6S124N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S6S124N006P004nsss(0) <='1';
          else
          cVar2S6S124N006P004nsss(0) <='0';
          end if;
        if(cVar1S7S124N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S7S124N006N004P007nsss(0) <='1';
          else
          cVar2S7S124N006N004P007nsss(0) <='0';
          end if;
        if(cVar1S8S124N042P045P027N024(0)='1' AND  B( 7)='1' AND E(15)='1' )then
          cVar2S8S124P025P043nsss(0) <='1';
          else
          cVar2S8S124P025P043nsss(0) <='0';
          end if;
        if(cVar1S9S124N042P045P027N024(0)='1' AND  B( 7)='1' AND E(15)='0' AND E( 6)='1' )then
          cVar2S9S124P025N043P046nsss(0) <='1';
          else
          cVar2S9S124P025N043P046nsss(0) <='0';
          end if;
        if(cVar1S10S124N042P045P027N024(0)='1' AND  B( 7)='0' AND A( 9)='1' )then
          cVar2S10S124N025P001nsss(0) <='1';
          else
          cVar2S10S124N025P001nsss(0) <='0';
          end if;
        if(cVar1S11S124N042P045P027N024(0)='1' AND  B( 7)='0' AND A( 9)='0' AND B(18)='1' )then
          cVar2S11S124N025N001P022nsss(0) <='1';
          else
          cVar2S11S124N025N001P022nsss(0) <='0';
          end if;
        if(cVar1S12S124N042N045P049P024(0)='1' AND  A(17)='1' )then
          cVar2S12S124P004nsss(0) <='1';
          else
          cVar2S12S124P004nsss(0) <='0';
          end if;
        if(cVar1S13S124N042N045P049P024(0)='1' AND  A(17)='0' AND A(16)='1' AND A(15)='0' )then
          cVar2S13S124N004P006P008nsss(0) <='1';
          else
          cVar2S13S124N004P006P008nsss(0) <='0';
          end if;
        if(cVar1S14S124N042N045P049P024(0)='1' AND  A(17)='0' AND A(16)='0' AND B(16)='0' )then
          cVar2S14S124N004N006P026nsss(0) <='1';
          else
          cVar2S14S124N004N006P026nsss(0) <='0';
          end if;
        if(cVar1S15S124N042N045P049N024(0)='1' AND  B(16)='1' )then
          cVar2S15S124P026nsss(0) <='1';
          else
          cVar2S15S124P026nsss(0) <='0';
          end if;
        if(cVar1S16S124N042N045P049N024(0)='1' AND  B(16)='0' AND B( 6)='1' )then
          cVar2S16S124N026P027nsss(0) <='1';
          else
          cVar2S16S124N026P027nsss(0) <='0';
          end if;
        if(cVar1S17S124N042N045P049N024(0)='1' AND  B(16)='0' AND B( 6)='0' AND E(14)='0' )then
          cVar2S17S124N026N027P047nsss(0) <='1';
          else
          cVar2S17S124N026N027P047nsss(0) <='0';
          end if;
        if(cVar1S18S124N042N045N049P047(0)='1' AND  A( 0)='1' AND E( 6)='0' )then
          cVar2S18S124P019P046nsss(0) <='1';
          else
          cVar2S18S124P019P046nsss(0) <='0';
          end if;
        if(cVar1S19S124N042N045N049P047(0)='1' AND  A( 0)='1' AND E( 6)='1' AND D( 1)='1' )then
          cVar2S19S124P019P046P064nsss(0) <='1';
          else
          cVar2S19S124P019P046P064nsss(0) <='0';
          end if;
        if(cVar1S20S124N042N045N049P047(0)='1' AND  A( 0)='0' AND A(11)='1' AND B( 9)='0' )then
          cVar2S20S124N019P016P021nsss(0) <='1';
          else
          cVar2S20S124N019P016P021nsss(0) <='0';
          end if;
        if(cVar1S21S124N042N045N049P047(0)='1' AND  A( 0)='0' AND A(11)='0' )then
          cVar2S21S124N019N016psss(0) <='1';
          else
          cVar2S21S124N019N016psss(0) <='0';
          end if;
        if(cVar1S22S124N042N045N049P047(0)='1' AND  B(16)='0' AND A(12)='0' AND E( 1)='1' )then
          cVar2S22S124P026P014P066nsss(0) <='1';
          else
          cVar2S22S124P026P014P066nsss(0) <='0';
          end if;
        if(cVar1S1S125N042P045P027P024(0)='1' AND  A(16)='1' )then
          cVar2S1S125P006nsss(0) <='1';
          else
          cVar2S1S125P006nsss(0) <='0';
          end if;
        if(cVar1S2S125N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S2S125N006P004nsss(0) <='1';
          else
          cVar2S2S125N006P004nsss(0) <='0';
          end if;
        if(cVar1S3S125N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S3S125N006N004P007nsss(0) <='1';
          else
          cVar2S3S125N006N004P007nsss(0) <='0';
          end if;
        if(cVar1S5S125N042N045P049P024(0)='1' AND  A(17)='1' )then
          cVar2S5S125P004nsss(0) <='1';
          else
          cVar2S5S125P004nsss(0) <='0';
          end if;
        if(cVar1S6S125N042N045P049P024(0)='1' AND  A(17)='0' AND A(16)='1' AND A(15)='0' )then
          cVar2S6S125N004P006P008nsss(0) <='1';
          else
          cVar2S6S125N004P006P008nsss(0) <='0';
          end if;
        if(cVar1S7S125N042N045P049P024(0)='1' AND  A(17)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S7S125N004N006P005nsss(0) <='1';
          else
          cVar2S7S125N004N006P005nsss(0) <='0';
          end if;
        if(cVar1S8S125N042N045P049N024(0)='1' AND  B(16)='1' )then
          cVar2S8S125P026nsss(0) <='1';
          else
          cVar2S8S125P026nsss(0) <='0';
          end if;
        if(cVar1S9S125N042N045P049N024(0)='1' AND  B(16)='0' AND B( 6)='1' )then
          cVar2S9S125N026P027nsss(0) <='1';
          else
          cVar2S9S125N026P027nsss(0) <='0';
          end if;
        if(cVar1S10S125N042N045N049P032(0)='1' AND  B(14)='0' AND D(11)='1' )then
          cVar2S10S125P030P057nsss(0) <='1';
          else
          cVar2S10S125P030P057nsss(0) <='0';
          end if;
        if(cVar1S11S125N042N045N049P032(0)='1' AND  B(14)='0' AND D(11)='0' AND D( 3)='0' )then
          cVar2S11S125P030N057P056nsss(0) <='1';
          else
          cVar2S11S125P030N057P056nsss(0) <='0';
          end if;
        if(cVar1S12S125N042N045N049N032(0)='1' AND  E(11)='0' AND B(10)='1' AND B( 9)='1' )then
          cVar2S12S125P059P038P021nsss(0) <='1';
          else
          cVar2S12S125P059P038P021nsss(0) <='0';
          end if;
        if(cVar1S13S125N042N045N049N032(0)='1' AND  E(11)='0' AND B(10)='0' AND B(15)='1' )then
          cVar2S13S125P059N038P028nsss(0) <='1';
          else
          cVar2S13S125P059N038P028nsss(0) <='0';
          end if;
        if(cVar1S2S126P042N051P023N005(0)='1' AND  A(17)='1' )then
          cVar2S2S126P004nsss(0) <='1';
          else
          cVar2S2S126P004nsss(0) <='0';
          end if;
        if(cVar1S3S126P042N051P023N005(0)='1' AND  A(17)='0' AND A( 6)='1' )then
          cVar2S3S126N004P007nsss(0) <='1';
          else
          cVar2S3S126N004P007nsss(0) <='0';
          end if;
        if(cVar1S4S126P042N051P023N005(0)='1' AND  A(17)='0' AND A( 6)='0' AND A(16)='1' )then
          cVar2S4S126N004N007P006nsss(0) <='1';
          else
          cVar2S4S126N004N007P006nsss(0) <='0';
          end if;
        if(cVar1S6S126P042N051N023N000(0)='1' AND  E( 5)='0' AND B( 0)='1' )then
          cVar2S6S126P050P039nsss(0) <='1';
          else
          cVar2S6S126P050P039nsss(0) <='0';
          end if;
        if(cVar1S7S126P042N051N023N000(0)='1' AND  E( 5)='0' AND B( 0)='0' AND B( 9)='1' )then
          cVar2S7S126P050N039P021nsss(0) <='1';
          else
          cVar2S7S126P050N039P021nsss(0) <='0';
          end if;
        if(cVar1S8S126N042P045P027P024(0)='1' AND  A(16)='1' )then
          cVar2S8S126P006nsss(0) <='1';
          else
          cVar2S8S126P006nsss(0) <='0';
          end if;
        if(cVar1S9S126N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S9S126N006P004nsss(0) <='1';
          else
          cVar2S9S126N006P004nsss(0) <='0';
          end if;
        if(cVar1S10S126N042P045P027P024(0)='1' AND  A(16)='0' AND A(17)='0' AND E(14)='1' )then
          cVar2S10S126N006N004P047nsss(0) <='1';
          else
          cVar2S10S126N006N004P047nsss(0) <='0';
          end if;
        if(cVar1S11S126N042P045P027N024(0)='1' AND  B( 7)='1' AND E(15)='1' )then
          cVar2S11S126P025P043nsss(0) <='1';
          else
          cVar2S11S126P025P043nsss(0) <='0';
          end if;
        if(cVar1S12S126N042P045P027N024(0)='1' AND  B( 7)='1' AND E(15)='0' AND E( 6)='1' )then
          cVar2S12S126P025N043P046nsss(0) <='1';
          else
          cVar2S12S126P025N043P046nsss(0) <='0';
          end if;
        if(cVar1S13S126N042P045P027N024(0)='1' AND  B( 7)='0' AND B(11)='1' )then
          cVar2S13S126N025P036nsss(0) <='1';
          else
          cVar2S13S126N025P036nsss(0) <='0';
          end if;
        if(cVar1S14S126N042P045P027N024(0)='1' AND  B( 7)='0' AND B(11)='0' AND D(10)='1' )then
          cVar2S14S126N025N036P061nsss(0) <='1';
          else
          cVar2S14S126N025N036P061nsss(0) <='0';
          end if;
        if(cVar1S15S126N042N045P049P007(0)='1' AND  A(16)='0' AND A( 0)='0' )then
          cVar2S15S126P006P019nsss(0) <='1';
          else
          cVar2S15S126P006P019nsss(0) <='0';
          end if;
        if(cVar1S16S126N042N045P049N007(0)='1' AND  A( 5)='1' AND E(13)='0' )then
          cVar2S16S126P009P051nsss(0) <='1';
          else
          cVar2S16S126P009P051nsss(0) <='0';
          end if;
        if(cVar1S17S126N042N045P049N007(0)='1' AND  A( 5)='1' AND E(13)='1' AND E(14)='0' )then
          cVar2S17S126P009P051P047nsss(0) <='1';
          else
          cVar2S17S126P009P051P047nsss(0) <='0';
          end if;
        if(cVar1S18S126N042N045P049N007(0)='1' AND  A( 5)='0' AND A(16)='1' AND A(12)='0' )then
          cVar2S18S126N009P006P014nsss(0) <='1';
          else
          cVar2S18S126N009P006P014nsss(0) <='0';
          end if;
        if(cVar1S19S126N042N045P049N007(0)='1' AND  A( 5)='0' AND A(16)='0' AND A( 7)='1' )then
          cVar2S19S126N009N006P005nsss(0) <='1';
          else
          cVar2S19S126N009N006P005nsss(0) <='0';
          end if;
        if(cVar1S20S126N042N045N049P059(0)='1' AND  E(15)='0' )then
          cVar2S20S126P043nsss(0) <='1';
          else
          cVar2S20S126P043nsss(0) <='0';
          end if;
        if(cVar1S21S126N042N045N049P059(0)='1' AND  E(15)='1' AND A( 8)='1' )then
          cVar2S21S126P043P003nsss(0) <='1';
          else
          cVar2S21S126P043P003nsss(0) <='0';
          end if;
        if(cVar1S22S126N042N045N049P059(0)='1' AND  E(15)='1' AND A( 8)='0' AND E( 9)='1' )then
          cVar2S22S126P043N003P067nsss(0) <='1';
          else
          cVar2S22S126P043N003P067nsss(0) <='0';
          end if;
        if(cVar1S23S126N042N045N049P059(0)='1' AND  E(15)='1' )then
          cVar2S23S126P043nsss(0) <='1';
          else
          cVar2S23S126P043nsss(0) <='0';
          end if;
        if(cVar1S24S126N042N045N049P059(0)='1' AND  E(15)='0' AND E( 9)='1' )then
          cVar2S24S126N043P067nsss(0) <='1';
          else
          cVar2S24S126N043P067nsss(0) <='0';
          end if;
        if(cVar1S1S127P042P050P004N040(0)='1' AND  D( 6)='1' )then
          cVar2S1S127P044nsss(0) <='1';
          else
          cVar2S1S127P044nsss(0) <='0';
          end if;
        if(cVar1S3S127P042P050N004N005(0)='1' AND  D(12)='1' )then
          cVar2S3S127P053nsss(0) <='1';
          else
          cVar2S3S127P053nsss(0) <='0';
          end if;
        if(cVar1S4S127P042P050N004N005(0)='1' AND  D(12)='0' AND A(18)='1' )then
          cVar2S4S127N053P002nsss(0) <='1';
          else
          cVar2S4S127N053P002nsss(0) <='0';
          end if;
        if(cVar1S5S127P042P050N004N005(0)='1' AND  D(12)='0' AND A(18)='0' AND E( 3)='1' )then
          cVar2S5S127N053N002P058nsss(0) <='1';
          else
          cVar2S5S127N053N002P058nsss(0) <='0';
          end if;
        if(cVar1S7S127N042P049P024N004(0)='1' AND  A(16)='1' AND A(12)='0' )then
          cVar2S7S127P006P014nsss(0) <='1';
          else
          cVar2S7S127P006P014nsss(0) <='0';
          end if;
        if(cVar1S8S127N042P049P024N004(0)='1' AND  A(16)='0' AND A( 7)='1' )then
          cVar2S8S127N006P005nsss(0) <='1';
          else
          cVar2S8S127N006P005nsss(0) <='0';
          end if;
        if(cVar1S9S127N042P049P024N004(0)='1' AND  A(16)='0' AND A( 7)='0' AND B(16)='0' )then
          cVar2S9S127N006N005P026nsss(0) <='1';
          else
          cVar2S9S127N006N005P026nsss(0) <='0';
          end if;
        if(cVar1S10S127N042P049N024P026(0)='1' AND  A( 6)='1' )then
          cVar2S10S127P007nsss(0) <='1';
          else
          cVar2S10S127P007nsss(0) <='0';
          end if;
        if(cVar1S11S127N042P049N024P026(0)='1' AND  A( 6)='0' AND A( 4)='1' )then
          cVar2S11S127N007P011nsss(0) <='1';
          else
          cVar2S11S127N007P011nsss(0) <='0';
          end if;
        if(cVar1S12S127N042P049N024P026(0)='1' AND  A( 6)='0' AND A( 4)='0' AND A(15)='1' )then
          cVar2S12S127N007N011P008nsss(0) <='1';
          else
          cVar2S12S127N007N011P008nsss(0) <='0';
          end if;
        if(cVar1S13S127N042P049N024N026(0)='1' AND  B( 6)='1' )then
          cVar2S13S127P027nsss(0) <='1';
          else
          cVar2S13S127P027nsss(0) <='0';
          end if;
        if(cVar1S14S127N042P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='0' AND E(15)='1' )then
          cVar2S14S127N027P047P043nsss(0) <='1';
          else
          cVar2S14S127N027P047P043nsss(0) <='0';
          end if;
        if(cVar1S15S127N042P049N024N026(0)='1' AND  B( 6)='0' AND E(14)='1' AND B( 7)='1' )then
          cVar2S15S127N027P047P025nsss(0) <='1';
          else
          cVar2S15S127N027P047P025nsss(0) <='0';
          end if;
        if(cVar1S16S127N042N049P045P024(0)='1' AND  A(16)='1' )then
          cVar2S16S127P006nsss(0) <='1';
          else
          cVar2S16S127P006nsss(0) <='0';
          end if;
        if(cVar1S17S127N042N049P045P024(0)='1' AND  A(16)='0' AND A(17)='1' )then
          cVar2S17S127N006P004nsss(0) <='1';
          else
          cVar2S17S127N006P004nsss(0) <='0';
          end if;
        if(cVar1S18S127N042N049P045P024(0)='1' AND  A(16)='0' AND A(17)='0' AND A( 6)='1' )then
          cVar2S18S127N006N004P007nsss(0) <='1';
          else
          cVar2S18S127N006N004P007nsss(0) <='0';
          end if;
        if(cVar1S19S127N042N049P045N024(0)='1' AND  B( 7)='1' AND E(15)='1' )then
          cVar2S19S127P025P043nsss(0) <='1';
          else
          cVar2S19S127P025P043nsss(0) <='0';
          end if;
        if(cVar1S20S127N042N049P045N024(0)='1' AND  B( 7)='1' AND E(15)='0' AND E( 6)='1' )then
          cVar2S20S127P025N043P046nsss(0) <='1';
          else
          cVar2S20S127P025N043P046nsss(0) <='0';
          end if;
        if(cVar1S21S127N042N049P045N024(0)='1' AND  B( 7)='0' AND A( 4)='1' )then
          cVar2S21S127N025P011nsss(0) <='1';
          else
          cVar2S21S127N025P011nsss(0) <='0';
          end if;
        if(cVar1S22S127N042N049P045N024(0)='1' AND  B( 7)='0' AND A( 4)='0' AND A( 3)='0' )then
          cVar2S22S127N025N011P013nsss(0) <='1';
          else
          cVar2S22S127N025N011P013nsss(0) <='0';
          end if;
        if(cVar1S23S127N042N049N045P020(0)='1' AND  A( 8)='1' )then
          cVar2S23S127P003nsss(0) <='1';
          else
          cVar2S23S127P003nsss(0) <='0';
          end if;
        if(cVar1S24S127N042N049N045P020(0)='1' AND  A( 8)='0' AND D( 5)='1' )then
          cVar2S24S127N003P048nsss(0) <='1';
          else
          cVar2S24S127N003P048nsss(0) <='0';
          end if;
        if(cVar1S25S127N042N049N045P020(0)='1' AND  A( 8)='0' AND D( 5)='0' AND A(18)='1' )then
          cVar2S25S127N003N048P002nsss(0) <='1';
          else
          cVar2S25S127N003N048P002nsss(0) <='0';
          end if;
        if(cVar1S26S127N042N049N045N020(0)='1' AND  B( 0)='0' AND E(14)='0' AND B(12)='1' )then
          cVar2S26S127P039P047P034nsss(0) <='1';
          else
          cVar2S26S127P039P047P034nsss(0) <='0';
          end if;
        if(cVar1S27S127N042N049N045N020(0)='1' AND  B( 0)='1' AND B( 9)='1' )then
          cVar2S27S127P039P021nsss(0) <='1';
          else
          cVar2S27S127P039P021nsss(0) <='0';
          end if;
        if(cVar1S28S127N042N049N045N020(0)='1' AND  B( 0)='1' AND B( 9)='0' AND A(11)='1' )then
          cVar2S28S127P039N021P016nsss(0) <='1';
          else
          cVar2S28S127P039N021P016nsss(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV3 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar1S0S0P055P030nsss(0)='1'  OR cVar1S1S0P055N030P031nsss(0)='1'  OR cVar1S2S0P055N030N031P028nsss(0)='1'  OR cVar2S3S0P029nsss(0)='1'  )then
          oVar1S0(0) <='1';
          else
          oVar1S0(0) <='0';
          end if;
        if(cVar2S4S0N029P061nsss(0)='1'  OR cVar2S5S0N029N061P049nsss(0)='1'  OR cVar1S6S0N055P059P061P032nsss(0)='1'  OR cVar2S7S0P060nsss(0)='1'  )then
          oVar1S1(0) <='1';
          else
          oVar1S1(0) <='0';
          end if;
        if(cVar2S8S0N060P033nsss(0)='1'  OR cVar2S9S0N060N033P034nsss(0)='1'  OR cVar1S10S0N055P059N061P058nsss(0)='1'  OR cVar2S11S0P063nsss(0)='1'  )then
          oVar1S2(0) <='1';
          else
          oVar1S2(0) <='0';
          end if;
        if(cVar2S12S0N063P030nsss(0)='1'  OR cVar2S13S0N063N030P067nsss(0)='1'  OR cVar1S14S0N055N059P052P029nsss(0)='1'  OR cVar2S15S0P027nsss(0)='1'  )then
          oVar1S3(0) <='1';
          else
          oVar1S3(0) <='0';
          end if;
        if(cVar2S16S0N027P051nsss(0)='1'  OR cVar2S17S0N027N051P028nsss(0)='1'  OR cVar2S18S0P049nsss(0)='1'  OR cVar2S19S0N049P024nsss(0)='1'  )then
          oVar1S4(0) <='1';
          else
          oVar1S4(0) <='0';
          end if;
        if(cVar2S20S0N049N024P025nsss(0)='1'  OR cVar2S21S0P065P063nsss(0)='1'  OR cVar2S22S0N065P043nsss(0)='1'  OR cVar2S23S0N065N043P067nsss(0)='1'  )then
          oVar1S5(0) <='1';
          else
          oVar1S5(0) <='0';
          end if;
        if(cVar1S0S1P058P033P060nsss(0)='1'  OR cVar2S1S1P056nsss(0)='1'  OR cVar2S2S1N056P059nsss(0)='1'  OR cVar1S3S1P058N033P031nsss(0)='1'  )then
          oVar1S7(0) <='1';
          else
          oVar1S7(0) <='0';
          end if;
        if(cVar1S4S1P058N033N031P032nsss(0)='1'  OR cVar2S5S1P030nsss(0)='1'  OR cVar2S6S1N030P035nsss(0)='1'  OR cVar2S7S1N030N035P053nsss(0)='1'  )then
          oVar1S8(0) <='1';
          else
          oVar1S8(0) <='0';
          end if;
        if(cVar1S8S1N058P051P053P028nsss(0)='1'  OR cVar2S9S1P026nsss(0)='1'  OR cVar2S10S1N026P029nsss(0)='1'  OR cVar2S11S1N026N029P027nsss(0)='1'  )then
          oVar1S9(0) <='1';
          else
          oVar1S9(0) <='0';
          end if;
        if(cVar1S12S1N058P051N053P026nsss(0)='1'  OR cVar2S13S1P027nsss(0)='1'  OR cVar2S14S1N027P054nsss(0)='1'  OR cVar2S15S1N027N054P032nsss(0)='1'  )then
          oVar1S10(0) <='1';
          else
          oVar1S10(0) <='0';
          end if;
        if(cVar1S16S1N058N051P046P025nsss(0)='1'  OR cVar2S17S1P027nsss(0)='1'  OR cVar2S18S1N027P024nsss(0)='1'  OR cVar2S19S1N027N024P026nsss(0)='1'  )then
          oVar1S11(0) <='1';
          else
          oVar1S11(0) <='0';
          end if;
        if(cVar2S20S1P035P062nsss(0)='1'  OR cVar2S21S1N035P037nsss(0)='1'  OR cVar2S22S1N035N037P034nsss(0)='1'  OR cVar2S23S1P054P056nsss(0)='1'  )then
          oVar1S12(0) <='1';
          else
          oVar1S12(0) <='0';
          end if;
        if(cVar2S24S1P054N056P029nsss(0)='1'  OR cVar2S25S1N054P042nsss(0)='1'  OR cVar2S26S1N054N042P039nsss(0)='1'  )then
          oVar1S13(0) <='1';
          else
          oVar1S13(0) <='0';
          end if;
        if(cVar1S0S2P068P019P015P066nsss(0)='1'  OR cVar2S1S2P013P067nsss(0)='1'  OR cVar2S2S2P066nsss(0)='1'  OR cVar2S3S2N066P016nsss(0)='1'  )then
          oVar1S14(0) <='1';
          else
          oVar1S14(0) <='0';
          end if;
        if(cVar2S4S2P062nsss(0)='1'  OR cVar1S5S2P068N019P011P018nsss(0)='1'  OR cVar2S6S2P017nsss(0)='1'  OR cVar2S7S2N017P067P064nsss(0)='1'  )then
          oVar1S15(0) <='1';
          else
          oVar1S15(0) <='0';
          end if;
        if(cVar2S8S2P065P052nsss(0)='1'  OR cVar2S9S2P065N052P017nsss(0)='1'  OR cVar2S10S2P037P018nsss(0)='1'  OR cVar1S11S2N068P040P038nsss(0)='1'  )then
          oVar1S16(0) <='1';
          else
          oVar1S16(0) <='0';
          end if;
        if(cVar1S12S2N068P040N038P023nsss(0)='1'  OR cVar2S13S2P021nsss(0)='1'  OR cVar2S14S2N021P004nsss(0)='1'  OR cVar2S15S2N021N004P046nsss(0)='1'  )then
          oVar1S17(0) <='1';
          else
          oVar1S17(0) <='0';
          end if;
        if(cVar1S16S2N068N040P050P027nsss(0)='1'  OR cVar2S17S2P052nsss(0)='1'  OR cVar2S18S2N052P026nsss(0)='1'  OR cVar2S19S2N052N026P051nsss(0)='1'  )then
          oVar1S18(0) <='1';
          else
          oVar1S18(0) <='0';
          end if;
        if(cVar2S20S2P025nsss(0)='1'  OR cVar2S21S2N025P036nsss(0)='1'  OR cVar2S22S2P060P033nsss(0)='1'  OR cVar2S23S2P060N033P067nsss(0)='1'  )then
          oVar1S19(0) <='1';
          else
          oVar1S19(0) <='0';
          end if;
        if(cVar2S24S2N060psss(0)='1'  )then
          oVar1S20(0) <='1';
          else
          oVar1S20(0) <='0';
          end if;
        if(cVar2S0S3P013nsss(0)='1'  OR cVar2S1S3P013P037nsss(0)='1'  OR cVar2S2S3P013N037P016nsss(0)='1'  OR cVar2S3S3P066P018nsss(0)='1'  )then
          oVar1S21(0) <='1';
          else
          oVar1S21(0) <='0';
          end if;
        if(cVar2S4S3P066P018P014nsss(0)='1'  OR cVar2S5S3N066P016nsss(0)='1'  OR cVar2S6S3P066P056nsss(0)='1'  OR cVar2S7S3N066P014P018nsss(0)='1'  )then
          oVar1S22(0) <='1';
          else
          oVar1S22(0) <='0';
          end if;
        if(cVar2S8S3P009P017nsss(0)='1'  OR cVar2S9S3P015P066nsss(0)='1'  OR cVar2S10S3P015N066P014nsss(0)='1'  OR cVar2S11S3P015P016nsss(0)='1'  )then
          oVar1S23(0) <='1';
          else
          oVar1S23(0) <='0';
          end if;
        if(cVar2S12S3P015P016P013nsss(0)='1'  OR cVar2S13S3P017P037P013nsss(0)='1'  OR cVar2S14S3P017N037P035nsss(0)='1'  OR cVar2S15S3N017P016P014nsss(0)='1'  )then
          oVar1S24(0) <='1';
          else
          oVar1S24(0) <='0';
          end if;
        if(cVar2S16S3N017N016P037nsss(0)='1'  OR cVar2S17S3P036P055nsss(0)='1'  OR cVar2S18S3P036N055P017nsss(0)='1'  OR cVar1S19S3N068P040P021nsss(0)='1'  )then
          oVar1S25(0) <='1';
          else
          oVar1S25(0) <='0';
          end if;
        if(cVar1S20S3N068P040N021P020nsss(0)='1'  OR cVar2S21S3P023nsss(0)='1'  OR cVar2S22S3N023P022nsss(0)='1'  OR cVar2S23S3N023N022P046nsss(0)='1'  )then
          oVar1S26(0) <='1';
          else
          oVar1S26(0) <='0';
          end if;
        if(cVar1S24S3N068N040P050nsss(0)='1'  OR cVar1S25S3N068N040N050P046nsss(0)='1'  OR cVar2S26S3P060nsss(0)='1'  OR cVar2S27S3N060P051P053nsss(0)='1'  )then
          oVar1S27(0) <='1';
          else
          oVar1S27(0) <='0';
          end if;
        if(cVar2S28S3N060N051P057nsss(0)='1'  )then
          oVar1S28(0) <='1';
          else
          oVar1S28(0) <='0';
          end if;
        if(cVar1S0S4P040P038nsss(0)='1'  OR cVar1S1S4P040N038P067P023nsss(0)='1'  OR cVar2S2S4P068nsss(0)='1'  OR cVar1S3S4N040P044P023nsss(0)='1'  )then
          oVar1S29(0) <='1';
          else
          oVar1S29(0) <='0';
          end if;
        if(cVar1S4S4N040P044N023P022nsss(0)='1'  OR cVar2S5S4P025nsss(0)='1'  OR cVar2S6S4N025P024nsss(0)='1'  OR cVar2S7S4N025N024P050nsss(0)='1'  )then
          oVar1S30(0) <='1';
          else
          oVar1S30(0) <='0';
          end if;
        if(cVar1S8S4N040N044P047P024nsss(0)='1'  OR cVar2S9S4P026nsss(0)='1'  OR cVar2S10S4N026P025nsss(0)='1'  OR cVar2S11S4N026N025P027nsss(0)='1'  )then
          oVar1S31(0) <='1';
          else
          oVar1S31(0) <='0';
          end if;
        if(cVar2S12S4P059P058nsss(0)='1'  OR cVar2S13S4P059P058P012nsss(0)='1'  OR cVar2S14S4N059P063P065nsss(0)='1'  OR cVar2S15S4N059N063P054nsss(0)='1'  )then
          oVar1S32(0) <='1';
          else
          oVar1S32(0) <='0';
          end if;
        if(cVar2S16S4P056P031nsss(0)='1'  OR cVar2S17S4P056N031P029nsss(0)='1'  OR cVar2S18S4N056psss(0)='1'  )then
          oVar1S33(0) <='1';
          else
          oVar1S33(0) <='0';
          end if;
        if(cVar1S0S5P044P023nsss(0)='1'  OR cVar1S1S5P044N023P022nsss(0)='1'  OR cVar1S2S5P044N023N022P025nsss(0)='1'  OR cVar2S3S5P024nsss(0)='1'  )then
          oVar1S34(0) <='1';
          else
          oVar1S34(0) <='0';
          end if;
        if(cVar2S4S5N024P054nsss(0)='1'  OR cVar1S5S5N044P040P021nsss(0)='1'  OR cVar1S6S5N044P040N021P020nsss(0)='1'  OR cVar2S7S5P023nsss(0)='1'  )then
          oVar1S35(0) <='1';
          else
          oVar1S35(0) <='0';
          end if;
        if(cVar2S8S5N023P000nsss(0)='1'  OR cVar2S9S5N023N000P015nsss(0)='1'  OR cVar1S10S5N044N040P047P006nsss(0)='1'  OR cVar2S11S5P066nsss(0)='1'  )then
          oVar1S36(0) <='1';
          else
          oVar1S36(0) <='0';
          end if;
        if(cVar2S12S5P066P064P067nsss(0)='1'  OR cVar2S13S5P031P013nsss(0)='1'  OR cVar2S14S5P031N013P055nsss(0)='1'  OR cVar2S15S5N031P030nsss(0)='1'  )then
          oVar1S37(0) <='1';
          else
          oVar1S37(0) <='0';
          end if;
        if(cVar2S16S5N031N030P029nsss(0)='1'  OR cVar2S17S5P061P032P058nsss(0)='1'  OR cVar2S18S5P061N032P059nsss(0)='1'  OR cVar2S19S5N061P041nsss(0)='1'  )then
          oVar1S38(0) <='1';
          else
          oVar1S38(0) <='0';
          end if;
        if(cVar2S20S5N061N041P045nsss(0)='1'  )then
          oVar1S39(0) <='1';
          else
          oVar1S39(0) <='0';
          end if;
        if(cVar1S0S6P044P023nsss(0)='1'  OR cVar1S1S6P044N023P004nsss(0)='1'  OR cVar1S2S6P044N023N004P006nsss(0)='1'  OR cVar2S3S6P007P025nsss(0)='1'  )then
          oVar1S40(0) <='1';
          else
          oVar1S40(0) <='0';
          end if;
        if(cVar2S4S6N007P014nsss(0)='1'  OR cVar1S5S6N044P015P050P027nsss(0)='1'  OR cVar2S6S6P026nsss(0)='1'  OR cVar2S7S6N026P029P048nsss(0)='1'  )then
          oVar1S41(0) <='1';
          else
          oVar1S41(0) <='0';
          end if;
        if(cVar2S8S6N026N029P010nsss(0)='1'  OR cVar2S9S6P031P009nsss(0)='1'  OR cVar2S10S6N031P013nsss(0)='1'  OR cVar2S11S6N031P013P029nsss(0)='1'  )then
          oVar1S42(0) <='1';
          else
          oVar1S42(0) <='0';
          end if;
        if(cVar2S12S6P040nsss(0)='1'  OR cVar2S13S6N040P042nsss(0)='1'  OR cVar2S14S6P012P037nsss(0)='1'  OR cVar2S15S6P012P037P014nsss(0)='1'  )then
          oVar1S43(0) <='1';
          else
          oVar1S43(0) <='0';
          end if;
        if(cVar2S16S6P012P063P017nsss(0)='1'  OR cVar2S17S6P058P012nsss(0)='1'  OR cVar2S18S6N058P037P033nsss(0)='1'  OR cVar2S19S6P033P017nsss(0)='1'  )then
          oVar1S44(0) <='1';
          else
          oVar1S44(0) <='0';
          end if;
        if(cVar2S20S6P033P017P016nsss(0)='1'  OR cVar2S21S6P061P059nsss(0)='1'  OR cVar2S22S6P061N059P018nsss(0)='1'  OR cVar2S23S6N061P040nsss(0)='1'  )then
          oVar1S45(0) <='1';
          else
          oVar1S45(0) <='0';
          end if;
        if(cVar2S24S6N061N040P065nsss(0)='1'  )then
          oVar1S46(0) <='1';
          else
          oVar1S46(0) <='0';
          end if;
        if(cVar1S0S7P050P027P048nsss(0)='1'  OR cVar1S1S7P050P027N048P009nsss(0)='1'  OR cVar2S2S7P008nsss(0)='1'  OR cVar2S3S7N008P011nsss(0)='1'  )then
          oVar1S47(0) <='1';
          else
          oVar1S47(0) <='0';
          end if;
        if(cVar1S4S7P050N027P052P008nsss(0)='1'  OR cVar2S5S7P029nsss(0)='1'  OR cVar2S6S7N029P010nsss(0)='1'  OR cVar2S7S7N029N010P006nsss(0)='1'  )then
          oVar1S48(0) <='1';
          else
          oVar1S48(0) <='0';
          end if;
        if(cVar2S8S7P026nsss(0)='1'  OR cVar2S9S7N026P015nsss(0)='1'  OR cVar2S10S7P057nsss(0)='1'  OR cVar1S11S7N050P044P023nsss(0)='1'  )then
          oVar1S49(0) <='1';
          else
          oVar1S49(0) <='0';
          end if;
        if(cVar1S12S7N050P044N023P004nsss(0)='1'  OR cVar2S13S7P006nsss(0)='1'  OR cVar2S14S7N006P007P025nsss(0)='1'  OR cVar2S15S7N006N007P002nsss(0)='1'  )then
          oVar1S50(0) <='1';
          else
          oVar1S50(0) <='0';
          end if;
        if(cVar2S16S7P013nsss(0)='1'  OR cVar2S17S7N013P067nsss(0)='1'  OR cVar2S18S7P067nsss(0)='1'  OR cVar2S19S7P067P065nsss(0)='1'  )then
          oVar1S51(0) <='1';
          else
          oVar1S51(0) <='0';
          end if;
        if(cVar2S20S7P021nsss(0)='1'  OR cVar2S21S7N021P020nsss(0)='1'  OR cVar2S22S7P062P067nsss(0)='1'  OR cVar2S23S7P062P067P065nsss(0)='1'  )then
          oVar1S52(0) <='1';
          else
          oVar1S52(0) <='0';
          end if;
        if(cVar2S24S7N062P066P068nsss(0)='1'  OR cVar2S25S7N062N066P047nsss(0)='1'  )then
          oVar1S53(0) <='1';
          else
          oVar1S53(0) <='0';
          end if;
        if(cVar1S0S8P044P023P005nsss(0)='1'  OR cVar1S1S8P044P023N005P004nsss(0)='1'  OR cVar2S2S8P015nsss(0)='1'  OR cVar1S3S8P044N023P004nsss(0)='1'  )then
          oVar1S54(0) <='1';
          else
          oVar1S54(0) <='0';
          end if;
        if(cVar1S4S8P044N023N004P006nsss(0)='1'  OR cVar2S5S8P007nsss(0)='1'  OR cVar2S6S8N007P042P046nsss(0)='1'  OR cVar2S7S8N007P042P002nsss(0)='1'  )then
          oVar1S55(0) <='1';
          else
          oVar1S55(0) <='0';
          end if;
        if(cVar1S8S8N044P050P027P009nsss(0)='1'  OR cVar2S9S8P048nsss(0)='1'  OR cVar2S10S8N048P006nsss(0)='1'  OR cVar2S11S8N048N006P008nsss(0)='1'  )then
          oVar1S56(0) <='1';
          else
          oVar1S56(0) <='0';
          end if;
        if(cVar2S12S8P008nsss(0)='1'  OR cVar2S13S8N008P010nsss(0)='1'  OR cVar2S14S8N008N010P006nsss(0)='1'  OR cVar2S15S8P029nsss(0)='1'  )then
          oVar1S57(0) <='1';
          else
          oVar1S57(0) <='0';
          end if;
        if(cVar2S16S8N029P009nsss(0)='1'  OR cVar2S17S8P028P054nsss(0)='1'  OR cVar2S18S8N028P008P026nsss(0)='1'  OR cVar2S19S8N028N008P009nsss(0)='1'  )then
          oVar1S58(0) <='1';
          else
          oVar1S58(0) <='0';
          end if;
        if(cVar2S20S8P022P043nsss(0)='1'  OR cVar2S21S8P022N043P039nsss(0)='1'  OR cVar2S22S8N022psss(0)='1'  OR cVar2S23S8P061P013nsss(0)='1'  )then
          oVar1S59(0) <='1';
          else
          oVar1S59(0) <='0';
          end if;
        if(cVar2S24S8P061P013P068nsss(0)='1'  OR cVar2S25S8N061P030nsss(0)='1'  OR cVar2S26S8P065P034nsss(0)='1'  OR cVar2S27S8P065N034P063nsss(0)='1'  )then
          oVar1S60(0) <='1';
          else
          oVar1S60(0) <='0';
          end if;
        if(cVar2S28S8N065P067P015nsss(0)='1'  )then
          oVar1S61(0) <='1';
          else
          oVar1S61(0) <='0';
          end if;
        if(cVar1S0S9P051P028P055nsss(0)='1'  OR cVar1S1S9P051P028P055P057nsss(0)='1'  OR cVar1S2S9P051N028P029nsss(0)='1'  OR cVar2S3S9P008P013nsss(0)='1'  )then
          oVar1S62(0) <='1';
          else
          oVar1S62(0) <='0';
          end if;
        if(cVar2S4S9N008P009nsss(0)='1'  OR cVar2S5S9N008N009P007nsss(0)='1'  OR cVar2S6S9P027P009nsss(0)='1'  OR cVar2S7S9N027P057P030nsss(0)='1'  )then
          oVar1S63(0) <='1';
          else
          oVar1S63(0) <='0';
          end if;
        if(cVar1S8S9N051P022P043P062nsss(0)='1'  OR cVar1S9S9N051P022N043P004nsss(0)='1'  OR cVar2S10S9P010P023nsss(0)='1'  OR cVar1S11S9N051N022P044P023nsss(0)='1'  )then
          oVar1S64(0) <='1';
          else
          oVar1S64(0) <='0';
          end if;
        if(cVar2S12S9P025P014nsss(0)='1'  OR cVar2S13S9N025P047nsss(0)='1'  OR cVar2S14S9N025N047P019nsss(0)='1'  OR cVar2S15S9P027nsss(0)='1'  )then
          oVar1S65(0) <='1';
          else
          oVar1S65(0) <='0';
          end if;
        if(cVar2S16S9N027P026nsss(0)='1'  OR cVar2S17S9N027N026P029nsss(0)='1'  OR cVar2S18S9P038P021nsss(0)='1'  OR cVar2S19S9P038N021P002nsss(0)='1'  )then
          oVar1S66(0) <='1';
          else
          oVar1S66(0) <='0';
          end if;
        if(cVar2S20S9N038P009P065nsss(0)='1'  OR cVar2S21S9N038P009P046nsss(0)='1'  )then
          oVar1S67(0) <='1';
          else
          oVar1S67(0) <='0';
          end if;
        if(cVar2S0S10P067P008nsss(0)='1'  OR cVar2S1S10P067N008P047nsss(0)='1'  OR cVar2S2S10P067P013nsss(0)='1'  OR cVar2S3S10P027nsss(0)='1'  )then
          oVar1S68(0) <='1';
          else
          oVar1S68(0) <='0';
          end if;
        if(cVar2S4S10N027P025nsss(0)='1'  OR cVar2S5S10N027N025P006nsss(0)='1'  OR cVar2S6S10P022P043nsss(0)='1'  OR cVar2S7S10P022N043P004nsss(0)='1'  )then
          oVar1S69(0) <='1';
          else
          oVar1S69(0) <='0';
          end if;
        if(cVar2S8S10N022psss(0)='1'  OR cVar2S9S10P066P018P010nsss(0)='1'  OR cVar2S10S10P066P018P033nsss(0)='1'  OR cVar2S11S10N066P069nsss(0)='1'  )then
          oVar1S70(0) <='1';
          else
          oVar1S70(0) <='0';
          end if;
        if(cVar2S12S10P068P066nsss(0)='1'  OR cVar2S13S10P068P065P014nsss(0)='1'  OR cVar2S14S10P068P067P015nsss(0)='1'  OR cVar2S15S10P016P012P034nsss(0)='1'  )then
          oVar1S71(0) <='1';
          else
          oVar1S71(0) <='0';
          end if;
        if(cVar2S16S10P003P035nsss(0)='1'  OR cVar2S17S10P003N035P037nsss(0)='1'  OR cVar2S18S10P066P067P015nsss(0)='1'  OR cVar2S19S10P016P018nsss(0)='1'  )then
          oVar1S72(0) <='1';
          else
          oVar1S72(0) <='0';
          end if;
        if(cVar2S20S10P016N018P037nsss(0)='1'  OR cVar2S21S10P016P068nsss(0)='1'  OR cVar2S22S10P003P035P067nsss(0)='1'  OR cVar2S23S10P067P051nsss(0)='1'  )then
          oVar1S73(0) <='1';
          else
          oVar1S73(0) <='0';
          end if;
        if(cVar2S24S10P067N051P043nsss(0)='1'  OR cVar2S25S10P067P069P011nsss(0)='1'  OR cVar2S26S10P034P066P019nsss(0)='1'  OR cVar2S27S10P066P012P008nsss(0)='1'  )then
          oVar1S74(0) <='1';
          else
          oVar1S74(0) <='0';
          end if;
        if(cVar2S28S10P066P012P018nsss(0)='1'  OR cVar2S29S10N066P069P016nsss(0)='1'  OR cVar2S30S10N066N069P008nsss(0)='1'  OR cVar2S31S10P034P063P012nsss(0)='1'  )then
          oVar1S75(0) <='1';
          else
          oVar1S75(0) <='0';
          end if;
        if(cVar2S32S10N034P031P013nsss(0)='1'  OR cVar2S33S10N034N031P038nsss(0)='1'  )then
          oVar1S76(0) <='1';
          else
          oVar1S76(0) <='0';
          end if;
        if(cVar1S0S11P048P025P007nsss(0)='1'  OR cVar1S1S11P048P025N007P006nsss(0)='1'  OR cVar2S2S11P009nsss(0)='1'  OR cVar2S3S11N009P005nsss(0)='1'  )then
          oVar1S77(0) <='1';
          else
          oVar1S77(0) <='0';
          end if;
        if(cVar2S4S11N009N005P008nsss(0)='1'  OR cVar2S5S11P009nsss(0)='1'  OR cVar2S6S11N009P007nsss(0)='1'  OR cVar2S7S11N009N007P008nsss(0)='1'  )then
          oVar1S78(0) <='1';
          else
          oVar1S78(0) <='0';
          end if;
        if(cVar2S8S11P046nsss(0)='1'  OR cVar2S9S11P006P024nsss(0)='1'  OR cVar2S10S11P006N024P026nsss(0)='1'  OR cVar2S11S11N006P026P008nsss(0)='1'  )then
          oVar1S79(0) <='1';
          else
          oVar1S79(0) <='0';
          end if;
        if(cVar2S12S11N006N026P058nsss(0)='1'  OR cVar1S13S11N048P051P028P055nsss(0)='1'  OR cVar1S14S11N048P051N028P029nsss(0)='1'  OR cVar2S15S11P026P008nsss(0)='1'  )then
          oVar1S80(0) <='1';
          else
          oVar1S80(0) <='0';
          end if;
        if(cVar2S16S11P026N008P047nsss(0)='1'  OR cVar2S17S11N026P027nsss(0)='1'  OR cVar2S18S11P035nsss(0)='1'  OR cVar2S19S11P044nsss(0)='1'  )then
          oVar1S81(0) <='1';
          else
          oVar1S81(0) <='0';
          end if;
        if(cVar2S20S11N044P040nsss(0)='1'  OR cVar2S21S11N044N040P014nsss(0)='1'  OR cVar2S22S11P042P008nsss(0)='1'  OR cVar2S23S11N042P043nsss(0)='1'  )then
          oVar1S82(0) <='1';
          else
          oVar1S82(0) <='0';
          end if;
        if(cVar2S24S11N042N043P064nsss(0)='1'  OR cVar2S25S11P043P007P031nsss(0)='1'  OR cVar2S26S11P043P007P047nsss(0)='1'  OR cVar2S27S11P043P024nsss(0)='1'  )then
          oVar1S83(0) <='1';
          else
          oVar1S83(0) <='0';
          end if;
        if(cVar2S28S11P043N024P025nsss(0)='1'  )then
          oVar1S84(0) <='1';
          else
          oVar1S84(0) <='0';
          end if;
        if(cVar1S0S12P048P025P007nsss(0)='1'  OR cVar1S1S12P048P025N007P006nsss(0)='1'  OR cVar2S2S12P009nsss(0)='1'  OR cVar2S3S12N009P005nsss(0)='1'  )then
          oVar1S85(0) <='1';
          else
          oVar1S85(0) <='0';
          end if;
        if(cVar2S4S12N009N005P008nsss(0)='1'  OR cVar1S5S12P048N025P027P052nsss(0)='1'  OR cVar2S6S12P024nsss(0)='1'  OR cVar2S7S12N024P026nsss(0)='1'  )then
          oVar1S86(0) <='1';
          else
          oVar1S86(0) <='0';
          end if;
        if(cVar2S8S12N024N026P008nsss(0)='1'  OR cVar2S9S12P008P026nsss(0)='1'  OR cVar2S10S12P008N026P028nsss(0)='1'  OR cVar2S11S12N008psss(0)='1'  )then
          oVar1S87(0) <='1';
          else
          oVar1S87(0) <='0';
          end if;
        if(cVar2S12S12P003P016nsss(0)='1'  OR cVar2S13S12P003P016P018nsss(0)='1'  OR cVar2S14S12P026nsss(0)='1'  OR cVar2S15S12P026P049nsss(0)='1'  )then
          oVar1S88(0) <='1';
          else
          oVar1S88(0) <='0';
          end if;
        if(cVar2S16S12P047P026nsss(0)='1'  OR cVar2S17S12P047N026P024nsss(0)='1'  OR cVar2S18S12N047P050P011nsss(0)='1'  OR cVar1S19S12N048P001P041nsss(0)='1'  )then
          oVar1S89(0) <='1';
          else
          oVar1S89(0) <='0';
          end if;
        if(cVar2S20S12P033P010nsss(0)='1'  OR cVar2S21S12P033N010P066nsss(0)='1'  OR cVar2S22S12P015P013P018nsss(0)='1'  )then
          oVar1S90(0) <='1';
          else
          oVar1S90(0) <='0';
          end if;
        if(cVar1S0S13P048P025P007nsss(0)='1'  OR cVar1S1S13P048P025N007P016nsss(0)='1'  OR cVar1S2S13P048N025P027P011nsss(0)='1'  OR cVar2S3S13P050nsss(0)='1'  )then
          oVar1S91(0) <='1';
          else
          oVar1S91(0) <='0';
          end if;
        if(cVar2S4S13P006P024nsss(0)='1'  OR cVar2S5S13P006N024P026nsss(0)='1'  OR cVar2S6S13N006P017P026nsss(0)='1'  OR cVar2S7S13N006P017P052nsss(0)='1'  )then
          oVar1S92(0) <='1';
          else
          oVar1S92(0) <='0';
          end if;
        if(cVar2S8S13P028nsss(0)='1'  OR cVar2S9S13N028P026nsss(0)='1'  OR cVar2S10S13P010P016P054nsss(0)='1'  OR cVar2S11S13P010P016psss(0)='1'  )then
          oVar1S93(0) <='1';
          else
          oVar1S93(0) <='0';
          end if;
        if(cVar2S12S13N010P011nsss(0)='1'  OR cVar2S13S13N010N011P009nsss(0)='1'  OR cVar2S14S13P029P011nsss(0)='1'  OR cVar2S15S13P029N011P009nsss(0)='1'  )then
          oVar1S94(0) <='1';
          else
          oVar1S94(0) <='0';
          end if;
        if(cVar2S16S13N029P009P011nsss(0)='1'  OR cVar1S17S13N048N051P038P021nsss(0)='1'  OR cVar2S18S13P000nsss(0)='1'  OR cVar2S19S13N000P020P002nsss(0)='1'  )then
          oVar1S95(0) <='1';
          else
          oVar1S95(0) <='0';
          end if;
        if(cVar2S20S13N000N020P023nsss(0)='1'  OR cVar2S21S13P032P066P004nsss(0)='1'  OR cVar2S22S13P032P066P014nsss(0)='1'  OR cVar2S23S13N032P030P012nsss(0)='1'  )then
          oVar1S96(0) <='1';
          else
          oVar1S96(0) <='0';
          end if;
        if(cVar2S24S13P055P030P035nsss(0)='1'  OR cVar2S25S13P055N030P028nsss(0)='1'  OR cVar2S26S13N055P022P043nsss(0)='1'  OR cVar2S27S13N055N022P017nsss(0)='1'  )then
          oVar1S97(0) <='1';
          else
          oVar1S97(0) <='0';
          end if;
        if(cVar1S0S14P017P048P025nsss(0)='1'  OR cVar2S1S14P009nsss(0)='1'  OR cVar2S2S14N009P007nsss(0)='1'  OR cVar2S3S14N009N007P008nsss(0)='1'  )then
          oVar1S99(0) <='1';
          else
          oVar1S99(0) <='0';
          end if;
        if(cVar2S4S14P007P011P037nsss(0)='1'  OR cVar2S5S14P007P011P050nsss(0)='1'  OR cVar1S6S14P017N048P044P023nsss(0)='1'  OR cVar2S7S14P022P006nsss(0)='1'  )then
          oVar1S100(0) <='1';
          else
          oVar1S100(0) <='0';
          end if;
        if(cVar2S8S14P022N006P004nsss(0)='1'  OR cVar2S9S14N022P025nsss(0)='1'  OR cVar2S10S14N022N025P058nsss(0)='1'  OR cVar2S11S14P021nsss(0)='1'  )then
          oVar1S101(0) <='1';
          else
          oVar1S101(0) <='0';
          end if;
        if(cVar2S12S14N021P020nsss(0)='1'  OR cVar2S13S14N021N020P013nsss(0)='1'  OR cVar2S14S14P003P046nsss(0)='1'  OR cVar2S15S14P003P039nsss(0)='1'  )then
          oVar1S102(0) <='1';
          else
          oVar1S102(0) <='0';
          end if;
        if(cVar2S16S14P035P068P012nsss(0)='1'  OR cVar2S17S14P035P068P018nsss(0)='1'  OR cVar2S18S14N035P003P011nsss(0)='1'  OR cVar1S19S14P017P064P019P050nsss(0)='1'  )then
          oVar1S103(0) <='1';
          else
          oVar1S103(0) <='0';
          end if;
        if(cVar2S20S14P056nsss(0)='1'  OR cVar2S21S14N056P015P008nsss(0)='1'  OR cVar2S22S14P019P059nsss(0)='1'  OR cVar2S23S14P019N059P063nsss(0)='1'  )then
          oVar1S104(0) <='1';
          else
          oVar1S104(0) <='0';
          end if;
        if(cVar2S24S14P019P014P016nsss(0)='1'  OR cVar2S25S14P019N014P012nsss(0)='1'  OR cVar2S26S14P028nsss(0)='1'  OR cVar2S27S14N028P008nsss(0)='1'  )then
          oVar1S105(0) <='1';
          else
          oVar1S105(0) <='0';
          end if;
        if(cVar2S28S14N028N008P029nsss(0)='1'  OR cVar2S29S14P055P029P031nsss(0)='1'  OR cVar2S30S14N055P048P007nsss(0)='1'  )then
          oVar1S106(0) <='1';
          else
          oVar1S106(0) <='0';
          end if;
        if(cVar1S0S15P044P023P005nsss(0)='1'  OR cVar1S1S15P044P023N005P004nsss(0)='1'  OR cVar2S2S15P007nsss(0)='1'  OR cVar2S3S15N007P006nsss(0)='1'  )then
          oVar1S107(0) <='1';
          else
          oVar1S107(0) <='0';
          end if;
        if(cVar1S4S15P044N023P022P015nsss(0)='1'  OR cVar2S5S15P007nsss(0)='1'  OR cVar2S6S15N007P006nsss(0)='1'  OR cVar2S7S15N007N006P005nsss(0)='1'  )then
          oVar1S108(0) <='1';
          else
          oVar1S108(0) <='0';
          end if;
        if(cVar2S8S15P042nsss(0)='1'  OR cVar2S9S15P042P018P017nsss(0)='1'  OR cVar1S10S15N044P048P025P007nsss(0)='1'  OR cVar2S11S15P006nsss(0)='1'  )then
          oVar1S109(0) <='1';
          else
          oVar1S109(0) <='0';
          end if;
        if(cVar2S12S15N006P009nsss(0)='1'  OR cVar2S13S15N006N009P008nsss(0)='1'  OR cVar2S14S15P052P050nsss(0)='1'  OR cVar2S15S15P052N050P018nsss(0)='1'  )then
          oVar1S110(0) <='1';
          else
          oVar1S110(0) <='0';
          end if;
        if(cVar2S16S15P006P024nsss(0)='1'  OR cVar2S17S15P006N024P016nsss(0)='1'  OR cVar2S18S15N006P065P008nsss(0)='1'  OR cVar2S19S15P002nsss(0)='1'  )then
          oVar1S111(0) <='1';
          else
          oVar1S111(0) <='0';
          end if;
        if(cVar2S20S15N002P004nsss(0)='1'  OR cVar2S21S15N002N004P005nsss(0)='1'  OR cVar2S22S15P042P069P035nsss(0)='1'  OR cVar2S23S15P042P064nsss(0)='1'  )then
          oVar1S112(0) <='1';
          else
          oVar1S112(0) <='0';
          end if;
        if(cVar2S24S15P042N064P005nsss(0)='1'  OR cVar2S25S15P022nsss(0)='1'  OR cVar2S26S15N022P023nsss(0)='1'  OR cVar2S27S15N022N023P025nsss(0)='1'  )then
          oVar1S113(0) <='1';
          else
          oVar1S113(0) <='0';
          end if;
        if(cVar2S28S15P049P025nsss(0)='1'  OR cVar2S29S15P049N025P024nsss(0)='1'  )then
          oVar1S114(0) <='1';
          else
          oVar1S114(0) <='0';
          end if;
        if(cVar1S0S16P067P048P025P050nsss(0)='1'  OR cVar1S1S16P067P048N025P027nsss(0)='1'  OR cVar2S2S16P024P006nsss(0)='1'  OR cVar2S3S16P024N006P046nsss(0)='1'  )then
          oVar1S115(0) <='1';
          else
          oVar1S115(0) <='0';
          end if;
        if(cVar2S4S16N024P007nsss(0)='1'  OR cVar2S5S16P013P028nsss(0)='1'  OR cVar2S6S16P013N028P026nsss(0)='1'  OR cVar2S7S16P013psss(0)='1'  )then
          oVar1S116(0) <='1';
          else
          oVar1S116(0) <='0';
          end if;
        if(cVar2S8S16P036nsss(0)='1'  OR cVar2S9S16P036P015nsss(0)='1'  OR cVar2S10S16P045nsss(0)='1'  OR cVar2S11S16N045P041nsss(0)='1'  )then
          oVar1S117(0) <='1';
          else
          oVar1S117(0) <='0';
          end if;
        if(cVar2S12S16N045N041P044nsss(0)='1'  OR cVar2S13S16P038P040nsss(0)='1'  OR cVar2S14S16P038N040P012nsss(0)='1'  OR cVar2S15S16N038P043nsss(0)='1'  )then
          oVar1S118(0) <='1';
          else
          oVar1S118(0) <='0';
          end if;
        if(cVar2S16S16N038P043P045nsss(0)='1'  OR cVar2S17S16P033P016P034nsss(0)='1'  OR cVar2S18S16P033P016P036nsss(0)='1'  OR cVar2S19S16P033P061nsss(0)='1'  )then
          oVar1S119(0) <='1';
          else
          oVar1S119(0) <='0';
          end if;
        if(cVar2S20S16P014P015nsss(0)='1'  OR cVar2S21S16P013P065nsss(0)='1'  OR cVar2S22S16P013N065P034nsss(0)='1'  OR cVar2S23S16P013P015nsss(0)='1'  )then
          oVar1S120(0) <='1';
          else
          oVar1S120(0) <='0';
          end if;
        if(cVar2S24S16P016P036P014nsss(0)='1'  OR cVar2S25S16P016N036P068nsss(0)='1'  OR cVar2S26S16N016P017P015nsss(0)='1'  OR cVar1S27S16P067N069P052nsss(0)='1'  )then
          oVar1S121(0) <='1';
          else
          oVar1S121(0) <='0';
          end if;
        if(cVar2S28S16P063P015nsss(0)='1'  OR cVar2S29S16P063P034nsss(0)='1'  OR cVar2S30S16P055nsss(0)='1'  )then
          oVar1S122(0) <='1';
          else
          oVar1S122(0) <='0';
          end if;
        if(cVar1S0S17P022P043P062nsss(0)='1'  OR cVar1S1S17P022N043P069P004nsss(0)='1'  OR cVar2S2S17P066P020nsss(0)='1'  OR cVar2S3S17P066N020P024nsss(0)='1'  )then
          oVar1S123(0) <='1';
          else
          oVar1S123(0) <='0';
          end if;
        if(cVar1S4S17N022P048P025P007nsss(0)='1'  OR cVar2S5S17P006nsss(0)='1'  OR cVar2S6S17N006P009nsss(0)='1'  OR cVar2S7S17N006N009P005nsss(0)='1'  )then
          oVar1S124(0) <='1';
          else
          oVar1S124(0) <='0';
          end if;
        if(cVar2S8S17P013nsss(0)='1'  OR cVar2S9S17P024P012nsss(0)='1'  OR cVar2S10S17N024P050P026nsss(0)='1'  OR cVar2S11S17N024N050P014nsss(0)='1'  )then
          oVar1S125(0) <='1';
          else
          oVar1S125(0) <='0';
          end if;
        if(cVar2S12S17P013P028nsss(0)='1'  OR cVar2S13S17P013N028P026nsss(0)='1'  OR cVar2S14S17P013P026nsss(0)='1'  OR cVar2S15S17P010P036nsss(0)='1'  )then
          oVar1S126(0) <='1';
          else
          oVar1S126(0) <='0';
          end if;
        if(cVar2S16S17N010P011nsss(0)='1'  OR cVar2S17S17N010N011P009nsss(0)='1'  OR cVar2S18S17P021P015nsss(0)='1'  OR cVar2S19S17N021P000nsss(0)='1'  )then
          oVar1S127(0) <='1';
          else
          oVar1S127(0) <='0';
          end if;
        if(cVar2S20S17N021N000P004nsss(0)='1'  OR cVar2S21S17P052P009P066nsss(0)='1'  OR cVar2S22S17P052N009P010nsss(0)='1'  OR cVar2S23S17N052P009P061nsss(0)='1'  )then
          oVar1S128(0) <='1';
          else
          oVar1S128(0) <='0';
          end if;
        if(cVar2S24S17N052P009P047nsss(0)='1'  )then
          oVar1S129(0) <='1';
          else
          oVar1S129(0) <='0';
          end if;
        if(cVar1S0S18P041P020nsss(0)='1'  OR cVar1S1S18P041N020P021P039nsss(0)='1'  OR cVar2S2S18P004nsss(0)='1'  OR cVar2S3S18N004P005nsss(0)='1'  )then
          oVar1S130(0) <='1';
          else
          oVar1S130(0) <='0';
          end if;
        if(cVar2S4S18P023nsss(0)='1'  OR cVar2S5S18N023P061nsss(0)='1'  OR cVar2S6S18P023nsss(0)='1'  OR cVar2S7S18N023P004nsss(0)='1'  )then
          oVar1S131(0) <='1';
          else
          oVar1S131(0) <='0';
          end if;
        if(cVar2S8S18N023N004P025nsss(0)='1'  OR cVar2S9S18P042P050nsss(0)='1'  OR cVar2S10S18P042N050P002nsss(0)='1'  OR cVar2S11S18P042P040nsss(0)='1'  )then
          oVar1S132(0) <='1';
          else
          oVar1S132(0) <='0';
          end if;
        if(cVar2S12S18P042N040P064nsss(0)='1'  OR cVar2S13S18P002nsss(0)='1'  OR cVar2S14S18P024nsss(0)='1'  OR cVar2S15S18N024P037P012nsss(0)='1'  )then
          oVar1S133(0) <='1';
          else
          oVar1S133(0) <='0';
          end if;
        if(cVar1S16S18N041P039P005nsss(0)='1'  OR cVar1S17S18N041P039N005P020nsss(0)='1'  OR cVar2S18S18P051nsss(0)='1'  )then
          oVar1S134(0) <='1';
          else
          oVar1S134(0) <='0';
          end if;
        if(cVar1S0S19P041P020nsss(0)='1'  OR cVar1S1S19P041N020P021P003nsss(0)='1'  OR cVar2S2S19P040nsss(0)='1'  OR cVar2S3S19P004nsss(0)='1'  )then
          oVar1S135(0) <='1';
          else
          oVar1S135(0) <='0';
          end if;
        if(cVar2S4S19N004P005nsss(0)='1'  OR cVar2S5S19P023nsss(0)='1'  OR cVar2S6S19N023P047nsss(0)='1'  OR cVar2S7S19N023N047P061nsss(0)='1'  )then
          oVar1S136(0) <='1';
          else
          oVar1S136(0) <='0';
          end if;
        if(cVar2S8S19P005nsss(0)='1'  OR cVar2S9S19N005P004nsss(0)='1'  OR cVar2S10S19N005N004P015nsss(0)='1'  OR cVar1S11S19N041P039P044N023psss(0)='1'  )then
          oVar1S137(0) <='1';
          else
          oVar1S137(0) <='0';
          end if;
        if(cVar2S12S19P009P027nsss(0)='1'  OR cVar2S13S19P009N027P029nsss(0)='1'  OR cVar2S14S19N009P008P011nsss(0)='1'  OR cVar2S15S19N009N008P011nsss(0)='1'  )then
          oVar1S138(0) <='1';
          else
          oVar1S138(0) <='0';
          end if;
        if(cVar2S16S19P000P015P033nsss(0)='1'  OR cVar2S17S19P000N015P054nsss(0)='1'  OR cVar2S18S19P000P040nsss(0)='1'  OR cVar1S19S19N041P039P005nsss(0)='1'  )then
          oVar1S139(0) <='1';
          else
          oVar1S139(0) <='0';
          end if;
        if(cVar2S20S19P020nsss(0)='1'  )then
          oVar1S140(0) <='1';
          else
          oVar1S140(0) <='0';
          end if;
        if(cVar2S0S20P007nsss(0)='1'  OR cVar2S1S20N007P004nsss(0)='1'  OR cVar2S2S20N007N004P006nsss(0)='1'  OR cVar1S3S20P011P029P048N025psss(0)='1'  )then
          oVar1S141(0) <='1';
          else
          oVar1S141(0) <='0';
          end if;
        if(cVar2S4S20P020nsss(0)='1'  OR cVar2S5S20N020P021nsss(0)='1'  OR cVar2S6S20N020N021P022nsss(0)='1'  OR cVar2S7S20P039P007nsss(0)='1'  )then
          oVar1S142(0) <='1';
          else
          oVar1S142(0) <='0';
          end if;
        if(cVar2S8S20P039P007P025nsss(0)='1'  OR cVar2S9S20P039P064nsss(0)='1'  OR cVar2S10S20P039N064P005nsss(0)='1'  OR cVar1S11S20P011P029P010P052nsss(0)='1'  )then
          oVar1S143(0) <='1';
          else
          oVar1S143(0) <='0';
          end if;
        if(cVar2S12S20P054nsss(0)='1'  OR cVar2S13S20P050nsss(0)='1'  OR cVar2S14S20N050P053nsss(0)='1'  OR cVar2S15S20P008P052nsss(0)='1'  )then
          oVar1S144(0) <='1';
          else
          oVar1S144(0) <='0';
          end if;
        if(cVar2S16S20P016P033nsss(0)='1'  OR cVar2S17S20P016P018nsss(0)='1'  OR cVar2S18S20P053nsss(0)='1'  OR cVar2S19S20N053P018nsss(0)='1'  )then
          oVar1S145(0) <='1';
          else
          oVar1S145(0) <='0';
          end if;
        if(cVar2S20S20P003P009nsss(0)='1'  OR cVar2S21S20N003P055nsss(0)='1'  OR cVar2S22S20N003N055P043nsss(0)='1'  OR cVar2S23S20P069P013nsss(0)='1'  )then
          oVar1S146(0) <='1';
          else
          oVar1S146(0) <='0';
          end if;
        if(cVar2S24S20P035P014P008nsss(0)='1'  OR cVar2S25S20P035N014P031nsss(0)='1'  OR cVar2S26S20P035P012P062nsss(0)='1'  OR cVar2S27S20P054P031nsss(0)='1'  )then
          oVar1S147(0) <='1';
          else
          oVar1S147(0) <='0';
          end if;
        if(cVar2S28S20N054P064P049nsss(0)='1'  )then
          oVar1S148(0) <='1';
          else
          oVar1S148(0) <='0';
          end if;
        if(cVar1S0S21P041P020nsss(0)='1'  OR cVar1S1S21P041N020P021P003nsss(0)='1'  OR cVar2S2S21P040nsss(0)='1'  OR cVar1S3S21P041N020N021P004nsss(0)='1'  )then
          oVar1S149(0) <='1';
          else
          oVar1S149(0) <='0';
          end if;
        if(cVar2S4S21P023nsss(0)='1'  OR cVar2S5S21N023P022P005nsss(0)='1'  OR cVar2S6S21N023N022P061nsss(0)='1'  OR cVar2S7S21P025nsss(0)='1'  )then
          oVar1S150(0) <='1';
          else
          oVar1S150(0) <='0';
          end if;
        if(cVar2S8S21N025P027nsss(0)='1'  OR cVar2S9S21N025N027P049nsss(0)='1'  OR cVar2S10S21P051P008P013nsss(0)='1'  OR cVar2S11S21P051N008P019nsss(0)='1'  )then
          oVar1S151(0) <='1';
          else
          oVar1S151(0) <='0';
          end if;
        if(cVar2S12S21N051P055P030nsss(0)='1'  OR cVar1S13S21N041P039P000P040nsss(0)='1'  OR cVar2S14S21P015P014P062nsss(0)='1'  OR cVar2S15S21N015P017P008nsss(0)='1'  )then
          oVar1S152(0) <='1';
          else
          oVar1S152(0) <='0';
          end if;
        if(cVar1S16S21N041P039P051nsss(0)='1'  OR cVar1S17S21N041P039N051P020nsss(0)='1'  )then
          oVar1S153(0) <='1';
          else
          oVar1S153(0) <='0';
          end if;
        if(cVar1S0S22P000P041P020P039nsss(0)='1'  OR cVar2S1S22P021nsss(0)='1'  OR cVar2S2S22N021P017nsss(0)='1'  OR cVar2S3S22P003P021nsss(0)='1'  )then
          oVar1S154(0) <='1';
          else
          oVar1S154(0) <='0';
          end if;
        if(cVar2S4S22N003P022nsss(0)='1'  OR cVar2S5S22N003N022P004nsss(0)='1'  OR cVar2S6S22P030P040nsss(0)='1'  OR cVar2S7S22P030N040P057nsss(0)='1'  )then
          oVar1S155(0) <='1';
          else
          oVar1S155(0) <='0';
          end if;
        if(cVar2S8S22P030P010P009nsss(0)='1'  OR cVar2S9S22P030P031P036nsss(0)='1'  OR cVar2S10S22N030P032P010nsss(0)='1'  OR cVar2S11S22N030N032P017nsss(0)='1'  )then
          oVar1S156(0) <='1';
          else
          oVar1S156(0) <='0';
          end if;
        if(cVar1S12S22P000N041P039P049nsss(0)='1'  OR cVar2S13S22P020nsss(0)='1'  OR cVar2S14S22N020P064nsss(0)='1'  OR cVar2S15S22N020N064P005nsss(0)='1'  )then
          oVar1S157(0) <='1';
          else
          oVar1S157(0) <='0';
          end if;
        if(cVar1S16S22P000P040nsss(0)='1'  OR cVar1S17S22P000N040P059P041nsss(0)='1'  OR cVar2S18S22P018P012P016nsss(0)='1'  OR cVar2S19S22N018P052nsss(0)='1'  )then
          oVar1S158(0) <='1';
          else
          oVar1S158(0) <='0';
          end if;
        if(cVar1S0S23P041P020P010nsss(0)='1'  OR cVar1S1S23P041N020P005P021nsss(0)='1'  OR cVar2S2S23P022nsss(0)='1'  OR cVar2S3S23N022P042nsss(0)='1'  )then
          oVar1S160(0) <='1';
          else
          oVar1S160(0) <='0';
          end if;
        if(cVar2S4S23P021nsss(0)='1'  OR cVar2S5S23P004nsss(0)='1'  OR cVar2S6S23P010P028nsss(0)='1'  OR cVar2S7S23P010N028P030nsss(0)='1'  )then
          oVar1S161(0) <='1';
          else
          oVar1S161(0) <='0';
          end if;
        if(cVar2S8S23N010P058nsss(0)='1'  OR cVar2S9S23P029P033nsss(0)='1'  OR cVar1S10S23N041P055P061P054nsss(0)='1'  OR cVar2S11S23P030nsss(0)='1'  )then
          oVar1S162(0) <='1';
          else
          oVar1S162(0) <='0';
          end if;
        if(cVar2S12S23P008P026nsss(0)='1'  OR cVar2S13S23P008N026P027nsss(0)='1'  OR cVar2S14S23N008P038nsss(0)='1'  OR cVar2S15S23N008N038P058nsss(0)='1'  )then
          oVar1S163(0) <='1';
          else
          oVar1S163(0) <='0';
          end if;
        if(cVar2S16S23P005nsss(0)='1'  OR cVar2S17S23P035P069nsss(0)='1'  OR cVar2S18S23P029P063P008nsss(0)='1'  OR cVar2S19S23N029P030P014nsss(0)='1'  )then
          oVar1S164(0) <='1';
          else
          oVar1S164(0) <='0';
          end if;
        if(cVar1S0S24P041P020P039nsss(0)='1'  OR cVar1S1S24P041N020P005P021nsss(0)='1'  OR cVar2S2S24P022nsss(0)='1'  OR cVar2S3S24N022P042nsss(0)='1'  )then
          oVar1S166(0) <='1';
          else
          oVar1S166(0) <='0';
          end if;
        if(cVar2S4S24P021nsss(0)='1'  OR cVar2S5S24P022P004nsss(0)='1'  OR cVar2S6S24N022P061nsss(0)='1'  OR cVar2S7S24P060P013nsss(0)='1'  )then
          oVar1S167(0) <='1';
          else
          oVar1S167(0) <='0';
          end if;
        if(cVar2S8S24P060P013P031nsss(0)='1'  OR cVar2S9S24P060P035P064nsss(0)='1'  OR cVar2S10S24P060N035P066nsss(0)='1'  OR cVar2S11S24P063P014P016nsss(0)='1'  )then
          oVar1S168(0) <='1';
          else
          oVar1S168(0) <='0';
          end if;
        if(cVar2S12S24P063N014P062nsss(0)='1'  OR cVar2S13S24P063P034P016nsss(0)='1'  OR cVar2S14S24P001P010nsss(0)='1'  OR cVar2S15S24P056P013nsss(0)='1'  )then
          oVar1S169(0) <='1';
          else
          oVar1S169(0) <='0';
          end if;
        if(cVar2S16S24P056N013P012nsss(0)='1'  OR cVar2S17S24N056P014P032nsss(0)='1'  OR cVar1S18S24N041P039P051nsss(0)='1'  OR cVar1S19S24N041P039N051P064nsss(0)='1'  )then
          oVar1S170(0) <='1';
          else
          oVar1S170(0) <='0';
          end if;
        if(cVar2S20S24P010P020nsss(0)='1'  )then
          oVar1S171(0) <='1';
          else
          oVar1S171(0) <='0';
          end if;
        if(cVar1S0S25P041P020nsss(0)='1'  OR cVar1S1S25P041N020P005P021nsss(0)='1'  OR cVar2S2S25P017nsss(0)='1'  OR cVar2S3S25P021nsss(0)='1'  )then
          oVar1S172(0) <='1';
          else
          oVar1S172(0) <='0';
          end if;
        if(cVar2S4S25P065P022nsss(0)='1'  OR cVar2S5S25P065N022P018nsss(0)='1'  OR cVar2S6S25P016P010nsss(0)='1'  OR cVar2S7S25P016P019nsss(0)='1'  )then
          oVar1S173(0) <='1';
          else
          oVar1S173(0) <='0';
          end if;
        if(cVar2S8S25P057nsss(0)='1'  OR cVar2S9S25N057P060P019nsss(0)='1'  OR cVar2S10S25P065P019P020nsss(0)='1'  OR cVar2S11S25P065N019psss(0)='1'  )then
          oVar1S174(0) <='1';
          else
          oVar1S174(0) <='0';
          end if;
        if(cVar2S12S25P065P059P017nsss(0)='1'  OR cVar2S13S25P062P017P047nsss(0)='1'  OR cVar2S14S25P062N017P057nsss(0)='1'  OR cVar2S15S25P023nsss(0)='1'  )then
          oVar1S175(0) <='1';
          else
          oVar1S175(0) <='0';
          end if;
        if(cVar2S16S25N023P022nsss(0)='1'  OR cVar2S17S25P064P037P062nsss(0)='1'  OR cVar2S18S25N064P037P068nsss(0)='1'  OR cVar2S19S25N064N037P022nsss(0)='1'  )then
          oVar1S176(0) <='1';
          else
          oVar1S176(0) <='0';
          end if;
        if(cVar2S20S25P016P054nsss(0)='1'  OR cVar2S21S25P016N054P057nsss(0)='1'  OR cVar2S22S25P012P056nsss(0)='1'  )then
          oVar1S177(0) <='1';
          else
          oVar1S177(0) <='0';
          end if;
        if(cVar1S0S26P068P041P020P016nsss(0)='1'  OR cVar2S1S26P039nsss(0)='1'  OR cVar2S2S26N039P023nsss(0)='1'  OR cVar2S3S26P003nsss(0)='1'  )then
          oVar1S178(0) <='1';
          else
          oVar1S178(0) <='0';
          end if;
        if(cVar2S4S26N003P022nsss(0)='1'  OR cVar2S5S26P047nsss(0)='1'  OR cVar2S6S26N047P045nsss(0)='1'  OR cVar2S7S26N047N045P046nsss(0)='1'  )then
          oVar1S179(0) <='1';
          else
          oVar1S179(0) <='0';
          end if;
        if(cVar2S8S26P007P045nsss(0)='1'  OR cVar2S9S26P007N045P049nsss(0)='1'  OR cVar2S10S26P005P042nsss(0)='1'  OR cVar2S11S26P005N042P045nsss(0)='1'  )then
          oVar1S180(0) <='1';
          else
          oVar1S180(0) <='0';
          end if;
        if(cVar2S12S26N005P042nsss(0)='1'  OR cVar2S13S26N005N042P007nsss(0)='1'  OR cVar2S14S26P045P043P042nsss(0)='1'  OR cVar2S15S26P045P022nsss(0)='1'  )then
          oVar1S181(0) <='1';
          else
          oVar1S181(0) <='0';
          end if;
        if(cVar2S16S26P045N022P025nsss(0)='1'  OR cVar2S17S26P045P027nsss(0)='1'  OR cVar2S18S26P045P027P015nsss(0)='1'  OR cVar2S19S26P067P007P061nsss(0)='1'  )then
          oVar1S182(0) <='1';
          else
          oVar1S182(0) <='0';
          end if;
        if(cVar2S20S26P067P007P012nsss(0)='1'  OR cVar2S21S26P067P062nsss(0)='1'  OR cVar2S22S26P018P062P006nsss(0)='1'  OR cVar2S23S26N018P069P016nsss(0)='1'  )then
          oVar1S183(0) <='1';
          else
          oVar1S183(0) <='0';
          end if;
        if(cVar2S24S26N018N069P057nsss(0)='1'  OR cVar2S25S26P019nsss(0)='1'  OR cVar2S26S26N019P017nsss(0)='1'  OR cVar2S27S26P064P016nsss(0)='1'  )then
          oVar1S184(0) <='1';
          else
          oVar1S184(0) <='0';
          end if;
        if(cVar2S28S26P034P064nsss(0)='1'  OR cVar2S29S26P034N064P019nsss(0)='1'  OR cVar2S30S26P014P034nsss(0)='1'  OR cVar2S31S26N014P063P018nsss(0)='1'  )then
          oVar1S185(0) <='1';
          else
          oVar1S185(0) <='0';
          end if;
        if(cVar1S0S27P041P020P003nsss(0)='1'  OR cVar1S1S27P041P020N003P002nsss(0)='1'  OR cVar2S2S27P004nsss(0)='1'  OR cVar2S3S27N004P005nsss(0)='1'  )then
          oVar1S187(0) <='1';
          else
          oVar1S187(0) <='0';
          end if;
        if(cVar2S4S27P039nsss(0)='1'  OR cVar2S5S27N039P023nsss(0)='1'  OR cVar2S6S27P034P065nsss(0)='1'  OR cVar2S7S27P019nsss(0)='1'  )then
          oVar1S188(0) <='1';
          else
          oVar1S188(0) <='0';
          end if;
        if(cVar1S8S27N041P024P006P047nsss(0)='1'  OR cVar2S9S27P045nsss(0)='1'  OR cVar2S10S27N045P044nsss(0)='1'  OR cVar2S11S27N045N044P046nsss(0)='1'  )then
          oVar1S189(0) <='1';
          else
          oVar1S189(0) <='0';
          end if;
        if(cVar2S12S27P068P007nsss(0)='1'  OR cVar2S13S27P068N007P017nsss(0)='1'  OR cVar2S14S27P045nsss(0)='1'  OR cVar2S15S27N045P068P011nsss(0)='1'  )then
          oVar1S190(0) <='1';
          else
          oVar1S190(0) <='0';
          end if;
        if(cVar2S16S27P042nsss(0)='1'  OR cVar2S17S27N042P045nsss(0)='1'  OR cVar2S18S27P042P004nsss(0)='1'  OR cVar2S19S27P042N004P017nsss(0)='1'  )then
          oVar1S191(0) <='1';
          else
          oVar1S191(0) <='0';
          end if;
        if(cVar2S20S27N042P007nsss(0)='1'  OR cVar2S21S27N042N007P008nsss(0)='1'  OR cVar2S22S27P009P027P011nsss(0)='1'  OR cVar2S23S27P009N027P029nsss(0)='1'  )then
          oVar1S192(0) <='1';
          else
          oVar1S192(0) <='0';
          end if;
        if(cVar2S24S27N009P026nsss(0)='1'  OR cVar2S25S27N009N026P055nsss(0)='1'  OR cVar2S26S27P005P069P036nsss(0)='1'  OR cVar2S27S27P005P022nsss(0)='1'  )then
          oVar1S193(0) <='1';
          else
          oVar1S193(0) <='0';
          end if;
        if(cVar2S28S27P005N022P025nsss(0)='1'  )then
          oVar1S194(0) <='1';
          else
          oVar1S194(0) <='0';
          end if;
        if(cVar1S0S28P024P006P047nsss(0)='1'  OR cVar1S1S28P024P006N047P045nsss(0)='1'  OR cVar2S2S28P044nsss(0)='1'  OR cVar2S3S28N044P048nsss(0)='1'  )then
          oVar1S195(0) <='1';
          else
          oVar1S195(0) <='0';
          end if;
        if(cVar2S4S28P007nsss(0)='1'  OR cVar2S5S28N007P025nsss(0)='1'  OR cVar2S6S28P015nsss(0)='1'  OR cVar1S7S28P024N006P068P047nsss(0)='1'  )then
          oVar1S196(0) <='1';
          else
          oVar1S196(0) <='0';
          end if;
        if(cVar1S8S28N024P040P002nsss(0)='1'  OR cVar1S9S28N024P040N002P004nsss(0)='1'  OR cVar2S10S28P005nsss(0)='1'  OR cVar2S11S28N005P003P015nsss(0)='1'  )then
          oVar1S197(0) <='1';
          else
          oVar1S197(0) <='0';
          end if;
        if(cVar2S12S28P005nsss(0)='1'  OR cVar2S13S28N005P004nsss(0)='1'  OR cVar2S14S28N005N004P007nsss(0)='1'  OR cVar2S15S28P025P014nsss(0)='1'  )then
          oVar1S198(0) <='1';
          else
          oVar1S198(0) <='0';
          end if;
        if(cVar2S16S28N025P054nsss(0)='1'  OR cVar2S17S28N025N054P022nsss(0)='1'  OR cVar2S18S28P021nsss(0)='1'  OR cVar2S19S28P021P039nsss(0)='1'  )then
          oVar1S199(0) <='1';
          else
          oVar1S199(0) <='0';
          end if;
        if(cVar2S20S28P021N039P055nsss(0)='1'  OR cVar2S21S28P058nsss(0)='1'  OR cVar2S22S28N058P043nsss(0)='1'  )then
          oVar1S200(0) <='1';
          else
          oVar1S200(0) <='0';
          end if;
        if(cVar1S0S29P024P006P047nsss(0)='1'  OR cVar1S1S29P024P006N047P045nsss(0)='1'  OR cVar2S2S29P044nsss(0)='1'  OR cVar2S3S29N044P048nsss(0)='1'  )then
          oVar1S201(0) <='1';
          else
          oVar1S201(0) <='0';
          end if;
        if(cVar2S4S29P045nsss(0)='1'  OR cVar2S5S29N045P049nsss(0)='1'  OR cVar2S6S29P025P057nsss(0)='1'  OR cVar1S7S29P024N006P068P012nsss(0)='1'  )then
          oVar1S202(0) <='1';
          else
          oVar1S202(0) <='0';
          end if;
        if(cVar2S8S29P008nsss(0)='1'  OR cVar1S9S29N024P040P002nsss(0)='1'  OR cVar2S10S29P021P003nsss(0)='1'  OR cVar2S11S29P021N003P005nsss(0)='1'  )then
          oVar1S203(0) <='1';
          else
          oVar1S203(0) <='0';
          end if;
        if(cVar2S12S29N021P066nsss(0)='1'  OR cVar2S13S29N021P066P017nsss(0)='1'  OR cVar2S14S29P005nsss(0)='1'  OR cVar2S15S29N005P004nsss(0)='1'  )then
          oVar1S204(0) <='1';
          else
          oVar1S204(0) <='0';
          end if;
        if(cVar2S16S29N005N004P007nsss(0)='1'  OR cVar2S17S29P025P015nsss(0)='1'  OR cVar2S18S29N025psss(0)='1'  OR cVar2S19S29P020P003nsss(0)='1'  )then
          oVar1S205(0) <='1';
          else
          oVar1S205(0) <='0';
          end if;
        if(cVar2S20S29P020N003P002nsss(0)='1'  OR cVar2S21S29N020P005nsss(0)='1'  OR cVar2S22S29N020N005P003nsss(0)='1'  OR cVar2S23S29P039P005P043nsss(0)='1'  )then
          oVar1S206(0) <='1';
          else
          oVar1S206(0) <='0';
          end if;
        if(cVar1S0S30P067P018P048P025nsss(0)='1'  OR cVar2S1S30P027nsss(0)='1'  OR cVar2S2S30N027P024nsss(0)='1'  OR cVar2S3S30N027N024P013nsss(0)='1'  )then
          oVar1S208(0) <='1';
          else
          oVar1S208(0) <='0';
          end if;
        if(cVar2S4S30P034P015P035nsss(0)='1'  OR cVar2S5S30P034P015P063nsss(0)='1'  OR cVar2S6S30N034P032P065nsss(0)='1'  OR cVar2S7S30N034N032psss(0)='1'  )then
          oVar1S209(0) <='1';
          else
          oVar1S209(0) <='0';
          end if;
        if(cVar2S8S30P030P031nsss(0)='1'  OR cVar2S9S30N030psss(0)='1'  OR cVar2S10S30P003nsss(0)='1'  OR cVar2S11S30N003P029nsss(0)='1'  )then
          oVar1S210(0) <='1';
          else
          oVar1S210(0) <='0';
          end if;
        if(cVar2S12S30N003N029P069nsss(0)='1'  OR cVar2S13S30P054P024nsss(0)='1'  OR cVar2S14S30P054N024P040nsss(0)='1'  OR cVar2S15S30P054P013P031nsss(0)='1'  )then
          oVar1S211(0) <='1';
          else
          oVar1S211(0) <='0';
          end if;
        if(cVar2S16S30P033nsss(0)='1'  OR cVar2S17S30N033P062P017nsss(0)='1'  OR cVar2S18S30P050nsss(0)='1'  OR cVar2S19S30N050P035P058nsss(0)='1'  )then
          oVar1S212(0) <='1';
          else
          oVar1S212(0) <='0';
          end if;
        if(cVar2S20S30P060P052nsss(0)='1'  OR cVar2S21S30P060N052P009nsss(0)='1'  OR cVar2S22S30P060P017nsss(0)='1'  OR cVar2S23S30P031P048P064nsss(0)='1'  )then
          oVar1S213(0) <='1';
          else
          oVar1S213(0) <='0';
          end if;
        if(cVar2S24S30P036nsss(0)='1'  OR cVar2S25S30P036P066P012nsss(0)='1'  OR cVar2S26S30P016P036P037nsss(0)='1'  OR cVar2S27S30P016N036P068nsss(0)='1'  )then
          oVar1S214(0) <='1';
          else
          oVar1S214(0) <='0';
          end if;
        if(cVar2S28S30N016P017P015nsss(0)='1'  OR cVar1S29S30P067N069P065P063nsss(0)='1'  OR cVar2S30S30P034nsss(0)='1'  OR cVar1S31S30P067N069N065P052nsss(0)='1'  )then
          oVar1S215(0) <='1';
          else
          oVar1S215(0) <='0';
          end if;
        if(cVar2S32S30P063P061nsss(0)='1'  )then
          oVar1S216(0) <='1';
          else
          oVar1S216(0) <='0';
          end if;
        if(cVar2S0S31P063P016nsss(0)='1'  OR cVar2S1S31P063P016P069nsss(0)='1'  OR cVar2S2S31P063P034P068nsss(0)='1'  OR cVar2S3S31P064P050nsss(0)='1'  )then
          oVar1S217(0) <='1';
          else
          oVar1S217(0) <='0';
          end if;
        if(cVar2S4S31P064N050P059nsss(0)='1'  OR cVar2S5S31N064P015P017nsss(0)='1'  OR cVar2S6S31P015nsss(0)='1'  OR cVar2S7S31P065P013P056nsss(0)='1'  )then
          oVar1S218(0) <='1';
          else
          oVar1S218(0) <='0';
          end if;
        if(cVar1S8S31P018P060P029P050nsss(0)='1'  OR cVar2S9S31P030P014P032nsss(0)='1'  OR cVar2S10S31P030N014P015nsss(0)='1'  OR cVar1S11S31N018P048P025P007nsss(0)='1'  )then
          oVar1S219(0) <='1';
          else
          oVar1S219(0) <='0';
          end if;
        if(cVar2S12S31P006nsss(0)='1'  OR cVar2S13S31N006P009nsss(0)='1'  OR cVar1S14S31N018P048N025P036nsss(0)='1'  OR cVar2S15S31P033P035nsss(0)='1'  )then
          oVar1S220(0) <='1';
          else
          oVar1S220(0) <='0';
          end if;
        if(cVar2S16S31P032P010nsss(0)='1'  OR cVar2S17S31N032P008P006nsss(0)='1'  OR cVar2S18S31N032N008P012nsss(0)='1'  OR cVar2S19S31P012P016P011nsss(0)='1'  )then
          oVar1S221(0) <='1';
          else
          oVar1S221(0) <='0';
          end if;
        if(cVar2S20S31P012P016P015nsss(0)='1'  OR cVar2S21S31N012P010nsss(0)='1'  OR cVar2S22S31N012N010P013nsss(0)='1'  OR cVar2S23S31P023P005nsss(0)='1'  )then
          oVar1S222(0) <='1';
          else
          oVar1S222(0) <='0';
          end if;
        if(cVar2S24S31P023N005P042nsss(0)='1'  OR cVar2S25S31N023P005P015nsss(0)='1'  OR cVar2S26S31N023P005P021nsss(0)='1'  )then
          oVar1S223(0) <='1';
          else
          oVar1S223(0) <='0';
          end if;
        if(cVar1S0S32P015P018P040P021nsss(0)='1'  OR cVar2S1S32P020nsss(0)='1'  OR cVar2S2S32N020P023nsss(0)='1'  OR cVar2S3S32N020N023P022nsss(0)='1'  )then
          oVar1S224(0) <='1';
          else
          oVar1S224(0) <='0';
          end if;
        if(cVar2S4S32P016P012P010nsss(0)='1'  OR cVar2S5S32P016P012P034nsss(0)='1'  OR cVar2S6S32N016P017P019nsss(0)='1'  OR cVar2S7S32N016N017P014nsss(0)='1'  )then
          oVar1S225(0) <='1';
          else
          oVar1S225(0) <='0';
          end if;
        if(cVar2S8S32P016P036nsss(0)='1'  OR cVar2S9S32P016P036P017nsss(0)='1'  OR cVar2S10S32P016P062P012nsss(0)='1'  OR cVar2S11S32P016N062P036nsss(0)='1'  )then
          oVar1S226(0) <='1';
          else
          oVar1S226(0) <='0';
          end if;
        if(cVar2S12S32P057P017nsss(0)='1'  OR cVar2S13S32P057N017P069nsss(0)='1'  OR cVar2S14S32P057P013P030nsss(0)='1'  OR cVar2S15S32P057N013P051nsss(0)='1'  )then
          oVar1S227(0) <='1';
          else
          oVar1S227(0) <='0';
          end if;
        if(cVar2S16S32P065P036P037nsss(0)='1'  OR cVar2S17S32P065P037P019nsss(0)='1'  OR cVar1S18S32P015P018P004P041nsss(0)='1'  OR cVar2S19S32P006nsss(0)='1'  )then
          oVar1S228(0) <='1';
          else
          oVar1S228(0) <='0';
          end if;
        if(cVar2S20S32N006P042nsss(0)='1'  OR cVar2S21S32N006N042P045nsss(0)='1'  OR cVar2S22S32P033P018P016nsss(0)='1'  OR cVar2S23S32P033P018P061nsss(0)='1'  )then
          oVar1S229(0) <='1';
          else
          oVar1S229(0) <='0';
          end if;
        if(cVar2S24S32N033P035P058nsss(0)='1'  OR cVar2S25S32N033N035P037nsss(0)='1'  OR cVar2S26S32P010nsss(0)='1'  OR cVar2S27S32P010P055nsss(0)='1'  )then
          oVar1S230(0) <='1';
          else
          oVar1S230(0) <='0';
          end if;
        if(cVar2S28S32P064P035P013nsss(0)='1'  OR cVar2S29S32P064N035P016nsss(0)='1'  OR cVar2S30S32N064P007nsss(0)='1'  OR cVar2S31S32N064N007P012nsss(0)='1'  )then
          oVar1S231(0) <='1';
          else
          oVar1S231(0) <='0';
          end if;
        if(cVar1S32S32P015P017P008P066nsss(0)='1'  OR cVar2S33S32P012P018nsss(0)='1'  OR cVar2S34S32P049P013nsss(0)='1'  OR cVar2S35S32N049P014P032nsss(0)='1'  )then
          oVar1S232(0) <='1';
          else
          oVar1S232(0) <='0';
          end if;
        if(cVar2S36S32P066nsss(0)='1'  )then
          oVar1S233(0) <='1';
          else
          oVar1S233(0) <='0';
          end if;
        if(cVar2S0S33P034P035nsss(0)='1'  OR cVar2S1S33P034P035P014nsss(0)='1'  OR cVar2S2S33N034P036P037nsss(0)='1'  OR cVar2S3S33N034N036P035nsss(0)='1'  )then
          oVar1S234(0) <='1';
          else
          oVar1S234(0) <='0';
          end if;
        if(cVar2S4S33P032P057P067nsss(0)='1'  OR cVar2S5S33P054nsss(0)='1'  OR cVar2S6S33P062P004nsss(0)='1'  OR cVar2S7S33P062N004P019nsss(0)='1'  )then
          oVar1S235(0) <='1';
          else
          oVar1S235(0) <='0';
          end if;
        if(cVar2S8S33P062P008P034nsss(0)='1'  OR cVar2S9S33P064P010P017nsss(0)='1'  OR cVar2S10S33N064P066P017nsss(0)='1'  OR cVar2S11S33N064N066P000nsss(0)='1'  )then
          oVar1S236(0) <='1';
          else
          oVar1S236(0) <='0';
          end if;
        if(cVar2S12S33P012P015nsss(0)='1'  OR cVar2S13S33N012P014P019nsss(0)='1'  OR cVar2S14S33P069P061nsss(0)='1'  OR cVar2S15S33N069P011P019nsss(0)='1'  )then
          oVar1S237(0) <='1';
          else
          oVar1S237(0) <='0';
          end if;
        if(cVar2S16S33P002nsss(0)='1'  OR cVar2S17S33N002P003nsss(0)='1'  OR cVar2S18S33N002N003P004nsss(0)='1'  OR cVar2S19S33P004nsss(0)='1'  )then
          oVar1S238(0) <='1';
          else
          oVar1S238(0) <='0';
          end if;
        if(cVar2S20S33N004P009nsss(0)='1'  OR cVar2S21S33P023nsss(0)='1'  OR cVar2S22S33N023P006nsss(0)='1'  OR cVar2S23S33N023N006P054nsss(0)='1'  )then
          oVar1S239(0) <='1';
          else
          oVar1S239(0) <='0';
          end if;
        if(cVar2S24S33P050P014nsss(0)='1'  OR cVar2S25S33P050P014P068nsss(0)='1'  OR cVar2S26S33N050P065P041nsss(0)='1'  OR cVar2S27S33N050P065P017nsss(0)='1'  )then
          oVar1S240(0) <='1';
          else
          oVar1S240(0) <='0';
          end if;
        if(cVar2S28S33P066P056P013nsss(0)='1'  OR cVar2S29S33P066P012nsss(0)='1'  OR cVar2S30S33P066N012P065nsss(0)='1'  OR cVar2S31S33P064P035P066nsss(0)='1'  )then
          oVar1S241(0) <='1';
          else
          oVar1S241(0) <='0';
          end if;
        if(cVar2S0S34P026nsss(0)='1'  OR cVar2S1S34N026P024nsss(0)='1'  OR cVar2S2S34P051P016P066nsss(0)='1'  OR cVar2S3S34P051P016P026nsss(0)='1'  )then
          oVar1S243(0) <='1';
          else
          oVar1S243(0) <='0';
          end if;
        if(cVar2S4S34N051P027nsss(0)='1'  OR cVar2S5S34N051N027P065nsss(0)='1'  OR cVar2S6S34P058P033P034nsss(0)='1'  OR cVar2S7S34P058N033P012nsss(0)='1'  )then
          oVar1S244(0) <='1';
          else
          oVar1S244(0) <='0';
          end if;
        if(cVar2S8S34N058P060nsss(0)='1'  OR cVar2S9S34N058P060P057nsss(0)='1'  OR cVar2S10S34P063P017P034nsss(0)='1'  OR cVar2S11S34P063N017P018nsss(0)='1'  )then
          oVar1S245(0) <='1';
          else
          oVar1S245(0) <='0';
          end if;
        if(cVar2S12S34N063P037P013nsss(0)='1'  OR cVar2S13S34N063N037P015nsss(0)='1'  OR cVar2S14S34P010P011P034nsss(0)='1'  OR cVar2S15S34P010P011P060nsss(0)='1'  )then
          oVar1S246(0) <='1';
          else
          oVar1S246(0) <='0';
          end if;
        if(cVar2S16S34P010P017P015nsss(0)='1'  OR cVar2S17S34P016P034nsss(0)='1'  OR cVar2S18S34P016N034P036nsss(0)='1'  OR cVar2S19S34N016P065P056nsss(0)='1'  )then
          oVar1S247(0) <='1';
          else
          oVar1S247(0) <='0';
          end if;
        if(cVar1S20S34P067P062P055P068nsss(0)='1'  OR cVar2S21S34P054P052nsss(0)='1'  OR cVar2S22S34P054N052P028nsss(0)='1'  OR cVar2S23S34P054P011nsss(0)='1'  )then
          oVar1S248(0) <='1';
          else
          oVar1S248(0) <='0';
          end if;
        if(cVar2S24S34P058P057nsss(0)='1'  OR cVar1S25S34P067P010N069P052nsss(0)='1'  OR cVar2S26S34P069P017nsss(0)='1'  OR cVar2S27S34P016nsss(0)='1'  )then
          oVar1S249(0) <='1';
          else
          oVar1S249(0) <='0';
          end if;
        if(cVar1S28S34P067P010N015P050nsss(0)='1'  OR cVar2S29S34P005P053nsss(0)='1'  )then
          oVar1S250(0) <='1';
          else
          oVar1S250(0) <='0';
          end if;
        if(cVar2S0S35P031nsss(0)='1'  OR cVar2S1S35N031P033nsss(0)='1'  OR cVar2S2S35N031N033P037nsss(0)='1'  OR cVar2S3S35P012P068nsss(0)='1'  )then
          oVar1S251(0) <='1';
          else
          oVar1S251(0) <='0';
          end if;
        if(cVar2S4S35P031P014P060nsss(0)='1'  OR cVar2S5S35P031N014P011nsss(0)='1'  OR cVar2S6S35P031P012nsss(0)='1'  OR cVar2S7S35P069P009P014nsss(0)='1'  )then
          oVar1S252(0) <='1';
          else
          oVar1S252(0) <='0';
          end if;
        if(cVar2S8S35P056nsss(0)='1'  OR cVar2S9S35N056P057nsss(0)='1'  OR cVar2S10S35N056N057P059nsss(0)='1'  OR cVar2S11S35P057nsss(0)='1'  )then
          oVar1S253(0) <='1';
          else
          oVar1S253(0) <='0';
          end if;
        if(cVar2S12S35N057P054nsss(0)='1'  OR cVar2S13S35P013P057nsss(0)='1'  OR cVar2S14S35P047nsss(0)='1'  OR cVar2S15S35N047P043nsss(0)='1'  )then
          oVar1S254(0) <='1';
          else
          oVar1S254(0) <='0';
          end if;
        if(cVar2S16S35N047N043P044nsss(0)='1'  OR cVar2S17S35P025P047P066nsss(0)='1'  OR cVar2S18S35P025N047P045nsss(0)='1'  OR cVar2S19S35P057P052P054nsss(0)='1'  )then
          oVar1S255(0) <='1';
          else
          oVar1S255(0) <='0';
          end if;
        if(cVar2S20S35P057P052P067nsss(0)='1'  OR cVar2S21S35P057P068P018nsss(0)='1'  OR cVar2S22S35P031P054nsss(0)='1'  OR cVar2S23S35P031N054P013nsss(0)='1'  )then
          oVar1S256(0) <='1';
          else
          oVar1S256(0) <='0';
          end if;
        if(cVar2S24S35N031P028P010nsss(0)='1'  OR cVar2S25S35N031N028P029nsss(0)='1'  )then
          oVar1S257(0) <='1';
          else
          oVar1S257(0) <='0';
          end if;
        if(cVar1S0S36P037P048P025P067nsss(0)='1'  OR cVar2S1S36P027nsss(0)='1'  OR cVar2S2S36N027P013nsss(0)='1'  OR cVar2S3S36P024P014nsss(0)='1'  )then
          oVar1S258(0) <='1';
          else
          oVar1S258(0) <='0';
          end if;
        if(cVar2S4S36N024P052P030nsss(0)='1'  OR cVar2S5S36P027P050nsss(0)='1'  OR cVar2S6S36P027P007nsss(0)='1'  OR cVar2S7S36P027N007P050nsss(0)='1'  )then
          oVar1S259(0) <='1';
          else
          oVar1S259(0) <='0';
          end if;
        if(cVar2S8S36P049P017nsss(0)='1'  OR cVar2S9S36N049P052P013nsss(0)='1'  OR cVar2S10S36N049N052P007nsss(0)='1'  OR cVar2S11S36P025P007nsss(0)='1'  )then
          oVar1S260(0) <='1';
          else
          oVar1S260(0) <='0';
          end if;
        if(cVar2S12S36P025N007P006nsss(0)='1'  OR cVar2S13S36N025P004nsss(0)='1'  OR cVar2S14S36N025N004P018nsss(0)='1'  OR cVar2S15S36P019P017nsss(0)='1'  )then
          oVar1S261(0) <='1';
          else
          oVar1S261(0) <='0';
          end if;
        if(cVar2S16S36P014nsss(0)='1'  OR cVar2S17S36N014P067P024nsss(0)='1'  OR cVar2S18S36P036P025P046nsss(0)='1'  OR cVar2S19S36P036P014P069nsss(0)='1'  )then
          oVar1S262(0) <='1';
          else
          oVar1S262(0) <='0';
          end if;
        if(cVar2S20S36P036N014P013nsss(0)='1'  OR cVar2S21S36P033P003P010nsss(0)='1'  OR cVar1S22S36P037P059P008nsss(0)='1'  OR cVar2S23S36P062nsss(0)='1'  )then
          oVar1S263(0) <='1';
          else
          oVar1S263(0) <='0';
          end if;
        if(cVar2S24S36P014P068P064nsss(0)='1'  )then
          oVar1S264(0) <='1';
          else
          oVar1S264(0) <='0';
          end if;
        if(cVar1S0S37P048P025P007nsss(0)='1'  OR cVar1S1S37P048P025N007P004nsss(0)='1'  OR cVar2S2S37P006nsss(0)='1'  OR cVar2S3S37N006P009nsss(0)='1'  )then
          oVar1S265(0) <='1';
          else
          oVar1S265(0) <='0';
          end if;
        if(cVar2S4S37N006N009P005nsss(0)='1'  OR cVar1S5S37P048N025P037P017nsss(0)='1'  OR cVar2S6S37P060nsss(0)='1'  OR cVar2S7S37N060P007nsss(0)='1'  )then
          oVar1S266(0) <='1';
          else
          oVar1S266(0) <='0';
          end if;
        if(cVar2S8S37N060N007P008nsss(0)='1'  OR cVar1S9S37P048N025P037P006nsss(0)='1'  OR cVar2S10S37P036P062nsss(0)='1'  OR cVar1S11S37N048P044P004nsss(0)='1'  )then
          oVar1S267(0) <='1';
          else
          oVar1S267(0) <='0';
          end if;
        if(cVar2S12S37P023nsss(0)='1'  OR cVar2S13S37N023P046nsss(0)='1'  OR cVar2S14S37P006P024nsss(0)='1'  OR cVar2S15S37P006N024P025nsss(0)='1'  )then
          oVar1S268(0) <='1';
          else
          oVar1S268(0) <='0';
          end if;
        if(cVar2S16S37N006P021nsss(0)='1'  OR cVar2S17S37N006N021P007nsss(0)='1'  OR cVar2S18S37P026P049nsss(0)='1'  OR cVar2S19S37P026N049P055nsss(0)='1'  )then
          oVar1S269(0) <='1';
          else
          oVar1S269(0) <='0';
          end if;
        if(cVar2S20S37N026P024P047nsss(0)='1'  OR cVar2S21S37P007P047nsss(0)='1'  OR cVar2S22S37P007N047P043nsss(0)='1'  OR cVar2S23S37N007P009nsss(0)='1'  )then
          oVar1S270(0) <='1';
          else
          oVar1S270(0) <='0';
          end if;
        if(cVar2S24S37P054nsss(0)='1'  )then
          oVar1S271(0) <='1';
          else
          oVar1S271(0) <='0';
          end if;
        if(cVar1S0S38P048P025P007nsss(0)='1'  OR cVar1S1S38P048P025N007P004nsss(0)='1'  OR cVar2S2S38P009nsss(0)='1'  OR cVar2S3S38N009P006nsss(0)='1'  )then
          oVar1S272(0) <='1';
          else
          oVar1S272(0) <='0';
          end if;
        if(cVar2S4S38N009N006P005nsss(0)='1'  OR cVar2S5S38P007nsss(0)='1'  OR cVar2S6S38N007P006nsss(0)='1'  OR cVar2S7S38N007N006P009nsss(0)='1'  )then
          oVar1S273(0) <='1';
          else
          oVar1S273(0) <='0';
          end if;
        if(cVar2S8S38P037P030nsss(0)='1'  OR cVar2S9S38P037N030P000nsss(0)='1'  OR cVar2S10S38P037P006nsss(0)='1'  OR cVar1S11S38P048N025P052P046nsss(0)='1'  )then
          oVar1S274(0) <='1';
          else
          oVar1S274(0) <='0';
          end if;
        if(cVar2S12S38P009nsss(0)='1'  OR cVar2S13S38P045P043nsss(0)='1'  OR cVar2S14S38P045P022nsss(0)='1'  OR cVar2S15S38P045N022P024nsss(0)='1'  )then
          oVar1S275(0) <='1';
          else
          oVar1S275(0) <='0';
          end if;
        if(cVar2S16S38P016P065P054nsss(0)='1'  OR cVar2S17S38P016N065P031nsss(0)='1'  OR cVar2S18S38N016P036nsss(0)='1'  OR cVar2S19S38N016P036P017nsss(0)='1'  )then
          oVar1S276(0) <='1';
          else
          oVar1S276(0) <='0';
          end if;
        if(cVar2S20S38P018P019nsss(0)='1'  OR cVar2S21S38N018P056nsss(0)='1'  OR cVar2S22S38N018N056P004nsss(0)='1'  OR cVar2S23S38P044nsss(0)='1'  )then
          oVar1S277(0) <='1';
          else
          oVar1S277(0) <='0';
          end if;
        if(cVar2S24S38N044P043nsss(0)='1'  OR cVar2S25S38N044N043P049nsss(0)='1'  OR cVar2S26S38P006nsss(0)='1'  OR cVar2S27S38P009nsss(0)='1'  )then
          oVar1S278(0) <='1';
          else
          oVar1S278(0) <='0';
          end if;
        if(cVar1S0S39P048P025P007nsss(0)='1'  OR cVar1S1S39P048P025N007P004nsss(0)='1'  OR cVar2S2S39P009nsss(0)='1'  OR cVar2S3S39N009P006nsss(0)='1'  )then
          oVar1S280(0) <='1';
          else
          oVar1S280(0) <='0';
          end if;
        if(cVar2S4S39N009N006P005nsss(0)='1'  OR cVar1S5S39P048N025P027P007nsss(0)='1'  OR cVar2S6S39P006nsss(0)='1'  OR cVar2S7S39N006P009P050nsss(0)='1'  )then
          oVar1S281(0) <='1';
          else
          oVar1S281(0) <='0';
          end if;
        if(cVar2S8S39N006N009P008nsss(0)='1'  OR cVar1S9S39P048N025N027P058nsss(0)='1'  OR cVar2S10S39P030nsss(0)='1'  OR cVar2S11S39N030P024P013nsss(0)='1'  )then
          oVar1S282(0) <='1';
          else
          oVar1S282(0) <='0';
          end if;
        if(cVar2S12S39N030N024P045nsss(0)='1'  OR cVar1S13S39N048P044P004nsss(0)='1'  OR cVar2S14S39P023nsss(0)='1'  OR cVar2S15S39N023P046nsss(0)='1'  )then
          oVar1S283(0) <='1';
          else
          oVar1S283(0) <='0';
          end if;
        if(cVar2S16S39P006P024nsss(0)='1'  OR cVar2S17S39P006N024P025nsss(0)='1'  OR cVar2S18S39N006P021nsss(0)='1'  OR cVar2S19S39N006N021P042nsss(0)='1'  )then
          oVar1S284(0) <='1';
          else
          oVar1S284(0) <='0';
          end if;
        if(cVar2S20S39P067P015nsss(0)='1'  OR cVar2S21S39P067N015P029nsss(0)='1'  OR cVar2S22S39N067P065nsss(0)='1'  OR cVar2S23S39N067N065P034nsss(0)='1'  )then
          oVar1S285(0) <='1';
          else
          oVar1S285(0) <='0';
          end if;
        if(cVar2S24S39P018P016P034nsss(0)='1'  OR cVar2S25S39P018P016P063nsss(0)='1'  OR cVar2S26S39N018P016P065nsss(0)='1'  OR cVar2S27S39P019P018nsss(0)='1'  )then
          oVar1S286(0) <='1';
          else
          oVar1S286(0) <='0';
          end if;
        if(cVar2S28S39P019N018P013nsss(0)='1'  )then
          oVar1S287(0) <='1';
          else
          oVar1S287(0) <='0';
          end if;
        if(cVar1S0S40P018P048P025nsss(0)='1'  OR cVar2S1S40P009nsss(0)='1'  OR cVar2S2S40N009P006nsss(0)='1'  OR cVar2S3S40N009N006P007nsss(0)='1'  )then
          oVar1S288(0) <='1';
          else
          oVar1S288(0) <='0';
          end if;
        if(cVar2S4S40P058nsss(0)='1'  OR cVar2S5S40N058P024P046nsss(0)='1'  OR cVar2S6S40P059P019P058nsss(0)='1'  OR cVar2S7S40P059P019P066nsss(0)='1'  )then
          oVar1S289(0) <='1';
          else
          oVar1S289(0) <='0';
          end if;
        if(cVar2S8S40N059P060nsss(0)='1'  OR cVar2S9S40N059N060P015nsss(0)='1'  OR cVar2S10S40P035P034P057nsss(0)='1'  OR cVar2S11S40P035P034P009nsss(0)='1'  )then
          oVar1S290(0) <='1';
          else
          oVar1S290(0) <='0';
          end if;
        if(cVar2S12S40N035P011nsss(0)='1'  OR cVar2S13S40N035N011P029nsss(0)='1'  OR cVar2S14S40P055nsss(0)='1'  OR cVar2S15S40N055P054nsss(0)='1'  )then
          oVar1S291(0) <='1';
          else
          oVar1S291(0) <='0';
          end if;
        if(cVar2S16S40N055N054P051nsss(0)='1'  OR cVar2S17S40P030P057nsss(0)='1'  OR cVar2S18S40P030N057P056nsss(0)='1'  OR cVar2S19S40N030P029P037nsss(0)='1'  )then
          oVar1S292(0) <='1';
          else
          oVar1S292(0) <='0';
          end if;
        if(cVar2S20S40P028P057P000nsss(0)='1'  OR cVar2S21S40P007nsss(0)='1'  OR cVar2S22S40N007P017P037nsss(0)='1'  OR cVar2S23S40P066P064nsss(0)='1'  )then
          oVar1S293(0) <='1';
          else
          oVar1S293(0) <='0';
          end if;
        if(cVar2S24S40P066P016P017nsss(0)='1'  OR cVar2S25S40P015P019P066nsss(0)='1'  OR cVar2S26S40P015P019P007nsss(0)='1'  OR cVar2S27S40P015P012nsss(0)='1'  )then
          oVar1S294(0) <='1';
          else
          oVar1S294(0) <='0';
          end if;
        if(cVar2S28S40P015N012P064nsss(0)='1'  OR cVar1S29S40P018P069P052P029nsss(0)='1'  )then
          oVar1S295(0) <='1';
          else
          oVar1S295(0) <='0';
          end if;
        if(cVar1S0S41P048P025P007nsss(0)='1'  OR cVar1S1S41P048P025N007P004nsss(0)='1'  OR cVar2S2S41P009nsss(0)='1'  OR cVar2S3S41N009P006nsss(0)='1'  )then
          oVar1S296(0) <='1';
          else
          oVar1S296(0) <='0';
          end if;
        if(cVar2S4S41N009N006P005nsss(0)='1'  OR cVar2S5S41P050P027nsss(0)='1'  OR cVar2S6S41P050N027P011nsss(0)='1'  OR cVar2S7S41N050P005P017nsss(0)='1'  )then
          oVar1S297(0) <='1';
          else
          oVar1S297(0) <='0';
          end if;
        if(cVar2S8S41P046nsss(0)='1'  OR cVar1S9S41P048N025P052P015nsss(0)='1'  OR cVar2S10S41P054nsss(0)='1'  OR cVar2S11S41N054P046nsss(0)='1'  )then
          oVar1S298(0) <='1';
          else
          oVar1S298(0) <='0';
          end if;
        if(cVar2S12S41P043P025P022nsss(0)='1'  OR cVar2S13S41P043P025P017nsss(0)='1'  OR cVar2S14S41P043P019P041nsss(0)='1'  OR cVar2S15S41P022nsss(0)='1'  )then
          oVar1S299(0) <='1';
          else
          oVar1S299(0) <='0';
          end if;
        if(cVar2S16S41N022P007nsss(0)='1'  OR cVar2S17S41N022N007P005nsss(0)='1'  OR cVar1S18S41N048P018P059P050nsss(0)='1'  OR cVar2S19S41P004P061P009nsss(0)='1'  )then
          oVar1S300(0) <='1';
          else
          oVar1S300(0) <='0';
          end if;
        if(cVar2S20S41P004N061P057nsss(0)='1'  OR cVar2S21S41P065P014nsss(0)='1'  OR cVar2S22S41P065N014P012nsss(0)='1'  OR cVar2S23S41P065P037nsss(0)='1'  )then
          oVar1S301(0) <='1';
          else
          oVar1S301(0) <='0';
          end if;
        if(cVar2S24S41P013P031nsss(0)='1'  OR cVar2S25S41P013N031P010nsss(0)='1'  OR cVar2S26S41N013P011nsss(0)='1'  OR cVar2S27S41N013N011P010nsss(0)='1'  )then
          oVar1S302(0) <='1';
          else
          oVar1S302(0) <='0';
          end if;
        if(cVar2S28S41P035P012P017nsss(0)='1'  OR cVar2S29S41P035P012P014nsss(0)='1'  OR cVar2S30S41N035P024P006nsss(0)='1'  )then
          oVar1S303(0) <='1';
          else
          oVar1S303(0) <='0';
          end if;
        if(cVar1S0S42P018P048P025nsss(0)='1'  OR cVar2S1S42P009nsss(0)='1'  OR cVar2S2S42N009P006nsss(0)='1'  OR cVar2S3S42N009N006P008nsss(0)='1'  )then
          oVar1S304(0) <='1';
          else
          oVar1S304(0) <='0';
          end if;
        if(cVar2S4S42P062P066nsss(0)='1'  OR cVar2S5S42N062P006nsss(0)='1'  OR cVar2S6S42N062N006P040nsss(0)='1'  OR cVar1S7S42P018N048P038P002nsss(0)='1'  )then
          oVar1S305(0) <='1';
          else
          oVar1S305(0) <='0';
          end if;
        if(cVar2S8S42P015P021nsss(0)='1'  OR cVar2S9S42P015N021P004nsss(0)='1'  OR cVar2S10S42P022P043P010nsss(0)='1'  OR cVar2S11S42P022N043P007nsss(0)='1'  )then
          oVar1S306(0) <='1';
          else
          oVar1S306(0) <='0';
          end if;
        if(cVar2S12S42N022P046P005nsss(0)='1'  OR cVar2S13S42N022P046P025nsss(0)='1'  OR cVar2S14S42P047P063P062nsss(0)='1'  OR cVar2S15S42P014nsss(0)='1'  )then
          oVar1S307(0) <='1';
          else
          oVar1S307(0) <='0';
          end if;
        if(cVar2S16S42N014P017nsss(0)='1'  OR cVar2S17S42N014P017P046nsss(0)='1'  OR cVar2S18S42P016nsss(0)='1'  OR cVar2S19S42P017nsss(0)='1'  )then
          oVar1S308(0) <='1';
          else
          oVar1S308(0) <='0';
          end if;
        if(cVar1S20S42P018N048P044P023nsss(0)='1'  OR cVar2S21S42P046nsss(0)='1'  OR cVar2S22S42N046P015nsss(0)='1'  OR cVar2S23S42P042P023P067nsss(0)='1'  )then
          oVar1S309(0) <='1';
          else
          oVar1S309(0) <='0';
          end if;
        if(cVar2S24S42P042P066P013nsss(0)='1'  OR cVar2S25S42P017P019P012nsss(0)='1'  OR cVar2S26S42N017P041nsss(0)='1'  OR cVar2S27S42N017N041P009nsss(0)='1'  )then
          oVar1S310(0) <='1';
          else
          oVar1S310(0) <='0';
          end if;
        if(cVar1S0S43P048P025P007nsss(0)='1'  OR cVar1S1S43P048P025N007P004nsss(0)='1'  OR cVar2S2S43P009nsss(0)='1'  OR cVar2S3S43N009P006nsss(0)='1'  )then
          oVar1S312(0) <='1';
          else
          oVar1S312(0) <='0';
          end if;
        if(cVar2S4S43N009N006P008nsss(0)='1'  OR cVar1S5S43P048N025P062P058nsss(0)='1'  OR cVar2S6S43P037nsss(0)='1'  OR cVar2S7S43P007nsss(0)='1'  )then
          oVar1S313(0) <='1';
          else
          oVar1S313(0) <='0';
          end if;
        if(cVar2S8S43N007P006nsss(0)='1'  OR cVar2S9S43N007N006P009nsss(0)='1'  OR cVar2S10S43P045nsss(0)='1'  OR cVar2S11S43N045P000nsss(0)='1'  )then
          oVar1S314(0) <='1';
          else
          oVar1S314(0) <='0';
          end if;
        if(cVar2S12S43P010nsss(0)='1'  OR cVar2S13S43P042nsss(0)='1'  OR cVar2S14S43P049P067P036nsss(0)='1'  OR cVar2S15S43P002nsss(0)='1'  )then
          oVar1S315(0) <='1';
          else
          oVar1S315(0) <='0';
          end if;
        if(cVar2S16S43N002P015nsss(0)='1'  OR cVar2S17S43P041nsss(0)='1'  OR cVar2S18S43N041P067P003nsss(0)='1'  OR cVar2S19S43P008P049nsss(0)='1'  )then
          oVar1S316(0) <='1';
          else
          oVar1S316(0) <='0';
          end if;
        if(cVar2S20S43P008N049P051nsss(0)='1'  OR cVar2S21S43N008P030P012nsss(0)='1'  OR cVar2S22S43P042nsss(0)='1'  OR cVar2S23S43N042P017P012nsss(0)='1'  )then
          oVar1S317(0) <='1';
          else
          oVar1S317(0) <='0';
          end if;
        if(cVar2S24S43N042N017P045nsss(0)='1'  )then
          oVar1S318(0) <='1';
          else
          oVar1S318(0) <='0';
          end if;
        if(cVar1S0S44P022P043P037P010nsss(0)='1'  OR cVar1S1S44P022P043P037P004nsss(0)='1'  OR cVar1S2S44P022N043P004nsss(0)='1'  OR cVar2S3S44P067P017nsss(0)='1'  )then
          oVar1S319(0) <='1';
          else
          oVar1S319(0) <='0';
          end if;
        if(cVar2S4S44P008nsss(0)='1'  OR cVar2S5S44N008P047P006nsss(0)='1'  OR cVar2S6S44N008P047P006nsss(0)='1'  OR cVar2S7S44P047P006nsss(0)='1'  )then
          oVar1S320(0) <='1';
          else
          oVar1S320(0) <='0';
          end if;
        if(cVar2S8S44P047N006P017nsss(0)='1'  OR cVar2S9S44N047P051nsss(0)='1'  OR cVar2S10S44N047N051P044nsss(0)='1'  OR cVar2S11S44P005nsss(0)='1'  )then
          oVar1S321(0) <='1';
          else
          oVar1S321(0) <='0';
          end if;
        if(cVar2S12S44N005P044nsss(0)='1'  OR cVar2S13S44P006nsss(0)='1'  OR cVar2S14S44N006P007nsss(0)='1'  OR cVar2S15S44N006N007P003nsss(0)='1'  )then
          oVar1S322(0) <='1';
          else
          oVar1S322(0) <='0';
          end if;
        if(cVar1S16S44N022P004P040nsss(0)='1'  OR cVar2S17S44P012P048nsss(0)='1'  OR cVar2S18S44P012N048P016nsss(0)='1'  OR cVar2S19S44P044P023nsss(0)='1'  )then
          oVar1S323(0) <='1';
          else
          oVar1S323(0) <='0';
          end if;
        if(cVar2S20S44N044P015P002nsss(0)='1'  OR cVar2S21S44N044N015P045nsss(0)='1'  )then
          oVar1S324(0) <='1';
          else
          oVar1S324(0) <='0';
          end if;
        if(cVar1S0S45P022P043P019nsss(0)='1'  OR cVar2S1S45P013nsss(0)='1'  OR cVar1S2S45P022N043P004P042nsss(0)='1'  OR cVar1S3S45P022N043N004P007nsss(0)='1'  )then
          oVar1S325(0) <='1';
          else
          oVar1S325(0) <='0';
          end if;
        if(cVar2S4S45P033nsss(0)='1'  OR cVar2S5S45N033P002nsss(0)='1'  OR cVar2S6S45N033N002P008nsss(0)='1'  OR cVar1S7S45N022P047P006nsss(0)='1'  )then
          oVar1S326(0) <='1';
          else
          oVar1S326(0) <='0';
          end if;
        if(cVar2S8S45P026P018nsss(0)='1'  OR cVar2S9S45P026N018P050nsss(0)='1'  OR cVar2S10S45N026P024nsss(0)='1'  OR cVar2S11S45P007P015nsss(0)='1'  )then
          oVar1S327(0) <='1';
          else
          oVar1S327(0) <='0';
          end if;
        if(cVar2S12S45N007P009P051nsss(0)='1'  OR cVar2S13S45N007N009P069nsss(0)='1'  OR cVar2S14S45P028nsss(0)='1'  OR cVar2S15S45N028P026P066nsss(0)='1'  )then
          oVar1S328(0) <='1';
          else
          oVar1S328(0) <='0';
          end if;
        if(cVar2S16S45N028N026P053nsss(0)='1'  OR cVar2S17S45P027P009nsss(0)='1'  OR cVar2S18S45P027N009P011nsss(0)='1'  OR cVar2S19S45N027P011nsss(0)='1'  )then
          oVar1S329(0) <='1';
          else
          oVar1S329(0) <='0';
          end if;
        if(cVar2S20S45P023P005P068nsss(0)='1'  OR cVar2S21S45P023N005P004nsss(0)='1'  OR cVar2S22S45N023P043P024nsss(0)='1'  OR cVar2S23S45P033nsss(0)='1'  )then
          oVar1S330(0) <='1';
          else
          oVar1S330(0) <='0';
          end if;
        if(cVar2S24S45N033P034nsss(0)='1'  )then
          oVar1S331(0) <='1';
          else
          oVar1S331(0) <='0';
          end if;
        if(cVar1S0S46P022P043P019nsss(0)='1'  OR cVar1S1S46P022P043N019P037nsss(0)='1'  OR cVar1S2S46P022N043P004nsss(0)='1'  OR cVar2S3S46P061nsss(0)='1'  )then
          oVar1S332(0) <='1';
          else
          oVar1S332(0) <='0';
          end if;
        if(cVar2S4S46N061P069P003nsss(0)='1'  OR cVar2S5S46P067nsss(0)='1'  OR cVar2S6S46P045nsss(0)='1'  OR cVar2S7S46N045P052nsss(0)='1'  )then
          oVar1S333(0) <='1';
          else
          oVar1S333(0) <='0';
          end if;
        if(cVar2S8S46N045P052P015nsss(0)='1'  OR cVar2S9S46P025P059P027nsss(0)='1'  OR cVar2S10S46P025P059P003nsss(0)='1'  OR cVar2S11S46P025P014nsss(0)='1'  )then
          oVar1S334(0) <='1';
          else
          oVar1S334(0) <='0';
          end if;
        if(cVar2S12S46P062P069P067nsss(0)='1'  OR cVar2S13S46P062N069P068nsss(0)='1'  OR cVar2S14S46P005P039nsss(0)='1'  OR cVar2S15S46N005P004nsss(0)='1'  )then
          oVar1S335(0) <='1';
          else
          oVar1S335(0) <='0';
          end if;
        if(cVar2S16S46N005N004P006nsss(0)='1'  OR cVar2S17S46P043P045nsss(0)='1'  OR cVar2S18S46P043P045P024nsss(0)='1'  OR cVar2S19S46P043P006nsss(0)='1'  )then
          oVar1S336(0) <='1';
          else
          oVar1S336(0) <='0';
          end if;
        if(cVar2S20S46P043N006P007nsss(0)='1'  )then
          oVar1S337(0) <='1';
          else
          oVar1S337(0) <='0';
          end if;
        if(cVar1S0S47P022P043P019nsss(0)='1'  OR cVar2S1S47P004nsss(0)='1'  OR cVar2S2S47N004P005nsss(0)='1'  OR cVar2S3S47N004N005P007nsss(0)='1'  )then
          oVar1S338(0) <='1';
          else
          oVar1S338(0) <='0';
          end if;
        if(cVar1S4S47P022N043P004P042nsss(0)='1'  OR cVar2S5S47P061nsss(0)='1'  OR cVar2S6S47N061P067P036nsss(0)='1'  OR cVar2S7S47P043nsss(0)='1'  )then
          oVar1S339(0) <='1';
          else
          oVar1S339(0) <='0';
          end if;
        if(cVar2S8S47N043P042nsss(0)='1'  OR cVar2S9S47P007nsss(0)='1'  OR cVar2S10S47N007P004nsss(0)='1'  OR cVar2S11S47N007N004P006nsss(0)='1'  )then
          oVar1S340(0) <='1';
          else
          oVar1S340(0) <='0';
          end if;
        if(cVar2S12S47P025P050P067nsss(0)='1'  OR cVar2S13S47N025P045nsss(0)='1'  OR cVar2S14S47N025N045P036nsss(0)='1'  OR cVar2S15S47P045P037P025nsss(0)='1'  )then
          oVar1S341(0) <='1';
          else
          oVar1S341(0) <='0';
          end if;
        if(cVar2S16S47P045N037P016nsss(0)='1'  OR cVar2S17S47P045P047nsss(0)='1'  OR cVar2S18S47P045N047P060nsss(0)='1'  OR cVar1S19S47N022N023P043P006nsss(0)='1'  )then
          oVar1S342(0) <='1';
          else
          oVar1S342(0) <='0';
          end if;
        if(cVar2S20S47P007P025nsss(0)='1'  OR cVar2S21S47P007N025P024nsss(0)='1'  OR cVar2S22S47N007P059nsss(0)='1'  OR cVar2S23S47N007N059P020nsss(0)='1'  )then
          oVar1S343(0) <='1';
          else
          oVar1S343(0) <='0';
          end if;
        if(cVar2S0S48P055P056P060nsss(0)='1'  OR cVar2S1S48P055P017nsss(0)='1'  OR cVar2S2S48P023P005nsss(0)='1'  OR cVar2S3S48P023N005P042nsss(0)='1'  )then
          oVar1S345(0) <='1';
          else
          oVar1S345(0) <='0';
          end if;
        if(cVar2S4S48N023P028P010nsss(0)='1'  OR cVar2S5S48N023N028psss(0)='1'  OR cVar2S6S48P062nsss(0)='1'  OR cVar2S7S48N062P059P032nsss(0)='1'  )then
          oVar1S346(0) <='1';
          else
          oVar1S346(0) <='0';
          end if;
        if(cVar2S8S48N062N059P037nsss(0)='1'  OR cVar2S9S48P064P002nsss(0)='1'  OR cVar1S10S48P016P065P067P063nsss(0)='1'  OR cVar2S11S48P035P018nsss(0)='1'  )then
          oVar1S347(0) <='1';
          else
          oVar1S347(0) <='0';
          end if;
        if(cVar2S12S48N035P062P034nsss(0)='1'  OR cVar2S13S48P034P014P015nsss(0)='1'  OR cVar2S14S48P034N014P017nsss(0)='1'  OR cVar2S15S48N034P035P063nsss(0)='1'  )then
          oVar1S348(0) <='1';
          else
          oVar1S348(0) <='0';
          end if;
        if(cVar2S16S48P015P018nsss(0)='1'  OR cVar2S17S48N015P012P014nsss(0)='1'  OR cVar2S18S48P066P032nsss(0)='1'  OR cVar2S19S48P066P018P036nsss(0)='1'  )then
          oVar1S349(0) <='1';
          else
          oVar1S349(0) <='0';
          end if;
        if(cVar2S20S48P066N018P067nsss(0)='1'  OR cVar2S21S48P018P062nsss(0)='1'  OR cVar2S22S48P018N062P066nsss(0)='1'  OR cVar2S23S48P018P013P019nsss(0)='1'  )then
          oVar1S350(0) <='1';
          else
          oVar1S350(0) <='0';
          end if;
        if(cVar2S24S48P004P022nsss(0)='1'  OR cVar2S25S48P004N022P019nsss(0)='1'  OR cVar2S26S48N004P062P055nsss(0)='1'  OR cVar2S27S48P018P015P014nsss(0)='1'  )then
          oVar1S351(0) <='1';
          else
          oVar1S351(0) <='0';
          end if;
        if(cVar2S28S48P018N015P014nsss(0)='1'  OR cVar2S29S48N018P032P015nsss(0)='1'  OR cVar2S30S48P029P017nsss(0)='1'  OR cVar2S31S48P029N017P009nsss(0)='1'  )then
          oVar1S352(0) <='1';
          else
          oVar1S352(0) <='0';
          end if;
        if(cVar1S0S49P023P005P042nsss(0)='1'  OR cVar1S1S49P023P005N042P043nsss(0)='1'  OR cVar2S2S49P043nsss(0)='1'  OR cVar2S3S49N043P044nsss(0)='1'  )then
          oVar1S354(0) <='1';
          else
          oVar1S354(0) <='0';
          end if;
        if(cVar2S4S49P054nsss(0)='1'  OR cVar2S5S49N054P004P044nsss(0)='1'  OR cVar2S6S49N054N004P003nsss(0)='1'  OR cVar1S7S49N023P022P043P005nsss(0)='1'  )then
          oVar1S355(0) <='1';
          else
          oVar1S355(0) <='0';
          end if;
        if(cVar2S8S49P019nsss(0)='1'  OR cVar2S9S49N019P004P018nsss(0)='1'  OR cVar2S10S49N019N004P007nsss(0)='1'  OR cVar1S11S49N023P022N043P004nsss(0)='1'  )then
          oVar1S356(0) <='1';
          else
          oVar1S356(0) <='0';
          end if;
        if(cVar2S12S49P007nsss(0)='1'  OR cVar2S13S49N007P002nsss(0)='1'  OR cVar2S14S49N007N002P018nsss(0)='1'  OR cVar2S15S49P034P063P036nsss(0)='1'  )then
          oVar1S357(0) <='1';
          else
          oVar1S357(0) <='0';
          end if;
        if(cVar2S16S49P034N063P062nsss(0)='1'  OR cVar2S17S49N034P036P037nsss(0)='1'  OR cVar2S18S49P051nsss(0)='1'  OR cVar2S19S49P010P055P012nsss(0)='1'  )then
          oVar1S358(0) <='1';
          else
          oVar1S358(0) <='0';
          end if;
        if(cVar2S20S49P010N055P051nsss(0)='1'  OR cVar2S21S49N010P029P008nsss(0)='1'  OR cVar2S22S49P059P032P035nsss(0)='1'  OR cVar2S23S49P059N032P013nsss(0)='1'  )then
          oVar1S359(0) <='1';
          else
          oVar1S359(0) <='0';
          end if;
        if(cVar2S24S49N059P047P006nsss(0)='1'  )then
          oVar1S360(0) <='1';
          else
          oVar1S360(0) <='0';
          end if;
        if(cVar1S0S50P023P005P042nsss(0)='1'  OR cVar1S1S50P023P005N042P043nsss(0)='1'  OR cVar2S2S50P043nsss(0)='1'  OR cVar2S3S50N043P018nsss(0)='1'  )then
          oVar1S361(0) <='1';
          else
          oVar1S361(0) <='0';
          end if;
        if(cVar2S4S50P064nsss(0)='1'  OR cVar2S5S50N064P006nsss(0)='1'  OR cVar2S6S50P031nsss(0)='1'  OR cVar2S7S50P008P014nsss(0)='1'  )then
          oVar1S362(0) <='1';
          else
          oVar1S362(0) <='0';
          end if;
        if(cVar2S8S50N008P063P011nsss(0)='1'  OR cVar2S9S50P007nsss(0)='1'  OR cVar2S10S50N007P046nsss(0)='1'  OR cVar2S11S50P024P006P011nsss(0)='1'  )then
          oVar1S363(0) <='1';
          else
          oVar1S363(0) <='0';
          end if;
        if(cVar2S12S50P024N006P010nsss(0)='1'  OR cVar2S13S50N024P045P043nsss(0)='1'  OR cVar2S14S50N024P045P022nsss(0)='1'  OR cVar2S15S50P011nsss(0)='1'  )then
          oVar1S364(0) <='1';
          else
          oVar1S364(0) <='0';
          end if;
        if(cVar2S16S50N011P009nsss(0)='1'  OR cVar2S17S50P026P036P011nsss(0)='1'  OR cVar2S18S50N026P027nsss(0)='1'  OR cVar2S19S50N026N027P035nsss(0)='1'  )then
          oVar1S365(0) <='1';
          else
          oVar1S365(0) <='0';
          end if;
        if(cVar2S0S51P053nsss(0)='1'  OR cVar2S1S51N053P055P012nsss(0)='1'  OR cVar2S2S51N053N055P054nsss(0)='1'  OR cVar1S3S51P028P029N010P008nsss(0)='1'  )then
          oVar1S367(0) <='1';
          else
          oVar1S367(0) <='0';
          end if;
        if(cVar2S4S51P063P068P014nsss(0)='1'  OR cVar1S5S51N028P023P005P042nsss(0)='1'  OR cVar2S6S51P043nsss(0)='1'  OR cVar2S7S51P026P007P015nsss(0)='1'  )then
          oVar1S368(0) <='1';
          else
          oVar1S368(0) <='0';
          end if;
        if(cVar2S8S51P026N007psss(0)='1'  OR cVar1S9S51N028N023P025P007nsss(0)='1'  OR cVar2S10S51P046nsss(0)='1'  OR cVar2S11S51N046P003P057nsss(0)='1'  )then
          oVar1S369(0) <='1';
          else
          oVar1S369(0) <='0';
          end if;
        if(cVar2S12S51P006P047nsss(0)='1'  OR cVar2S13S51P006N047P043nsss(0)='1'  OR cVar2S14S51N006P047nsss(0)='1'  OR cVar2S15S51P041P020nsss(0)='1'  )then
          oVar1S370(0) <='1';
          else
          oVar1S370(0) <='0';
          end if;
        if(cVar2S16S51P041N020P001nsss(0)='1'  OR cVar2S17S51N041P039P064nsss(0)='1'  )then
          oVar1S371(0) <='1';
          else
          oVar1S371(0) <='0';
          end if;
        if(cVar1S0S52P045P043P005P068nsss(0)='1'  OR cVar1S1S52P045P043N005P004nsss(0)='1'  OR cVar2S2S52P006nsss(0)='1'  OR cVar2S3S52N006P007P015nsss(0)='1'  )then
          oVar1S372(0) <='1';
          else
          oVar1S372(0) <='0';
          end if;
        if(cVar2S4S52N006N007P003nsss(0)='1'  OR cVar1S5S52P045N043P047P006nsss(0)='1'  OR cVar2S6S52P024nsss(0)='1'  OR cVar2S7S52N024P016nsss(0)='1'  )then
          oVar1S373(0) <='1';
          else
          oVar1S373(0) <='0';
          end if;
        if(cVar1S8S52P045N043N047P048nsss(0)='1'  OR cVar2S9S52P060nsss(0)='1'  OR cVar2S10S52N060P044nsss(0)='1'  OR cVar2S11S52N060N044P063nsss(0)='1'  )then
          oVar1S374(0) <='1';
          else
          oVar1S374(0) <='0';
          end if;
        if(cVar2S12S52P012nsss(0)='1'  OR cVar2S13S52P034P054nsss(0)='1'  OR cVar2S14S52P034N054P053nsss(0)='1'  OR cVar2S15S52P053nsss(0)='1'  )then
          oVar1S375(0) <='1';
          else
          oVar1S375(0) <='0';
          end if;
        if(cVar2S16S52N053P057nsss(0)='1'  OR cVar2S17S52N053N057P016nsss(0)='1'  OR cVar2S18S52P029P008nsss(0)='1'  OR cVar2S19S52P029N008P012nsss(0)='1'  )then
          oVar1S376(0) <='1';
          else
          oVar1S376(0) <='0';
          end if;
        if(cVar2S20S52P002nsss(0)='1'  OR cVar2S21S52N002P016P017nsss(0)='1'  OR cVar2S22S52P020nsss(0)='1'  OR cVar2S23S52N020P066P050nsss(0)='1'  )then
          oVar1S377(0) <='1';
          else
          oVar1S377(0) <='0';
          end if;
        if(cVar2S24S52P046P066nsss(0)='1'  OR cVar2S25S52P046P066P018nsss(0)='1'  OR cVar2S26S52N046P007P047nsss(0)='1'  OR cVar2S27S52P015P056nsss(0)='1'  )then
          oVar1S378(0) <='1';
          else
          oVar1S378(0) <='0';
          end if;
        if(cVar2S28S52P015P056P068nsss(0)='1'  OR cVar2S29S52N015P005nsss(0)='1'  OR cVar2S30S52N015P005P023nsss(0)='1'  )then
          oVar1S379(0) <='1';
          else
          oVar1S379(0) <='0';
          end if;
        if(cVar1S0S53P025P007P066nsss(0)='1'  OR cVar1S1S53P025P007P066P037nsss(0)='1'  OR cVar1S2S53P025N007P046P004nsss(0)='1'  OR cVar2S3S53P006nsss(0)='1'  )then
          oVar1S380(0) <='1';
          else
          oVar1S380(0) <='0';
          end if;
        if(cVar2S4S53N006P048nsss(0)='1'  OR cVar2S5S53P057nsss(0)='1'  OR cVar2S6S53N057P037P034nsss(0)='1'  OR cVar1S7S53N025P028P010P055nsss(0)='1'  )then
          oVar1S381(0) <='1';
          else
          oVar1S381(0) <='0';
          end if;
        if(cVar2S8S53P005P017nsss(0)='1'  OR cVar2S9S53P005N017P026nsss(0)='1'  OR cVar2S10S53P063P053P014nsss(0)='1'  OR cVar2S11S53P063N053P012nsss(0)='1'  )then
          oVar1S382(0) <='1';
          else
          oVar1S382(0) <='0';
          end if;
        if(cVar2S12S53P011nsss(0)='1'  OR cVar2S13S53P002nsss(0)='1'  OR cVar2S14S53N002P015nsss(0)='1'  OR cVar2S15S53P066P020nsss(0)='1'  )then
          oVar1S383(0) <='1';
          else
          oVar1S383(0) <='0';
          end if;
        if(cVar2S16S53P066N020P047nsss(0)='1'  OR cVar2S17S53P022nsss(0)='1'  OR cVar2S18S53N022P024nsss(0)='1'  OR cVar2S19S53N022N024P023nsss(0)='1'  )then
          oVar1S384(0) <='1';
          else
          oVar1S384(0) <='0';
          end if;
        if(cVar2S20S53P015P047P060nsss(0)='1'  OR cVar2S21S53P015P047P026nsss(0)='1'  OR cVar2S22S53N015P018P004nsss(0)='1'  OR cVar2S23S53N015N018P016nsss(0)='1'  )then
          oVar1S385(0) <='1';
          else
          oVar1S385(0) <='0';
          end if;
        if(cVar1S0S54P018P040P002nsss(0)='1'  OR cVar1S1S54P018P040N002P004nsss(0)='1'  OR cVar2S2S54P003P014nsss(0)='1'  OR cVar2S3S54N003P005nsss(0)='1'  )then
          oVar1S387(0) <='1';
          else
          oVar1S387(0) <='0';
          end if;
        if(cVar2S4S54N003N005P050nsss(0)='1'  OR cVar1S5S54P018N040P045P004nsss(0)='1'  OR cVar2S6S54P023nsss(0)='1'  OR cVar2S7S54N023P006nsss(0)='1'  )then
          oVar1S388(0) <='1';
          else
          oVar1S388(0) <='0';
          end if;
        if(cVar2S8S54N023N006P007nsss(0)='1'  OR cVar2S9S54P036P047nsss(0)='1'  OR cVar2S10S54P036P009P019nsss(0)='1'  OR cVar2S11S54P028P029nsss(0)='1'  )then
          oVar1S389(0) <='1';
          else
          oVar1S389(0) <='0';
          end if;
        if(cVar2S12S54N028P025nsss(0)='1'  OR cVar2S13S54N028N025P016nsss(0)='1'  OR cVar2S14S54P027nsss(0)='1'  OR cVar2S15S54N027P045nsss(0)='1'  )then
          oVar1S390(0) <='1';
          else
          oVar1S390(0) <='0';
          end if;
        if(cVar2S16S54N027N045P023nsss(0)='1'  OR cVar2S17S54P012nsss(0)='1'  OR cVar1S18S54P018P015N019P053nsss(0)='1'  OR cVar2S19S54P006P066P069nsss(0)='1'  )then
          oVar1S391(0) <='1';
          else
          oVar1S391(0) <='0';
          end if;
        if(cVar2S20S54N006P033P067nsss(0)='1'  OR cVar2S21S54P025nsss(0)='1'  OR cVar2S22S54N025P034P012nsss(0)='1'  OR cVar2S23S54P013nsss(0)='1'  )then
          oVar1S392(0) <='1';
          else
          oVar1S392(0) <='0';
          end if;
        if(cVar2S24S54N013P014nsss(0)='1'  OR cVar2S25S54P007P011P066nsss(0)='1'  OR cVar2S26S54N007P021nsss(0)='1'  )then
          oVar1S393(0) <='1';
          else
          oVar1S393(0) <='0';
          end if;
        if(cVar1S0S55P040P002nsss(0)='1'  OR cVar2S1S55P003nsss(0)='1'  OR cVar2S2S55N003P005P038nsss(0)='1'  OR cVar2S3S55P004nsss(0)='1'  )then
          oVar1S394(0) <='1';
          else
          oVar1S394(0) <='0';
          end if;
        if(cVar2S4S55N004P050nsss(0)='1'  OR cVar2S5S55N004N050P068nsss(0)='1'  OR cVar1S6S55P040N002P015P013nsss(0)='1'  OR cVar2S7S55P019nsss(0)='1'  )then
          oVar1S395(0) <='1';
          else
          oVar1S395(0) <='0';
          end if;
        if(cVar2S8S55P012nsss(0)='1'  OR cVar2S9S55P013P022nsss(0)='1'  OR cVar2S10S55P013N022P043nsss(0)='1'  OR cVar2S11S55P006P024nsss(0)='1'  )then
          oVar1S396(0) <='1';
          else
          oVar1S396(0) <='0';
          end if;
        if(cVar2S12S55P006N024P022nsss(0)='1'  OR cVar2S13S55N006P007P068nsss(0)='1'  OR cVar2S14S55N006N007P051nsss(0)='1'  OR cVar2S15S55P042P032P033nsss(0)='1'  )then
          oVar1S397(0) <='1';
          else
          oVar1S397(0) <='0';
          end if;
        if(cVar2S16S55P042N032psss(0)='1'  OR cVar2S17S55P042P016P044nsss(0)='1'  OR cVar2S18S55P042N016P023nsss(0)='1'  OR cVar2S19S55P033P049P037nsss(0)='1'  )then
          oVar1S398(0) <='1';
          else
          oVar1S398(0) <='0';
          end if;
        if(cVar2S20S55P029P031nsss(0)='1'  OR cVar2S21S55P029P011nsss(0)='1'  OR cVar2S22S55P025P046P066nsss(0)='1'  OR cVar2S23S55P025N046P007nsss(0)='1'  )then
          oVar1S399(0) <='1';
          else
          oVar1S399(0) <='0';
          end if;
        if(cVar2S24S55N025P018P019nsss(0)='1'  OR cVar2S25S55N025N018P011nsss(0)='1'  )then
          oVar1S400(0) <='1';
          else
          oVar1S400(0) <='0';
          end if;
        if(cVar1S0S56P045P005P068P012nsss(0)='1'  OR cVar1S1S56P045N005P004P013nsss(0)='1'  OR cVar2S2S56P024nsss(0)='1'  OR cVar2S3S56N024P022nsss(0)='1'  )then
          oVar1S401(0) <='1';
          else
          oVar1S401(0) <='0';
          end if;
        if(cVar2S4S56P007P068nsss(0)='1'  OR cVar2S5S56N007P003P043nsss(0)='1'  OR cVar2S6S56N007N003P048nsss(0)='1'  OR cVar1S7S56N045P040P021P002nsss(0)='1'  )then
          oVar1S402(0) <='1';
          else
          oVar1S402(0) <='0';
          end if;
        if(cVar2S8S56P015P016nsss(0)='1'  OR cVar2S9S56P020nsss(0)='1'  OR cVar2S10S56N020P008nsss(0)='1'  OR cVar2S11S56P015P003nsss(0)='1'  )then
          oVar1S403(0) <='1';
          else
          oVar1S403(0) <='0';
          end if;
        if(cVar2S12S56P015P003P039nsss(0)='1'  OR cVar2S13S56P015P016P035nsss(0)='1'  OR cVar2S14S56P041nsss(0)='1'  OR cVar2S15S56N041P011nsss(0)='1'  )then
          oVar1S404(0) <='1';
          else
          oVar1S404(0) <='0';
          end if;
        if(cVar2S16S56N041N011P049nsss(0)='1'  OR cVar2S17S56P011P029P013nsss(0)='1'  OR cVar2S18S56P011P029P052nsss(0)='1'  OR cVar2S19S56P011N029P003nsss(0)='1'  )then
          oVar1S405(0) <='1';
          else
          oVar1S405(0) <='0';
          end if;
        if(cVar2S20S56P026P035P058nsss(0)='1'  OR cVar2S21S56P026N035P013nsss(0)='1'  )then
          oVar1S406(0) <='1';
          else
          oVar1S406(0) <='0';
          end if;
        if(cVar1S0S57P045P005P037nsss(0)='1'  OR cVar1S1S57P045N005P004P013nsss(0)='1'  OR cVar2S2S57P024nsss(0)='1'  OR cVar2S3S57N024P022nsss(0)='1'  )then
          oVar1S407(0) <='1';
          else
          oVar1S407(0) <='0';
          end if;
        if(cVar2S4S57P007P068nsss(0)='1'  OR cVar2S5S57N007P014P043nsss(0)='1'  OR cVar2S6S57N007N014P051nsss(0)='1'  OR cVar1S7S57N045P040P021P002nsss(0)='1'  )then
          oVar1S408(0) <='1';
          else
          oVar1S408(0) <='0';
          end if;
        if(cVar2S8S57P003nsss(0)='1'  OR cVar2S9S57N003P004nsss(0)='1'  OR cVar2S10S57N003N004P005nsss(0)='1'  OR cVar2S11S57P002nsss(0)='1'  )then
          oVar1S409(0) <='1';
          else
          oVar1S409(0) <='0';
          end if;
        if(cVar2S12S57P008P060nsss(0)='1'  OR cVar2S13S57P008N060P023nsss(0)='1'  OR cVar2S14S57P011P029P042nsss(0)='1'  OR cVar2S15S57P011P029P013nsss(0)='1'  )then
          oVar1S410(0) <='1';
          else
          oVar1S410(0) <='0';
          end if;
        if(cVar2S16S57P011P053nsss(0)='1'  OR cVar2S17S57P011N053P054nsss(0)='1'  OR cVar2S18S57P001P017P003nsss(0)='1'  OR cVar2S19S57P001N017P016nsss(0)='1'  )then
          oVar1S411(0) <='1';
          else
          oVar1S411(0) <='0';
          end if;
        if(cVar2S20S57P008P049nsss(0)='1'  OR cVar2S21S57P008N049P064nsss(0)='1'  OR cVar2S22S57N008P021P003nsss(0)='1'  OR cVar2S23S57P041nsss(0)='1'  )then
          oVar1S412(0) <='1';
          else
          oVar1S412(0) <='0';
          end if;
        if(cVar2S24S57N041P049nsss(0)='1'  )then
          oVar1S413(0) <='1';
          else
          oVar1S413(0) <='0';
          end if;
        if(cVar1S0S58P045P005P068nsss(0)='1'  OR cVar2S1S58P008nsss(0)='1'  OR cVar2S2S58P004P018nsss(0)='1'  OR cVar2S3S58N004P007P068nsss(0)='1'  )then
          oVar1S414(0) <='1';
          else
          oVar1S414(0) <='0';
          end if;
        if(cVar2S4S58N004N007P048nsss(0)='1'  OR cVar1S5S58N045P018P040P002nsss(0)='1'  OR cVar2S6S58P038P015nsss(0)='1'  OR cVar2S7S58N038P062nsss(0)='1'  )then
          oVar1S415(0) <='1';
          else
          oVar1S415(0) <='0';
          end if;
        if(cVar2S8S58N038N062P023nsss(0)='1'  OR cVar2S9S58P021P038P012nsss(0)='1'  OR cVar2S10S58P021P038P037nsss(0)='1'  OR cVar2S11S58P021P003nsss(0)='1'  )then
          oVar1S416(0) <='1';
          else
          oVar1S416(0) <='0';
          end if;
        if(cVar2S12S58P021N003P006nsss(0)='1'  OR cVar2S13S58P041P005nsss(0)='1'  OR cVar2S14S58P041N005P020nsss(0)='1'  OR cVar2S15S58N041P011nsss(0)='1'  )then
          oVar1S417(0) <='1';
          else
          oVar1S417(0) <='0';
          end if;
        if(cVar2S16S58N041N011P016nsss(0)='1'  OR cVar2S17S58P035P065nsss(0)='1'  OR cVar2S18S58P035N065P068nsss(0)='1'  OR cVar2S19S58N035P039nsss(0)='1'  )then
          oVar1S418(0) <='1';
          else
          oVar1S418(0) <='0';
          end if;
        if(cVar2S20S58N035N039P021nsss(0)='1'  OR cVar2S21S58P064nsss(0)='1'  OR cVar2S22S58N064P055nsss(0)='1'  OR cVar2S23S58P028P009nsss(0)='1'  )then
          oVar1S419(0) <='1';
          else
          oVar1S419(0) <='0';
          end if;
        if(cVar2S24S58N028P055P013nsss(0)='1'  OR cVar2S25S58P036P012nsss(0)='1'  OR cVar2S26S58P036N012P049nsss(0)='1'  )then
          oVar1S420(0) <='1';
          else
          oVar1S420(0) <='0';
          end if;
        if(cVar1S0S59P045P022P019nsss(0)='1'  OR cVar1S1S59P045P022N019P013nsss(0)='1'  OR cVar1S2S59P045N022P023nsss(0)='1'  OR cVar2S3S59P024nsss(0)='1'  )then
          oVar1S421(0) <='1';
          else
          oVar1S421(0) <='0';
          end if;
        if(cVar2S4S59P044nsss(0)='1'  OR cVar2S5S59N044P067nsss(0)='1'  OR cVar2S6S59N044N067P004nsss(0)='1'  OR cVar1S7S59N045P040P021P002nsss(0)='1'  )then
          oVar1S422(0) <='1';
          else
          oVar1S422(0) <='0';
          end if;
        if(cVar2S8S59P003nsss(0)='1'  OR cVar2S9S59N003P004nsss(0)='1'  OR cVar2S10S59N003N004P005nsss(0)='1'  OR cVar1S11S59N045P040N021P066nsss(0)='1'  )then
          oVar1S423(0) <='1';
          else
          oVar1S423(0) <='0';
          end if;
        if(cVar2S12S59P018P037nsss(0)='1'  OR cVar2S13S59P066nsss(0)='1'  OR cVar2S14S59P046P004nsss(0)='1'  OR cVar2S15S59P046N004P006nsss(0)='1'  )then
          oVar1S424(0) <='1';
          else
          oVar1S424(0) <='0';
          end if;
        if(cVar2S16S59N046P003P058nsss(0)='1'  OR cVar2S17S59P022P057P032nsss(0)='1'  OR cVar2S18S59P022P057P068nsss(0)='1'  OR cVar2S19S59P030P031P012nsss(0)='1'  )then
          oVar1S425(0) <='1';
          else
          oVar1S425(0) <='0';
          end if;
        if(cVar2S20S59N030P057P063nsss(0)='1'  OR cVar2S21S59N030P057P031nsss(0)='1'  )then
          oVar1S426(0) <='1';
          else
          oVar1S426(0) <='0';
          end if;
        if(cVar1S0S60P045P005P037nsss(0)='1'  OR cVar2S1S60P006nsss(0)='1'  OR cVar2S2S60N006P004nsss(0)='1'  OR cVar2S3S60N006N004P007nsss(0)='1'  )then
          oVar1S427(0) <='1';
          else
          oVar1S427(0) <='0';
          end if;
        if(cVar1S4S60P045N005P021N024psss(0)='1'  OR cVar2S5S60P021nsss(0)='1'  OR cVar2S6S60N021P039nsss(0)='1'  OR cVar2S7S60N021N039P038nsss(0)='1'  )then
          oVar1S428(0) <='1';
          else
          oVar1S428(0) <='0';
          end if;
        if(cVar2S8S60P049nsss(0)='1'  OR cVar2S9S60N049P021nsss(0)='1'  OR cVar2S10S60N049N021P062nsss(0)='1'  OR cVar2S11S60P065P030P031nsss(0)='1'  )then
          oVar1S429(0) <='1';
          else
          oVar1S429(0) <='0';
          end if;
        if(cVar2S12S60P065N030psss(0)='1'  OR cVar2S13S60P065P066P058nsss(0)='1'  OR cVar2S14S60P065P066P069nsss(0)='1'  OR cVar2S15S60P041P022nsss(0)='1'  )then
          oVar1S430(0) <='1';
          else
          oVar1S430(0) <='0';
          end if;
        if(cVar2S16S60P041N022P020nsss(0)='1'  OR cVar2S17S60N041P049nsss(0)='1'  OR cVar1S18S60N045P018P025P035nsss(0)='1'  OR cVar2S19S60P066P046nsss(0)='1'  )then
          oVar1S431(0) <='1';
          else
          oVar1S431(0) <='0';
          end if;
        if(cVar2S20S60P066N046P014nsss(0)='1'  OR cVar2S21S60P066P036nsss(0)='1'  OR cVar2S22S60N066P040nsss(0)='1'  OR cVar2S23S60P066P006P016nsss(0)='1'  )then
          oVar1S432(0) <='1';
          else
          oVar1S432(0) <='0';
          end if;
        if(cVar2S24S60P066N006P058nsss(0)='1'  OR cVar2S25S60P066P053nsss(0)='1'  )then
          oVar1S433(0) <='1';
          else
          oVar1S433(0) <='0';
          end if;
        if(cVar1S0S61P045P005P068P012nsss(0)='1'  OR cVar2S1S61P013nsss(0)='1'  OR cVar2S2S61N013P068nsss(0)='1'  OR cVar2S3S61P022nsss(0)='1'  )then
          oVar1S434(0) <='1';
          else
          oVar1S434(0) <='0';
          end if;
        if(cVar2S4S61N022P044nsss(0)='1'  OR cVar2S5S61N022N044P025nsss(0)='1'  OR cVar2S6S61P017P036nsss(0)='1'  OR cVar2S7S61N017P009nsss(0)='1'  )then
          oVar1S435(0) <='1';
          else
          oVar1S435(0) <='0';
          end if;
        if(cVar2S8S61N017N009P036nsss(0)='1'  OR cVar2S9S61P059P068P014nsss(0)='1'  OR cVar2S10S61P059N068psss(0)='1'  OR cVar2S11S61P059P055nsss(0)='1'  )then
          oVar1S436(0) <='1';
          else
          oVar1S436(0) <='0';
          end if;
        if(cVar2S12S61P006P016nsss(0)='1'  OR cVar2S13S61N006P068P054nsss(0)='1'  OR cVar2S14S61P016P003nsss(0)='1'  OR cVar2S15S61N016P024P031nsss(0)='1'  )then
          oVar1S437(0) <='1';
          else
          oVar1S437(0) <='0';
          end if;
        if(cVar1S16S61N045N018P040P002nsss(0)='1'  OR cVar2S17S61P049nsss(0)='1'  OR cVar2S18S61N049P034nsss(0)='1'  OR cVar2S19S61P028P010nsss(0)='1'  )then
          oVar1S438(0) <='1';
          else
          oVar1S438(0) <='0';
          end if;
        if(cVar2S20S61P028N010P011nsss(0)='1'  OR cVar2S21S61N028P029P011nsss(0)='1'  OR cVar2S22S61P063P060P036nsss(0)='1'  )then
          oVar1S439(0) <='1';
          else
          oVar1S439(0) <='0';
          end if;
        if(cVar1S0S62P045P005P068nsss(0)='1'  OR cVar2S1S62P006nsss(0)='1'  OR cVar2S2S62N006P004nsss(0)='1'  OR cVar2S3S62N006N004P047nsss(0)='1'  )then
          oVar1S440(0) <='1';
          else
          oVar1S440(0) <='0';
          end if;
        if(cVar2S4S62P014P022nsss(0)='1'  OR cVar2S5S62P014N022P013nsss(0)='1'  OR cVar2S6S62N014P061nsss(0)='1'  OR cVar2S7S62N014N061P003nsss(0)='1'  )then
          oVar1S441(0) <='1';
          else
          oVar1S441(0) <='0';
          end if;
        if(cVar2S8S62P031P012nsss(0)='1'  OR cVar2S9S62P031N012P010nsss(0)='1'  OR cVar2S10S62P031P013nsss(0)='1'  OR cVar2S11S62P031N013P011nsss(0)='1'  )then
          oVar1S442(0) <='1';
          else
          oVar1S442(0) <='0';
          end if;
        if(cVar2S12S62N031P054P011nsss(0)='1'  OR cVar2S13S62N031P054P029nsss(0)='1'  OR cVar1S14S62N045P018P000P040nsss(0)='1'  OR cVar2S15S62P035P013P019nsss(0)='1'  )then
          oVar1S443(0) <='1';
          else
          oVar1S443(0) <='0';
          end if;
        if(cVar2S16S62P035N013P003nsss(0)='1'  OR cVar1S17S62N045P018P061P035nsss(0)='1'  OR cVar2S18S62P014P034nsss(0)='1'  OR cVar2S19S62P014N034P037nsss(0)='1'  )then
          oVar1S444(0) <='1';
          else
          oVar1S444(0) <='0';
          end if;
        if(cVar2S20S62N014P015nsss(0)='1'  OR cVar2S21S62P035nsss(0)='1'  OR cVar2S22S62N035P011nsss(0)='1'  OR cVar2S23S62P063P065P067nsss(0)='1'  )then
          oVar1S445(0) <='1';
          else
          oVar1S445(0) <='0';
          end if;
        if(cVar2S24S62P063N065P006nsss(0)='1'  )then
          oVar1S446(0) <='1';
          else
          oVar1S446(0) <='0';
          end if;
        if(cVar1S0S63P045P005P037nsss(0)='1'  OR cVar2S1S63P068nsss(0)='1'  OR cVar2S2S63P006P004nsss(0)='1'  OR cVar2S3S63N006P004P018nsss(0)='1'  )then
          oVar1S447(0) <='1';
          else
          oVar1S447(0) <='0';
          end if;
        if(cVar2S4S63N006N004psss(0)='1'  OR cVar2S5S63P033P027P066nsss(0)='1'  OR cVar2S6S63P033N027psss(0)='1'  OR cVar2S7S63P033P059nsss(0)='1'  )then
          oVar1S448(0) <='1';
          else
          oVar1S448(0) <='0';
          end if;
        if(cVar2S8S63P033N059P036nsss(0)='1'  OR cVar2S9S63P064nsss(0)='1'  OR cVar2S10S63N064P013P031nsss(0)='1'  OR cVar2S11S63N064N013P030nsss(0)='1'  )then
          oVar1S449(0) <='1';
          else
          oVar1S449(0) <='0';
          end if;
        if(cVar2S12S63P007P031P013nsss(0)='1'  OR cVar2S13S63P007N031P004nsss(0)='1'  OR cVar2S14S63P007P049nsss(0)='1'  OR cVar2S15S63P007N049P025nsss(0)='1'  )then
          oVar1S450(0) <='1';
          else
          oVar1S450(0) <='0';
          end if;
        if(cVar2S16S63P036P014nsss(0)='1'  OR cVar2S17S63P035P063nsss(0)='1'  OR cVar2S18S63P035P011P019nsss(0)='1'  OR cVar2S19S63P013nsss(0)='1'  )then
          oVar1S451(0) <='1';
          else
          oVar1S451(0) <='0';
          end if;
        if(cVar2S20S63N013P011P016nsss(0)='1'  OR cVar2S21S63N013N011P012nsss(0)='1'  OR cVar2S22S63P057P014P060nsss(0)='1'  OR cVar2S23S63P057N014P069nsss(0)='1'  )then
          oVar1S452(0) <='1';
          else
          oVar1S452(0) <='0';
          end if;
        if(cVar2S24S63P057P028P010nsss(0)='1'  OR cVar2S25S63P057N028P060nsss(0)='1'  )then
          oVar1S453(0) <='1';
          else
          oVar1S453(0) <='0';
          end if;
        if(cVar2S0S64P053nsss(0)='1'  OR cVar2S1S64N053P054P057nsss(0)='1'  OR cVar2S2S64N053N054P052nsss(0)='1'  OR cVar2S3S64P020nsss(0)='1'  )then
          oVar1S454(0) <='1';
          else
          oVar1S454(0) <='0';
          end if;
        if(cVar2S4S64N020P014P056nsss(0)='1'  OR cVar2S5S64N020N014P063nsss(0)='1'  OR cVar2S6S64P045P004P006nsss(0)='1'  OR cVar2S7S64P045N004psss(0)='1'  )then
          oVar1S455(0) <='1';
          else
          oVar1S455(0) <='0';
          end if;
        if(cVar2S8S64N045P041P020nsss(0)='1'  OR cVar2S9S64N045N041P043nsss(0)='1'  OR cVar2S10S64P009nsss(0)='1'  OR cVar2S11S64N009P010P019nsss(0)='1'  )then
          oVar1S456(0) <='1';
          else
          oVar1S456(0) <='0';
          end if;
        if(cVar2S12S64P065nsss(0)='1'  OR cVar2S13S64N065P017P013nsss(0)='1'  OR cVar2S14S64N065P017P036nsss(0)='1'  OR cVar2S15S64P066P037nsss(0)='1'  )then
          oVar1S457(0) <='1';
          else
          oVar1S457(0) <='0';
          end if;
        if(cVar2S16S64P059nsss(0)='1'  OR cVar2S17S64N059P065nsss(0)='1'  OR cVar2S18S64P035P067P052nsss(0)='1'  OR cVar2S19S64P035P017P064nsss(0)='1'  )then
          oVar1S458(0) <='1';
          else
          oVar1S458(0) <='0';
          end if;
        if(cVar2S20S64P054nsss(0)='1'  OR cVar2S21S64N054P057nsss(0)='1'  OR cVar2S22S64N054N057P058nsss(0)='1'  OR cVar2S23S64P057P037nsss(0)='1'  )then
          oVar1S459(0) <='1';
          else
          oVar1S459(0) <='0';
          end if;
        if(cVar2S24S64P057N037P012nsss(0)='1'  OR cVar1S25S64P018N031P007P051nsss(0)='1'  OR cVar2S26S64P013P043nsss(0)='1'  OR cVar2S27S64P013N043P034nsss(0)='1'  )then
          oVar1S460(0) <='1';
          else
          oVar1S460(0) <='0';
          end if;
        if(cVar2S28S64P013P068nsss(0)='1'  OR cVar2S29S64P068P062nsss(0)='1'  OR cVar2S30S64P068P062P035nsss(0)='1'  OR cVar2S31S64P066P036P067nsss(0)='1'  )then
          oVar1S461(0) <='1';
          else
          oVar1S461(0) <='0';
          end if;
        if(cVar2S32S64P066N036P028nsss(0)='1'  OR cVar2S33S64N066P036P014nsss(0)='1'  OR cVar2S34S64N066P036P059nsss(0)='1'  )then
          oVar1S462(0) <='1';
          else
          oVar1S462(0) <='0';
          end if;
        if(cVar2S0S65P037P029P012nsss(0)='1'  OR cVar2S1S65P037P024P056nsss(0)='1'  OR cVar2S2S65P012P065nsss(0)='1'  OR cVar2S3S65N012P056P060nsss(0)='1'  )then
          oVar1S463(0) <='1';
          else
          oVar1S463(0) <='0';
          end if;
        if(cVar1S4S65P018P014P042P004nsss(0)='1'  OR cVar2S5S65P005nsss(0)='1'  OR cVar2S6S65N005P069nsss(0)='1'  OR cVar1S7S65P018P014P045nsss(0)='1'  )then
          oVar1S464(0) <='1';
          else
          oVar1S464(0) <='0';
          end if;
        if(cVar1S8S65P018P014N045P046nsss(0)='1'  OR cVar2S9S65P031P036nsss(0)='1'  OR cVar2S10S65P031N036P019nsss(0)='1'  OR cVar2S11S65N031P032nsss(0)='1'  )then
          oVar1S465(0) <='1';
          else
          oVar1S465(0) <='0';
          end if;
        if(cVar2S12S65N031N032P020nsss(0)='1'  OR cVar1S13S65N018P041P020P002nsss(0)='1'  OR cVar2S14S65P003nsss(0)='1'  OR cVar2S15S65N003P005nsss(0)='1'  )then
          oVar1S466(0) <='1';
          else
          oVar1S466(0) <='0';
          end if;
        if(cVar2S16S65P042nsss(0)='1'  OR cVar2S17S65P009P021nsss(0)='1'  OR cVar2S18S65P009N021P016nsss(0)='1'  OR cVar2S19S65P004P016nsss(0)='1'  )then
          oVar1S467(0) <='1';
          else
          oVar1S467(0) <='0';
          end if;
        if(cVar2S20S65N004psss(0)='1'  OR cVar2S21S65P011P029P010nsss(0)='1'  OR cVar2S22S65P011N029P014nsss(0)='1'  OR cVar2S23S65N011P020P040nsss(0)='1'  )then
          oVar1S468(0) <='1';
          else
          oVar1S468(0) <='0';
          end if;
        if(cVar1S24S65N018N041P039P049nsss(0)='1'  OR cVar2S25S65P005nsss(0)='1'  )then
          oVar1S469(0) <='1';
          else
          oVar1S469(0) <='0';
          end if;
        if(cVar1S0S66P018P041P020P002nsss(0)='1'  OR cVar2S1S66P003nsss(0)='1'  OR cVar2S2S66N003P005nsss(0)='1'  OR cVar2S3S66P042nsss(0)='1'  )then
          oVar1S470(0) <='1';
          else
          oVar1S470(0) <='0';
          end if;
        if(cVar2S4S66P009P021nsss(0)='1'  OR cVar2S5S66P009N021P047nsss(0)='1'  OR cVar2S6S66P009P027P066nsss(0)='1'  OR cVar2S7S66P009N027P049nsss(0)='1'  )then
          oVar1S471(0) <='1';
          else
          oVar1S471(0) <='0';
          end if;
        if(cVar2S8S66N009P027P007nsss(0)='1'  OR cVar2S9S66N009P027P007nsss(0)='1'  OR cVar2S10S66P011nsss(0)='1'  OR cVar2S11S66N011P007nsss(0)='1'  )then
          oVar1S472(0) <='1';
          else
          oVar1S472(0) <='0';
          end if;
        if(cVar2S12S66N011N007P040nsss(0)='1'  OR cVar2S13S66P005nsss(0)='1'  OR cVar1S14S66P018P068P057nsss(0)='1'  OR cVar2S15S66P041P036P035nsss(0)='1'  )then
          oVar1S473(0) <='1';
          else
          oVar1S473(0) <='0';
          end if;
        if(cVar2S16S66P041N036P032nsss(0)='1'  OR cVar2S17S66P017P036nsss(0)='1'  OR cVar2S18S66P017P036P019nsss(0)='1'  OR cVar2S19S66N017P016nsss(0)='1'  )then
          oVar1S474(0) <='1';
          else
          oVar1S474(0) <='0';
          end if;
        if(cVar2S20S66P010nsss(0)='1'  OR cVar2S21S66P057P012nsss(0)='1'  OR cVar2S22S66P057N012P014nsss(0)='1'  OR cVar2S23S66P069P063P046nsss(0)='1'  )then
          oVar1S475(0) <='1';
          else
          oVar1S475(0) <='0';
          end if;
        if(cVar2S24S66P002P034nsss(0)='1'  OR cVar2S25S66P002N034P013nsss(0)='1'  OR cVar2S26S66N002P038P027nsss(0)='1'  )then
          oVar1S476(0) <='1';
          else
          oVar1S476(0) <='0';
          end if;
        if(cVar1S0S67P009P027P063P018nsss(0)='1'  OR cVar2S1S67P019nsss(0)='1'  OR cVar2S2S67N019P052P048nsss(0)='1'  OR cVar1S3S67P009N027P049P026nsss(0)='1'  )then
          oVar1S477(0) <='1';
          else
          oVar1S477(0) <='0';
          end if;
        if(cVar2S4S67P025nsss(0)='1'  OR cVar2S5S67N025P024nsss(0)='1'  OR cVar2S6S67P001nsss(0)='1'  OR cVar2S7S67N001P000nsss(0)='1'  )then
          oVar1S478(0) <='1';
          else
          oVar1S478(0) <='0';
          end if;
        if(cVar2S8S67P012P065nsss(0)='1'  OR cVar2S9S67P012N065P006nsss(0)='1'  OR cVar2S10S67N012P017P050nsss(0)='1'  OR cVar1S11S67N009P041P020P039nsss(0)='1'  )then
          oVar1S479(0) <='1';
          else
          oVar1S479(0) <='0';
          end if;
        if(cVar1S12S67N009P041N020P021nsss(0)='1'  OR cVar2S13S67P018P007nsss(0)='1'  OR cVar2S14S67P018N007P068nsss(0)='1'  OR cVar2S15S67P018P012P043nsss(0)='1'  )then
          oVar1S480(0) <='1';
          else
          oVar1S480(0) <='0';
          end if;
        if(cVar2S16S67P003P036P067nsss(0)='1'  OR cVar2S17S67P003P036P019nsss(0)='1'  OR cVar2S18S67P031P013P068nsss(0)='1'  OR cVar2S19S67P031N013P057nsss(0)='1'  )then
          oVar1S481(0) <='1';
          else
          oVar1S481(0) <='0';
          end if;
        if(cVar2S20S67N031P004P038nsss(0)='1'  OR cVar2S21S67N031P004P017nsss(0)='1'  OR cVar2S22S67P020P015P008nsss(0)='1'  OR cVar2S23S67P020N015P016nsss(0)='1'  )then
          oVar1S482(0) <='1';
          else
          oVar1S482(0) <='0';
          end if;
        if(cVar2S24S67P020P019P015nsss(0)='1'  OR cVar2S25S67P020N019P011nsss(0)='1'  OR cVar2S26S67P011P005nsss(0)='1'  )then
          oVar1S483(0) <='1';
          else
          oVar1S483(0) <='0';
          end if;
        if(cVar1S0S68P009P027P063P018nsss(0)='1'  OR cVar2S1S68P019nsss(0)='1'  OR cVar1S2S68P009N027P049P026nsss(0)='1'  OR cVar2S3S68P025nsss(0)='1'  )then
          oVar1S484(0) <='1';
          else
          oVar1S484(0) <='0';
          end if;
        if(cVar2S4S68N025P019P024nsss(0)='1'  OR cVar2S5S68P029nsss(0)='1'  OR cVar2S6S68N029P051P015nsss(0)='1'  OR cVar2S7S68P015P064P033nsss(0)='1'  )then
          oVar1S485(0) <='1';
          else
          oVar1S485(0) <='0';
          end if;
        if(cVar2S8S68P015P064P063nsss(0)='1'  OR cVar2S9S68N015P034nsss(0)='1'  OR cVar2S10S68N015N034P023nsss(0)='1'  OR cVar1S11S68N009P041P020P003nsss(0)='1'  )then
          oVar1S486(0) <='1';
          else
          oVar1S486(0) <='0';
          end if;
        if(cVar2S12S68P002nsss(0)='1'  OR cVar2S13S68N002P004nsss(0)='1'  OR cVar2S14S68N002N004P005nsss(0)='1'  OR cVar2S15S68P038nsss(0)='1'  )then
          oVar1S487(0) <='1';
          else
          oVar1S487(0) <='0';
          end if;
        if(cVar2S16S68N038P042nsss(0)='1'  OR cVar2S17S68P018P007nsss(0)='1'  OR cVar2S18S68P018N007P047nsss(0)='1'  OR cVar2S19S68P018P012P043nsss(0)='1'  )then
          oVar1S488(0) <='1';
          else
          oVar1S488(0) <='0';
          end if;
        if(cVar2S20S68P054P013nsss(0)='1'  OR cVar2S21S68P054N013P019nsss(0)='1'  OR cVar2S22S68N054P013nsss(0)='1'  OR cVar2S23S68N054N013P011nsss(0)='1'  )then
          oVar1S489(0) <='1';
          else
          oVar1S489(0) <='0';
          end if;
        if(cVar2S24S68P020P039nsss(0)='1'  OR cVar2S25S68P020P039P045nsss(0)='1'  OR cVar2S26S68P020P050P003nsss(0)='1'  OR cVar2S27S68P035P053P030nsss(0)='1'  )then
          oVar1S490(0) <='1';
          else
          oVar1S490(0) <='0';
          end if;
        if(cVar2S28S68P035P029P037nsss(0)='1'  OR cVar2S29S68P018P014nsss(0)='1'  OR cVar2S30S68P018P014P017nsss(0)='1'  OR cVar2S31S68N018P069P019nsss(0)='1'  )then
          oVar1S491(0) <='1';
          else
          oVar1S491(0) <='0';
          end if;
        if(cVar2S0S69P013P051nsss(0)='1'  OR cVar2S1S69P013P051P047nsss(0)='1'  OR cVar2S2S69P013psss(0)='1'  OR cVar1S3S69P009N049P053P029nsss(0)='1'  )then
          oVar1S493(0) <='1';
          else
          oVar1S493(0) <='0';
          end if;
        if(cVar2S4S69P051P007nsss(0)='1'  OR cVar2S5S69N051P019nsss(0)='1'  OR cVar2S6S69P027P013nsss(0)='1'  OR cVar2S7S69N027P029P011nsss(0)='1'  )then
          oVar1S494(0) <='1';
          else
          oVar1S494(0) <='0';
          end if;
        if(cVar2S8S69N027N029P015nsss(0)='1'  OR cVar2S9S69P051P019P002nsss(0)='1'  OR cVar2S10S69P051N019P066nsss(0)='1'  OR cVar1S11S69N009P041P020P003nsss(0)='1'  )then
          oVar1S495(0) <='1';
          else
          oVar1S495(0) <='0';
          end if;
        if(cVar2S12S69P002nsss(0)='1'  OR cVar2S13S69N002P004nsss(0)='1'  OR cVar2S14S69N002N004P005nsss(0)='1'  OR cVar1S15S69N009P041N020P001nsss(0)='1'  )then
          oVar1S496(0) <='1';
          else
          oVar1S496(0) <='0';
          end if;
        if(cVar2S16S69P021P040nsss(0)='1'  OR cVar2S17S69P021P040P042nsss(0)='1'  OR cVar2S18S69N021P039P043nsss(0)='1'  OR cVar2S19S69P054P012P065nsss(0)='1'  )then
          oVar1S497(0) <='1';
          else
          oVar1S497(0) <='0';
          end if;
        if(cVar2S20S69P054P012psss(0)='1'  OR cVar2S21S69N054P057nsss(0)='1'  OR cVar2S22S69N054N057P058nsss(0)='1'  OR cVar2S23S69P054P016nsss(0)='1'  )then
          oVar1S498(0) <='1';
          else
          oVar1S498(0) <='0';
          end if;
        if(cVar2S24S69N054P018P012nsss(0)='1'  OR cVar2S25S69P039P016P059nsss(0)='1'  OR cVar2S26S69P039N016P025nsss(0)='1'  OR cVar2S27S69P039P011P064nsss(0)='1'  )then
          oVar1S499(0) <='1';
          else
          oVar1S499(0) <='0';
          end if;
        if(cVar2S28S69P011P029nsss(0)='1'  OR cVar2S29S69P011N029P012nsss(0)='1'  OR cVar2S30S69N011P010nsss(0)='1'  OR cVar2S31S69N011N010P030nsss(0)='1'  )then
          oVar1S500(0) <='1';
          else
          oVar1S500(0) <='0';
          end if;
        if(cVar2S0S70P014P028P015nsss(0)='1'  OR cVar2S1S70P014N028psss(0)='1'  OR cVar2S2S70P014P009nsss(0)='1'  OR cVar2S3S70P023P005nsss(0)='1'  )then
          oVar1S502(0) <='1';
          else
          oVar1S502(0) <='0';
          end if;
        if(cVar2S4S70P023N005P017nsss(0)='1'  OR cVar2S5S70N023P049P026nsss(0)='1'  OR cVar2S6S70N023N049P047nsss(0)='1'  OR cVar2S7S70P037P056nsss(0)='1'  )then
          oVar1S503(0) <='1';
          else
          oVar1S503(0) <='0';
          end if;
        if(cVar2S8S70P037P019nsss(0)='1'  OR cVar2S9S70P019P065nsss(0)='1'  OR cVar2S10S70P019N065P015nsss(0)='1'  OR cVar2S11S70N019P065P011nsss(0)='1'  )then
          oVar1S504(0) <='1';
          else
          oVar1S504(0) <='0';
          end if;
        if(cVar2S12S70P013nsss(0)='1'  OR cVar2S13S70P047P009nsss(0)='1'  OR cVar2S14S70P047P009nsss(0)='1'  OR cVar2S15S70P047N009P017nsss(0)='1'  )then
          oVar1S505(0) <='1';
          else
          oVar1S505(0) <='0';
          end if;
        if(cVar2S16S70P049nsss(0)='1'  OR cVar2S17S70N049P052nsss(0)='1'  OR cVar2S18S70P040nsss(0)='1'  OR cVar2S19S70N040P012nsss(0)='1'  )then
          oVar1S506(0) <='1';
          else
          oVar1S506(0) <='0';
          end if;
        if(cVar2S20S70P042P047P068nsss(0)='1'  OR cVar2S21S70P042P005nsss(0)='1'  OR cVar2S22S70P042N005P012nsss(0)='1'  OR cVar2S23S70P019nsss(0)='1'  )then
          oVar1S507(0) <='1';
          else
          oVar1S507(0) <='0';
          end if;
        if(cVar2S24S70P036P015P019nsss(0)='1'  OR cVar2S25S70P036N015P009nsss(0)='1'  OR cVar1S26S70P016P035P032P018nsss(0)='1'  OR cVar2S27S70P010P009P015nsss(0)='1'  )then
          oVar1S508(0) <='1';
          else
          oVar1S508(0) <='0';
          end if;
        if(cVar1S0S71P041P020P003nsss(0)='1'  OR cVar1S1S71P041P020N003P002nsss(0)='1'  OR cVar2S2S71P004nsss(0)='1'  OR cVar2S3S71N004P005nsss(0)='1'  )then
          oVar1S510(0) <='1';
          else
          oVar1S510(0) <='0';
          end if;
        if(cVar1S4S71P041N020P001nsss(0)='1'  OR cVar2S5S71P021P040nsss(0)='1'  OR cVar2S6S71N021P022nsss(0)='1'  OR cVar2S7S71N021N022P042nsss(0)='1'  )then
          oVar1S511(0) <='1';
          else
          oVar1S511(0) <='0';
          end if;
        if(cVar2S8S71P039P067nsss(0)='1'  OR cVar2S9S71P039N067P022nsss(0)='1'  OR cVar2S10S71P039P017P021nsss(0)='1'  OR cVar2S11S71P024nsss(0)='1'  )then
          oVar1S512(0) <='1';
          else
          oVar1S512(0) <='0';
          end if;
        if(cVar2S12S71P006nsss(0)='1'  OR cVar2S13S71N006P016nsss(0)='1'  OR cVar2S14S71P027P048nsss(0)='1'  OR cVar2S15S71P027P048P047nsss(0)='1'  )then
          oVar1S513(0) <='1';
          else
          oVar1S513(0) <='0';
          end if;
        if(cVar2S16S71N027P025nsss(0)='1'  OR cVar2S17S71P007P037nsss(0)='1'  OR cVar2S18S71N007P004P013nsss(0)='1'  OR cVar2S19S71N007N004P005nsss(0)='1'  )then
          oVar1S514(0) <='1';
          else
          oVar1S514(0) <='0';
          end if;
        if(cVar2S20S71P047P016P035nsss(0)='1'  OR cVar2S21S71P047N016P053nsss(0)='1'  OR cVar2S22S71P047P069nsss(0)='1'  OR cVar2S23S71P047N069P008nsss(0)='1'  )then
          oVar1S515(0) <='1';
          else
          oVar1S515(0) <='0';
          end if;
        if(cVar1S24S71N041N049P039P036nsss(0)='1'  OR cVar2S25S71P011P020nsss(0)='1'  OR cVar2S26S71P011N020P013nsss(0)='1'  )then
          oVar1S516(0) <='1';
          else
          oVar1S516(0) <='0';
          end if;
        if(cVar1S0S72P016P018P023P042nsss(0)='1'  OR cVar2S1S72P043nsss(0)='1'  OR cVar2S2S72N043P017P019nsss(0)='1'  OR cVar2S3S72P006nsss(0)='1'  )then
          oVar1S517(0) <='1';
          else
          oVar1S517(0) <='0';
          end if;
        if(cVar2S4S72N006P008nsss(0)='1'  OR cVar2S5S72N006N008P007nsss(0)='1'  OR cVar2S6S72P028P032nsss(0)='1'  OR cVar2S7S72N028P031P054nsss(0)='1'  )then
          oVar1S518(0) <='1';
          else
          oVar1S518(0) <='0';
          end if;
        if(cVar2S8S72N028N031P054nsss(0)='1'  OR cVar1S9S72P016P018P045P015nsss(0)='1'  OR cVar2S10S72P017nsss(0)='1'  OR cVar2S11S72P047P028nsss(0)='1'  )then
          oVar1S519(0) <='1';
          else
          oVar1S519(0) <='0';
          end if;
        if(cVar2S12S72P047N028P054nsss(0)='1'  OR cVar2S13S72P047P009nsss(0)='1'  OR cVar2S14S72P047N009P017nsss(0)='1'  OR cVar2S15S72P031nsss(0)='1'  )then
          oVar1S520(0) <='1';
          else
          oVar1S520(0) <='0';
          end if;
        if(cVar2S16S72N031P046nsss(0)='1'  OR cVar2S17S72N031N046P029nsss(0)='1'  OR cVar2S18S72P019P020nsss(0)='1'  OR cVar2S19S72P019P039nsss(0)='1'  )then
          oVar1S521(0) <='1';
          else
          oVar1S521(0) <='0';
          end if;
        if(cVar2S20S72P029nsss(0)='1'  OR cVar2S21S72N029P007nsss(0)='1'  OR cVar2S22S72N029P007P014nsss(0)='1'  OR cVar2S23S72P053P004nsss(0)='1'  )then
          oVar1S522(0) <='1';
          else
          oVar1S522(0) <='0';
          end if;
        if(cVar2S24S72P053P011P019nsss(0)='1'  OR cVar2S25S72P013nsss(0)='1'  OR cVar2S26S72N013P015nsss(0)='1'  OR cVar2S27S72P007nsss(0)='1'  )then
          oVar1S523(0) <='1';
          else
          oVar1S523(0) <='0';
          end if;
        if(cVar2S28S72N007P018P003nsss(0)='1'  OR cVar2S29S72N007N018P037nsss(0)='1'  OR cVar2S30S72P036nsss(0)='1'  )then
          oVar1S524(0) <='1';
          else
          oVar1S524(0) <='0';
          end if;
        if(cVar1S0S73P047P006P024nsss(0)='1'  OR cVar1S1S73P047P006N024P026nsss(0)='1'  OR cVar1S2S73P047N006P008P026nsss(0)='1'  OR cVar2S3S73P049nsss(0)='1'  )then
          oVar1S525(0) <='1';
          else
          oVar1S525(0) <='0';
          end if;
        if(cVar2S4S73P015P068nsss(0)='1'  OR cVar2S5S73P009P017nsss(0)='1'  OR cVar2S6S73N009P005nsss(0)='1'  OR cVar2S7S73N009N005P069nsss(0)='1'  )then
          oVar1S526(0) <='1';
          else
          oVar1S526(0) <='0';
          end if;
        if(cVar2S8S73P012nsss(0)='1'  OR cVar2S9S73P012P017nsss(0)='1'  OR cVar2S10S73P057nsss(0)='1'  OR cVar2S11S73N057P060P015nsss(0)='1'  )then
          oVar1S527(0) <='1';
          else
          oVar1S527(0) <='0';
          end if;
        if(cVar2S12S73N057N060P016nsss(0)='1'  OR cVar2S13S73P008P055nsss(0)='1'  OR cVar2S14S73P008N055P016nsss(0)='1'  OR cVar2S15S73P055P012nsss(0)='1'  )then
          oVar1S528(0) <='1';
          else
          oVar1S528(0) <='0';
          end if;
        if(cVar2S16S73P055N012P018nsss(0)='1'  OR cVar2S17S73P056nsss(0)='1'  OR cVar2S18S73N056P057P065nsss(0)='1'  OR cVar2S19S73N056N057P059nsss(0)='1'  )then
          oVar1S529(0) <='1';
          else
          oVar1S529(0) <='0';
          end if;
        if(cVar2S20S73P010P057nsss(0)='1'  OR cVar2S21S73P010N057P017nsss(0)='1'  OR cVar2S22S73N010P013P057nsss(0)='1'  OR cVar2S23S73P019P066P065nsss(0)='1'  )then
          oVar1S530(0) <='1';
          else
          oVar1S530(0) <='0';
          end if;
        if(cVar2S24S73P019N066P013nsss(0)='1'  OR cVar2S25S73N019P068P064nsss(0)='1'  OR cVar2S26S73P032nsss(0)='1'  OR cVar2S27S73N032P028P010nsss(0)='1'  )then
          oVar1S531(0) <='1';
          else
          oVar1S531(0) <='0';
          end if;
        if(cVar2S28S73N032N028P068nsss(0)='1'  )then
          oVar1S532(0) <='1';
          else
          oVar1S532(0) <='0';
          end if;
        if(cVar2S0S74P017P015nsss(0)='1'  OR cVar2S1S74P017P015P048nsss(0)='1'  OR cVar2S2S74P017P052nsss(0)='1'  OR cVar2S3S74P017N052P019nsss(0)='1'  )then
          oVar1S533(0) <='1';
          else
          oVar1S533(0) <='0';
          end if;
        if(cVar2S4S74P007nsss(0)='1'  OR cVar2S5S74N007P008nsss(0)='1'  OR cVar2S6S74N007N008P011nsss(0)='1'  OR cVar2S7S74P020P003nsss(0)='1'  )then
          oVar1S534(0) <='1';
          else
          oVar1S534(0) <='0';
          end if;
        if(cVar2S8S74P020N003P002nsss(0)='1'  OR cVar2S9S74N020P005nsss(0)='1'  OR cVar2S10S74N020N005P012nsss(0)='1'  OR cVar2S11S74P029P011P008nsss(0)='1'  )then
          oVar1S535(0) <='1';
          else
          oVar1S535(0) <='0';
          end if;
        if(cVar2S12S74P029N011P009nsss(0)='1'  OR cVar2S13S74N029P028nsss(0)='1'  OR cVar2S14S74N029N028P053nsss(0)='1'  OR cVar2S15S74P023P042P012nsss(0)='1'  )then
          oVar1S536(0) <='1';
          else
          oVar1S536(0) <='0';
          end if;
        if(cVar2S16S74P023P042nsss(0)='1'  OR cVar2S17S74P068P013nsss(0)='1'  OR cVar2S18S74P012P018nsss(0)='1'  OR cVar2S19S74N012P011nsss(0)='1'  )then
          oVar1S537(0) <='1';
          else
          oVar1S537(0) <='0';
          end if;
        if(cVar1S20S74P064P011P042P017nsss(0)='1'  OR cVar2S21S74P029P009P067nsss(0)='1'  OR cVar2S22S74P029P009P027nsss(0)='1'  OR cVar2S23S74P010nsss(0)='1'  )then
          oVar1S538(0) <='1';
          else
          oVar1S538(0) <='0';
          end if;
        if(cVar2S24S74N010P009nsss(0)='1'  OR cVar1S25S74P064P011P017P054nsss(0)='1'  OR cVar2S26S74P033P062P018nsss(0)='1'  OR cVar2S27S74P033N062P066nsss(0)='1'  )then
          oVar1S539(0) <='1';
          else
          oVar1S539(0) <='0';
          end if;
        if(cVar2S28S74P014nsss(0)='1'  OR cVar2S29S74P016P066nsss(0)='1'  )then
          oVar1S540(0) <='1';
          else
          oVar1S540(0) <='0';
          end if;
        if(cVar1S0S75P029P011P051nsss(0)='1'  OR cVar2S1S75P050P057nsss(0)='1'  OR cVar2S2S75P050P056nsss(0)='1'  OR cVar2S3S75P008P068nsss(0)='1'  )then
          oVar1S541(0) <='1';
          else
          oVar1S541(0) <='0';
          end if;
        if(cVar1S4S75P029N011P010P052nsss(0)='1'  OR cVar2S5S75P054nsss(0)='1'  OR cVar2S6S75P050nsss(0)='1'  OR cVar2S7S75N050P053nsss(0)='1'  )then
          oVar1S542(0) <='1';
          else
          oVar1S542(0) <='0';
          end if;
        if(cVar2S8S75N050N053P054nsss(0)='1'  OR cVar2S9S75P015P019nsss(0)='1'  OR cVar2S10S75N015P013nsss(0)='1'  OR cVar1S11S75N029P041P020P003nsss(0)='1'  )then
          oVar1S543(0) <='1';
          else
          oVar1S543(0) <='0';
          end if;
        if(cVar2S12S75P002nsss(0)='1'  OR cVar2S13S75N002P004nsss(0)='1'  OR cVar2S14S75N002N004P005nsss(0)='1'  OR cVar2S15S75P021P040nsss(0)='1'  )then
          oVar1S544(0) <='1';
          else
          oVar1S544(0) <='0';
          end if;
        if(cVar2S16S75N021P022nsss(0)='1'  OR cVar2S17S75N021N022P042nsss(0)='1'  OR cVar2S18S75P001nsss(0)='1'  OR cVar2S19S75N001P039P033nsss(0)='1'  )then
          oVar1S545(0) <='1';
          else
          oVar1S545(0) <='0';
          end if;
        if(cVar1S20S75N029N041P045P023nsss(0)='1'  OR cVar2S21S75P022nsss(0)='1'  OR cVar2S22S75N022P024nsss(0)='1'  OR cVar2S23S75N022N024P036nsss(0)='1'  )then
          oVar1S546(0) <='1';
          else
          oVar1S546(0) <='0';
          end if;
        if(cVar2S24S75P049nsss(0)='1'  OR cVar2S25S75N049P066P009nsss(0)='1'  OR cVar2S26S75P028P010P031nsss(0)='1'  OR cVar2S27S75N028P040P021nsss(0)='1'  )then
          oVar1S547(0) <='1';
          else
          oVar1S547(0) <='0';
          end if;
        if(cVar2S0S76P050P013nsss(0)='1'  OR cVar2S1S76N050P017nsss(0)='1'  OR cVar2S2S76P033nsss(0)='1'  OR cVar1S3S76P064P027P066P068nsss(0)='1'  )then
          oVar1S549(0) <='1';
          else
          oVar1S549(0) <='0';
          end if;
        if(cVar2S4S76P013nsss(0)='1'  OR cVar2S5S76N013P050nsss(0)='1'  OR cVar2S6S76P003nsss(0)='1'  OR cVar2S7S76N003P002nsss(0)='1'  )then
          oVar1S550(0) <='1';
          else
          oVar1S550(0) <='0';
          end if;
        if(cVar2S8S76N003N002P019nsss(0)='1'  OR cVar2S9S76P005P040nsss(0)='1'  OR cVar2S10S76N005P001nsss(0)='1'  OR cVar2S11S76N005N001P022nsss(0)='1'  )then
          oVar1S551(0) <='1';
          else
          oVar1S551(0) <='0';
          end if;
        if(cVar2S12S76P034P063P006nsss(0)='1'  OR cVar2S13S76P034N063P062nsss(0)='1'  OR cVar2S14S76N034P063P017nsss(0)='1'  OR cVar2S15S76N034P063P036nsss(0)='1'  )then
          oVar1S552(0) <='1';
          else
          oVar1S552(0) <='0';
          end if;
        if(cVar2S16S76P042nsss(0)='1'  OR cVar2S17S76N042P033nsss(0)='1'  OR cVar1S18S76P064P042nsss(0)='1'  OR cVar2S19S76P046nsss(0)='1'  )then
          oVar1S553(0) <='1';
          else
          oVar1S553(0) <='0';
          end if;
        if(cVar2S20S76N046P034P068nsss(0)='1'  OR cVar2S21S76N046P034P014nsss(0)='1'  OR cVar2S22S76P014nsss(0)='1'  OR cVar2S23S76P019P016nsss(0)='1'  )then
          oVar1S554(0) <='1';
          else
          oVar1S554(0) <='0';
          end if;
        if(cVar2S24S76N019P068nsss(0)='1'  )then
          oVar1S555(0) <='1';
          else
          oVar1S555(0) <='0';
          end if;
        if(cVar2S0S77P057P068P013nsss(0)='1'  OR cVar2S1S77P057P068P013nsss(0)='1'  OR cVar2S2S77P018nsss(0)='1'  OR cVar2S3S77P067nsss(0)='1'  )then
          oVar1S556(0) <='1';
          else
          oVar1S556(0) <='0';
          end if;
        if(cVar2S4S77N067P003nsss(0)='1'  OR cVar2S5S77N067N003P037nsss(0)='1'  OR cVar2S6S77P039P016P063nsss(0)='1'  OR cVar2S7S77P039N016P002nsss(0)='1'  )then
          oVar1S557(0) <='1';
          else
          oVar1S557(0) <='0';
          end if;
        if(cVar2S8S77P039P015nsss(0)='1'  OR cVar1S9S77P017P064P050P016nsss(0)='1'  OR cVar2S10S77P015P052P055nsss(0)='1'  OR cVar2S11S77P015P018P065nsss(0)='1'  )then
          oVar1S558(0) <='1';
          else
          oVar1S558(0) <='0';
          end if;
        if(cVar2S12S77P015N018P033nsss(0)='1'  OR cVar1S13S77N017P041P020P003nsss(0)='1'  OR cVar2S14S77P002nsss(0)='1'  OR cVar2S15S77N002P004nsss(0)='1'  )then
          oVar1S559(0) <='1';
          else
          oVar1S559(0) <='0';
          end if;
        if(cVar2S16S77P039nsss(0)='1'  OR cVar2S17S77N039P043nsss(0)='1'  OR cVar2S18S77N039N043P016nsss(0)='1'  OR cVar2S19S77P019nsss(0)='1'  )then
          oVar1S560(0) <='1';
          else
          oVar1S560(0) <='0';
          end if;
        if(cVar2S20S77P009nsss(0)='1'  OR cVar2S21S77N009P008nsss(0)='1'  OR cVar2S22S77N009N008P006nsss(0)='1'  OR cVar2S23S77P023P042P008nsss(0)='1'  )then
          oVar1S561(0) <='1';
          else
          oVar1S561(0) <='0';
          end if;
        if(cVar2S24S77P023N042P037nsss(0)='1'  OR cVar2S25S77N023P013P031nsss(0)='1'  OR cVar2S26S77N023N013P065nsss(0)='1'  OR cVar2S27S77P003P052nsss(0)='1'  )then
          oVar1S562(0) <='1';
          else
          oVar1S562(0) <='0';
          end if;
        if(cVar2S28S77P003N052P016nsss(0)='1'  OR cVar2S29S77P003N034P013nsss(0)='1'  OR cVar2S30S77P008P058nsss(0)='1'  )then
          oVar1S563(0) <='1';
          else
          oVar1S563(0) <='0';
          end if;
        if(cVar2S0S78P049nsss(0)='1'  OR cVar2S1S78N049P066nsss(0)='1'  OR cVar2S2S78P011P068nsss(0)='1'  OR cVar2S3S78P011P068P019nsss(0)='1'  )then
          oVar1S564(0) <='1';
          else
          oVar1S564(0) <='0';
          end if;
        if(cVar2S4S78P011P015P003nsss(0)='1'  OR cVar2S5S78P011N015P012nsss(0)='1'  OR cVar2S6S78P011P033nsss(0)='1'  OR cVar2S7S78N011P015P013nsss(0)='1'  )then
          oVar1S565(0) <='1';
          else
          oVar1S565(0) <='0';
          end if;
        if(cVar2S8S78N011N015P018nsss(0)='1'  OR cVar2S9S78P028P053P012nsss(0)='1'  OR cVar2S10S78P028N053P054nsss(0)='1'  OR cVar2S11S78N028P026nsss(0)='1'  )then
          oVar1S566(0) <='1';
          else
          oVar1S566(0) <='0';
          end if;
        if(cVar2S12S78N028N026P051nsss(0)='1'  OR cVar2S13S78P036P034nsss(0)='1'  OR cVar2S14S78P036P034P016nsss(0)='1'  OR cVar2S15S78P036P016nsss(0)='1'  )then
          oVar1S567(0) <='1';
          else
          oVar1S567(0) <='0';
          end if;
        if(cVar2S16S78P064P006P031nsss(0)='1'  OR cVar2S17S78P064P014nsss(0)='1'  OR cVar2S18S78P036P007P015nsss(0)='1'  OR cVar2S19S78N036P065P066nsss(0)='1'  )then
          oVar1S568(0) <='1';
          else
          oVar1S568(0) <='0';
          end if;
        if(cVar2S20S78N036P065P037nsss(0)='1'  OR cVar2S21S78P064P010nsss(0)='1'  OR cVar2S22S78P064P068nsss(0)='1'  OR cVar2S23S78P064N068P061nsss(0)='1'  )then
          oVar1S569(0) <='1';
          else
          oVar1S569(0) <='0';
          end if;
        if(cVar2S24S78P064P059P014nsss(0)='1'  OR cVar2S25S78P064P059P063nsss(0)='1'  OR cVar2S26S78N064P052nsss(0)='1'  OR cVar2S27S78N064N052P051nsss(0)='1'  )then
          oVar1S570(0) <='1';
          else
          oVar1S570(0) <='0';
          end if;
        if(cVar1S28S78P062P026P068nsss(0)='1'  )then
          oVar1S571(0) <='1';
          else
          oVar1S571(0) <='0';
          end if;
        if(cVar1S0S79P051P008P065P028nsss(0)='1'  OR cVar2S1S79P026P068nsss(0)='1'  OR cVar2S2S79N026P053nsss(0)='1'  OR cVar1S3S79P051N008P042nsss(0)='1'  )then
          oVar1S572(0) <='1';
          else
          oVar1S572(0) <='0';
          end if;
        if(cVar2S4S79P053P029nsss(0)='1'  OR cVar2S5S79P053N029P052nsss(0)='1'  OR cVar2S6S79N053P049nsss(0)='1'  OR cVar2S7S79P011P053P012nsss(0)='1'  )then
          oVar1S573(0) <='1';
          else
          oVar1S573(0) <='0';
          end if;
        if(cVar2S8S79N011P007nsss(0)='1'  OR cVar2S9S79N011N007P034nsss(0)='1'  OR cVar1S10S79N051P041P020P003nsss(0)='1'  OR cVar2S11S79P002nsss(0)='1'  )then
          oVar1S574(0) <='1';
          else
          oVar1S574(0) <='0';
          end if;
        if(cVar2S12S79N002P005nsss(0)='1'  OR cVar2S13S79N002N005P004nsss(0)='1'  OR cVar1S14S79N051P041N020P001nsss(0)='1'  OR cVar2S15S79P021P005P040nsss(0)='1'  )then
          oVar1S575(0) <='1';
          else
          oVar1S575(0) <='0';
          end if;
        if(cVar2S16S79P021N005psss(0)='1'  OR cVar2S17S79N021P039P067nsss(0)='1'  OR cVar2S18S79P009nsss(0)='1'  OR cVar2S19S79N009P024P012nsss(0)='1'  )then
          oVar1S576(0) <='1';
          else
          oVar1S576(0) <='0';
          end if;
        if(cVar2S20S79P024P006P008nsss(0)='1'  OR cVar2S21S79P024N006psss(0)='1'  OR cVar2S22S79N024P027nsss(0)='1'  OR cVar2S23S79N024N027P025nsss(0)='1'  )then
          oVar1S577(0) <='1';
          else
          oVar1S577(0) <='0';
          end if;
        if(cVar2S24S79P032P011P019nsss(0)='1'  OR cVar2S25S79P032P011P057nsss(0)='1'  OR cVar2S26S79N032P028P010nsss(0)='1'  OR cVar2S27S79P034nsss(0)='1'  )then
          oVar1S578(0) <='1';
          else
          oVar1S578(0) <='0';
          end if;
        if(cVar2S28S79N034P033nsss(0)='1'  OR cVar2S29S79N034N033P035nsss(0)='1'  )then
          oVar1S579(0) <='1';
          else
          oVar1S579(0) <='0';
          end if;
        if(cVar1S0S80P040P002P021nsss(0)='1'  OR cVar1S1S80P040P002N021P041nsss(0)='1'  OR cVar2S2S80P038nsss(0)='1'  OR cVar1S3S80P040N002P057nsss(0)='1'  )then
          oVar1S580(0) <='1';
          else
          oVar1S580(0) <='0';
          end if;
        if(cVar2S4S80P023nsss(0)='1'  OR cVar2S5S80N023P022nsss(0)='1'  OR cVar2S6S80N023N022P038nsss(0)='1'  OR cVar2S7S80P000nsss(0)='1'  )then
          oVar1S581(0) <='1';
          else
          oVar1S581(0) <='0';
          end if;
        if(cVar2S8S80N000P050nsss(0)='1'  OR cVar2S9S80N000N050P005nsss(0)='1'  OR cVar2S10S80P066nsss(0)='1'  OR cVar2S11S80P066P018nsss(0)='1'  )then
          oVar1S582(0) <='1';
          else
          oVar1S582(0) <='0';
          end if;
        if(cVar2S12S80P055nsss(0)='1'  OR cVar2S13S80P055P010nsss(0)='1'  OR cVar2S14S80P053P064P012nsss(0)='1'  OR cVar2S15S80N053P002P005nsss(0)='1'  )then
          oVar1S583(0) <='1';
          else
          oVar1S583(0) <='0';
          end if;
        if(cVar2S16S80P029P011P058nsss(0)='1'  OR cVar2S17S80P029N011P063nsss(0)='1'  OR cVar2S18S80N029P062P027nsss(0)='1'  OR cVar2S19S80N029N062psss(0)='1'  )then
          oVar1S584(0) <='1';
          else
          oVar1S584(0) <='0';
          end if;
        if(cVar1S20S80N040P021P042nsss(0)='1'  OR cVar2S21S80P019nsss(0)='1'  OR cVar2S22S80N019P039nsss(0)='1'  OR cVar2S23S80P008P015nsss(0)='1'  )then
          oVar1S585(0) <='1';
          else
          oVar1S585(0) <='0';
          end if;
        if(cVar2S24S80N008P015P066nsss(0)='1'  )then
          oVar1S586(0) <='1';
          else
          oVar1S586(0) <='0';
          end if;
        if(cVar1S0S81P040P002nsss(0)='1'  OR cVar1S1S81P040N002P057nsss(0)='1'  OR cVar2S2S81P023nsss(0)='1'  OR cVar2S3S81N023P022nsss(0)='1'  )then
          oVar1S587(0) <='1';
          else
          oVar1S587(0) <='0';
          end if;
        if(cVar2S4S81N023N022P038nsss(0)='1'  OR cVar2S5S81P020P015nsss(0)='1'  OR cVar2S6S81P014nsss(0)='1'  OR cVar2S7S81P014P010nsss(0)='1'  )then
          oVar1S588(0) <='1';
          else
          oVar1S588(0) <='0';
          end if;
        if(cVar2S8S81P068P031nsss(0)='1'  OR cVar2S9S81P068P018P037nsss(0)='1'  OR cVar2S10S81P054P057P050nsss(0)='1'  OR cVar2S11S81N054P053nsss(0)='1'  )then
          oVar1S589(0) <='1';
          else
          oVar1S589(0) <='0';
          end if;
        if(cVar2S12S81N054N053P052nsss(0)='1'  OR cVar2S13S81P010P052nsss(0)='1'  OR cVar2S14S81P010N052P054nsss(0)='1'  OR cVar2S15S81N010P009nsss(0)='1'  )then
          oVar1S590(0) <='1';
          else
          oVar1S590(0) <='0';
          end if;
        if(cVar2S16S81N010N009P013nsss(0)='1'  OR cVar2S17S81P025P008nsss(0)='1'  OR cVar2S18S81N025P027nsss(0)='1'  OR cVar2S19S81N025N027P023nsss(0)='1'  )then
          oVar1S591(0) <='1';
          else
          oVar1S591(0) <='0';
          end if;
        if(cVar2S20S81P062P026P027nsss(0)='1'  OR cVar2S21S81P062P026P068nsss(0)='1'  OR cVar2S22S81N062P015P067nsss(0)='1'  )then
          oVar1S592(0) <='1';
          else
          oVar1S592(0) <='0';
          end if;
        if(cVar2S0S82P066nsss(0)='1'  OR cVar2S1S82P048nsss(0)='1'  OR cVar2S2S82P018P014nsss(0)='1'  OR cVar2S3S82P018P014nsss(0)='1'  )then
          oVar1S593(0) <='1';
          else
          oVar1S593(0) <='0';
          end if;
        if(cVar2S4S82P049P026nsss(0)='1'  OR cVar2S5S82P049N026P019nsss(0)='1'  OR cVar2S6S82N049P023P015nsss(0)='1'  OR cVar2S7S82N049N023P012nsss(0)='1'  )then
          oVar1S594(0) <='1';
          else
          oVar1S594(0) <='0';
          end if;
        if(cVar2S8S82P021P002nsss(0)='1'  OR cVar2S9S82P021N002P003nsss(0)='1'  OR cVar2S10S82N021P064nsss(0)='1'  OR cVar2S11S82P012P059P030nsss(0)='1'  )then
          oVar1S595(0) <='1';
          else
          oVar1S595(0) <='0';
          end if;
        if(cVar2S12S82P012N059P060nsss(0)='1'  OR cVar2S13S82N012P014nsss(0)='1'  OR cVar2S14S82N012N014P013nsss(0)='1'  OR cVar2S15S82P036nsss(0)='1'  )then
          oVar1S596(0) <='1';
          else
          oVar1S596(0) <='0';
          end if;
        if(cVar2S16S82P058P035nsss(0)='1'  OR cVar2S17S82P058P035P017nsss(0)='1'  OR cVar2S18S82N058P059P010nsss(0)='1'  OR cVar2S19S82P018nsss(0)='1'  )then
          oVar1S597(0) <='1';
          else
          oVar1S597(0) <='0';
          end if;
        if(cVar2S20S82N018P014nsss(0)='1'  OR cVar2S21S82P055P027P065nsss(0)='1'  OR cVar2S22S82P055P068nsss(0)='1'  OR cVar2S23S82P015P011nsss(0)='1'  )then
          oVar1S598(0) <='1';
          else
          oVar1S598(0) <='0';
          end if;
        if(cVar1S24S82P062P026P037P019nsss(0)='1'  )then
          oVar1S599(0) <='1';
          else
          oVar1S599(0) <='0';
          end if;
        if(cVar1S0S83P007P025P046P011nsss(0)='1'  OR cVar2S1S83P043nsss(0)='1'  OR cVar2S2S83N043P042nsss(0)='1'  OR cVar2S3S83N043N042P049nsss(0)='1'  )then
          oVar1S600(0) <='1';
          else
          oVar1S600(0) <='0';
          end if;
        if(cVar2S4S83P066P027P011nsss(0)='1'  OR cVar2S5S83P066N027psss(0)='1'  OR cVar2S6S83P066P019P014nsss(0)='1'  OR cVar2S7S83P066nsss(0)='1'  )then
          oVar1S601(0) <='1';
          else
          oVar1S601(0) <='0';
          end if;
        if(cVar2S8S83N066P035nsss(0)='1'  OR cVar2S9S83P062P013nsss(0)='1'  OR cVar2S10S83P009nsss(0)='1'  OR cVar1S11S83N007P040P002nsss(0)='1'  )then
          oVar1S602(0) <='1';
          else
          oVar1S602(0) <='0';
          end if;
        if(cVar1S12S83N007P040N002P047nsss(0)='1'  OR cVar2S13S83P039nsss(0)='1'  OR cVar2S14S83N039P004nsss(0)='1'  OR cVar2S15S83N039N004P000nsss(0)='1'  )then
          oVar1S603(0) <='1';
          else
          oVar1S603(0) <='0';
          end if;
        if(cVar2S16S83P062P029P035nsss(0)='1'  OR cVar2S17S83P062N029P006nsss(0)='1'  OR cVar2S18S83P014P033nsss(0)='1'  OR cVar2S19S83N014P064P059nsss(0)='1'  )then
          oVar1S604(0) <='1';
          else
          oVar1S604(0) <='0';
          end if;
        if(cVar2S20S83P001P003P050nsss(0)='1'  OR cVar2S21S83P001P003P039nsss(0)='1'  OR cVar2S22S83P001P039nsss(0)='1'  OR cVar2S23S83P001N039P010nsss(0)='1'  )then
          oVar1S605(0) <='1';
          else
          oVar1S605(0) <='0';
          end if;
        if(cVar1S0S84P040P021P002nsss(0)='1'  OR cVar2S1S84P003nsss(0)='1'  OR cVar2S2S84N003P004nsss(0)='1'  OR cVar2S3S84N003N004P005nsss(0)='1'  )then
          oVar1S607(0) <='1';
          else
          oVar1S607(0) <='0';
          end if;
        if(cVar1S4S84P040N021P057nsss(0)='1'  OR cVar2S5S84P039nsss(0)='1'  OR cVar2S6S84N039P060nsss(0)='1'  OR cVar2S7S84N039N060P009nsss(0)='1'  )then
          oVar1S608(0) <='1';
          else
          oVar1S608(0) <='0';
          end if;
        if(cVar2S8S84P011nsss(0)='1'  OR cVar2S9S84P047nsss(0)='1'  OR cVar2S10S84N047P042nsss(0)='1'  OR cVar2S11S84N047N042P043nsss(0)='1'  )then
          oVar1S609(0) <='1';
          else
          oVar1S609(0) <='0';
          end if;
        if(cVar2S12S84P011nsss(0)='1'  OR cVar2S13S84P011P015P012nsss(0)='1'  OR cVar2S14S84P011N015P012nsss(0)='1'  OR cVar2S15S84P010nsss(0)='1'  )then
          oVar1S610(0) <='1';
          else
          oVar1S610(0) <='0';
          end if;
        if(cVar2S16S84P003P020P039nsss(0)='1'  OR cVar2S17S84P003P020P002nsss(0)='1'  OR cVar2S18S84P003P020nsss(0)='1'  OR cVar2S19S84P039nsss(0)='1'  )then
          oVar1S611(0) <='1';
          else
          oVar1S611(0) <='0';
          end if;
        if(cVar2S20S84N039P003nsss(0)='1'  OR cVar2S21S84N039N003P066nsss(0)='1'  OR cVar2S22S84P065P058nsss(0)='1'  OR cVar2S23S84N065P017P068nsss(0)='1'  )then
          oVar1S612(0) <='1';
          else
          oVar1S612(0) <='0';
          end if;
        if(cVar2S24S84N065P017P018nsss(0)='1'  OR cVar2S25S84P029P051nsss(0)='1'  OR cVar2S26S84P029N051P028nsss(0)='1'  OR cVar2S27S84N029P067nsss(0)='1'  )then
          oVar1S613(0) <='1';
          else
          oVar1S613(0) <='0';
          end if;
        if(cVar2S28S84N029N067P026nsss(0)='1'  )then
          oVar1S614(0) <='1';
          else
          oVar1S614(0) <='0';
          end if;
        if(cVar1S0S85P015P032P005nsss(0)='1'  OR cVar2S1S85P011P012nsss(0)='1'  OR cVar2S2S85P011P012P058nsss(0)='1'  OR cVar2S3S85P021nsss(0)='1'  )then
          oVar1S615(0) <='1';
          else
          oVar1S615(0) <='0';
          end if;
        if(cVar2S4S85P018P019nsss(0)='1'  OR cVar2S5S85P010nsss(0)='1'  OR cVar2S6S85N010P037nsss(0)='1'  OR cVar2S7S85N010N037P019nsss(0)='1'  )then
          oVar1S616(0) <='1';
          else
          oVar1S616(0) <='0';
          end if;
        if(cVar2S8S85P038P054P036nsss(0)='1'  OR cVar2S9S85P038P002nsss(0)='1'  OR cVar1S10S85N015P021P038nsss(0)='1'  OR cVar2S11S85P042nsss(0)='1'  )then
          oVar1S617(0) <='1';
          else
          oVar1S617(0) <='0';
          end if;
        if(cVar2S12S85N042P037nsss(0)='1'  OR cVar2S13S85N042N037P039nsss(0)='1'  OR cVar2S14S85P016P018nsss(0)='1'  OR cVar1S15S85N015N021P044P004nsss(0)='1'  )then
          oVar1S618(0) <='1';
          else
          oVar1S618(0) <='0';
          end if;
        if(cVar2S16S85P025P017nsss(0)='1'  OR cVar2S17S85N025P005nsss(0)='1'  OR cVar2S18S85N025N005P043nsss(0)='1'  OR cVar2S19S85P013P056nsss(0)='1'  )then
          oVar1S619(0) <='1';
          else
          oVar1S619(0) <='0';
          end if;
        if(cVar2S20S85P013N056P060nsss(0)='1'  OR cVar2S21S85N013P057P011nsss(0)='1'  OR cVar2S22S85P049nsss(0)='1'  OR cVar2S23S85N049P043P019nsss(0)='1'  )then
          oVar1S620(0) <='1';
          else
          oVar1S620(0) <='0';
          end if;
        if(cVar1S0S86P021P038P002nsss(0)='1'  OR cVar1S1S86P021P038N002P004nsss(0)='1'  OR cVar2S2S86P003nsss(0)='1'  OR cVar2S3S86N003P005nsss(0)='1'  )then
          oVar1S622(0) <='1';
          else
          oVar1S622(0) <='0';
          end if;
        if(cVar1S4S86P021N038P010P042nsss(0)='1'  OR cVar2S5S86P011nsss(0)='1'  OR cVar1S6S86P021N038P010P019nsss(0)='1'  OR cVar1S7S86N021P020P039P003nsss(0)='1'  )then
          oVar1S623(0) <='1';
          else
          oVar1S623(0) <='0';
          end if;
        if(cVar2S8S86P002nsss(0)='1'  OR cVar2S9S86N002P005nsss(0)='1'  OR cVar2S10S86N002N005P004nsss(0)='1'  OR cVar2S11S86P013P066nsss(0)='1'  )then
          oVar1S624(0) <='1';
          else
          oVar1S624(0) <='0';
          end if;
        if(cVar2S12S86P013N066P018nsss(0)='1'  OR cVar2S13S86N013P003nsss(0)='1'  OR cVar2S14S86N013N003P053nsss(0)='1'  OR cVar2S15S86P014P055P019nsss(0)='1'  )then
          oVar1S625(0) <='1';
          else
          oVar1S625(0) <='0';
          end if;
        if(cVar2S16S86P014N055P011nsss(0)='1'  OR cVar2S17S86P014P005nsss(0)='1'  OR cVar2S18S86P005nsss(0)='1'  OR cVar2S19S86P005P049nsss(0)='1'  )then
          oVar1S626(0) <='1';
          else
          oVar1S626(0) <='0';
          end if;
        if(cVar2S20S86P005N049P023nsss(0)='1'  OR cVar2S21S86P019nsss(0)='1'  OR cVar2S22S86N019P010nsss(0)='1'  OR cVar2S23S86P006P015nsss(0)='1'  )then
          oVar1S627(0) <='1';
          else
          oVar1S627(0) <='0';
          end if;
        if(cVar2S24S86N006P055P024nsss(0)='1'  )then
          oVar1S628(0) <='1';
          else
          oVar1S628(0) <='0';
          end if;
        if(cVar1S0S87P015P055P061P032nsss(0)='1'  OR cVar2S1S87P067nsss(0)='1'  OR cVar2S2S87N067P019P056nsss(0)='1'  OR cVar2S3S87N067P019P010nsss(0)='1'  )then
          oVar1S629(0) <='1';
          else
          oVar1S629(0) <='0';
          end if;
        if(cVar2S4S87P033P039nsss(0)='1'  OR cVar2S5S87P033N039P019nsss(0)='1'  OR cVar2S6S87P039P007P056nsss(0)='1'  OR cVar2S7S87P039N007psss(0)='1'  )then
          oVar1S630(0) <='1';
          else
          oVar1S630(0) <='0';
          end if;
        if(cVar2S8S87P039P017nsss(0)='1'  OR cVar1S9S87P015N055P021P066nsss(0)='1'  OR cVar2S10S87P014P016nsss(0)='1'  OR cVar2S11S87N014P018nsss(0)='1'  )then
          oVar1S631(0) <='1';
          else
          oVar1S631(0) <='0';
          end if;
        if(cVar1S12S87N015P021P038nsss(0)='1'  OR cVar2S13S87P042P002nsss(0)='1'  OR cVar2S14S87P042N002P041nsss(0)='1'  OR cVar2S15S87N042P003nsss(0)='1'  )then
          oVar1S632(0) <='1';
          else
          oVar1S632(0) <='0';
          end if;
        if(cVar2S16S87N042N003P009nsss(0)='1'  OR cVar2S17S87P016P018nsss(0)='1'  OR cVar1S18S87N015N021P020P039nsss(0)='1'  OR cVar2S19S87P035P013nsss(0)='1'  )then
          oVar1S633(0) <='1';
          else
          oVar1S633(0) <='0';
          end if;
        if(cVar2S20S87P035N013P003nsss(0)='1'  OR cVar2S21S87P055P026P049nsss(0)='1'  OR cVar2S22S87P055P069nsss(0)='1'  OR cVar2S23S87P055N069P010nsss(0)='1'  )then
          oVar1S634(0) <='1';
          else
          oVar1S634(0) <='0';
          end if;
        if(cVar2S24S87P030P010nsss(0)='1'  OR cVar2S25S87P030N010P054nsss(0)='1'  OR cVar2S26S87N030P011P055nsss(0)='1'  OR cVar2S27S87N030N011P013nsss(0)='1'  )then
          oVar1S635(0) <='1';
          else
          oVar1S635(0) <='0';
          end if;
        if(cVar2S0S88P034P020nsss(0)='1'  OR cVar2S1S88P034N020P017nsss(0)='1'  OR cVar2S2S88P035P003P066nsss(0)='1'  OR cVar2S3S88P035N003psss(0)='1'  )then
          oVar1S637(0) <='1';
          else
          oVar1S637(0) <='0';
          end if;
        if(cVar2S4S88P035P017nsss(0)='1'  OR cVar2S5S88P035N017P014nsss(0)='1'  OR cVar1S6S88P015P057P055P069nsss(0)='1'  OR cVar2S7S88P053P010nsss(0)='1'  )then
          oVar1S638(0) <='1';
          else
          oVar1S638(0) <='0';
          end if;
        if(cVar2S8S88P053N010P051nsss(0)='1'  OR cVar2S9S88N053P063nsss(0)='1'  OR cVar2S10S88P036P012nsss(0)='1'  OR cVar2S11S88P036P012P030nsss(0)='1'  )then
          oVar1S639(0) <='1';
          else
          oVar1S639(0) <='0';
          end if;
        if(cVar2S12S88P031P017nsss(0)='1'  OR cVar2S13S88N031P030nsss(0)='1'  OR cVar2S14S88P068P019nsss(0)='1'  OR cVar2S15S88P068N019P037nsss(0)='1'  )then
          oVar1S640(0) <='1';
          else
          oVar1S640(0) <='0';
          end if;
        if(cVar2S16S88N068P012P065nsss(0)='1'  OR cVar2S17S88N068N012P011nsss(0)='1'  OR cVar1S18S88P015P055P061P032nsss(0)='1'  OR cVar2S19S88P057nsss(0)='1'  )then
          oVar1S641(0) <='1';
          else
          oVar1S641(0) <='0';
          end if;
        if(cVar2S20S88N057P017nsss(0)='1'  OR cVar1S21S88P015N055P020P002nsss(0)='1'  OR cVar2S22S88P033P007P019nsss(0)='1'  OR cVar2S23S88P024P005P013nsss(0)='1'  )then
          oVar1S642(0) <='1';
          else
          oVar1S642(0) <='0';
          end if;
        if(cVar2S24S88P024N005psss(0)='1'  OR cVar2S25S88P039P007nsss(0)='1'  OR cVar2S26S88P039P017nsss(0)='1'  )then
          oVar1S643(0) <='1';
          else
          oVar1S643(0) <='0';
          end if;
        if(cVar2S0S89P033nsss(0)='1'  OR cVar2S1S89N033P037P019nsss(0)='1'  OR cVar2S2S89N033P037P018nsss(0)='1'  OR cVar2S3S89P012P033P046nsss(0)='1'  )then
          oVar1S644(0) <='1';
          else
          oVar1S644(0) <='0';
          end if;
        if(cVar2S4S89N012P032P033nsss(0)='1'  OR cVar2S5S89N012N032P035nsss(0)='1'  OR cVar2S6S89P063nsss(0)='1'  OR cVar2S7S89N063P035P014nsss(0)='1'  )then
          oVar1S645(0) <='1';
          else
          oVar1S645(0) <='0';
          end if;
        if(cVar2S8S89P052nsss(0)='1'  OR cVar2S9S89P057nsss(0)='1'  OR cVar2S10S89P005P019nsss(0)='1'  OR cVar2S11S89P005P019P014nsss(0)='1'  )then
          oVar1S646(0) <='1';
          else
          oVar1S646(0) <='0';
          end if;
        if(cVar2S12S89N005P019P018nsss(0)='1'  OR cVar2S13S89N005N019P068nsss(0)='1'  OR cVar2S14S89P058nsss(0)='1'  OR cVar2S15S89N058P032nsss(0)='1'  )then
          oVar1S647(0) <='1';
          else
          oVar1S647(0) <='0';
          end if;
        if(cVar1S16S89N015P039P020P003nsss(0)='1'  OR cVar2S17S89P002nsss(0)='1'  OR cVar2S18S89N002P005nsss(0)='1'  OR cVar2S19S89P021nsss(0)='1'  )then
          oVar1S648(0) <='1';
          else
          oVar1S648(0) <='0';
          end if;
        if(cVar2S20S89N021P011nsss(0)='1'  OR cVar2S21S89P017P014nsss(0)='1'  OR cVar2S22S89P005P023nsss(0)='1'  OR cVar2S23S89N005P004P042nsss(0)='1'  )then
          oVar1S649(0) <='1';
          else
          oVar1S649(0) <='0';
          end if;
        if(cVar2S24S89N005N004P006nsss(0)='1'  OR cVar2S25S89P021nsss(0)='1'  OR cVar2S26S89N021P017P012nsss(0)='1'  OR cVar2S27S89P027P009nsss(0)='1'  )then
          oVar1S650(0) <='1';
          else
          oVar1S650(0) <='0';
          end if;
        if(cVar2S28S89P027N009P037nsss(0)='1'  OR cVar2S29S89N027P042P064nsss(0)='1'  )then
          oVar1S651(0) <='1';
          else
          oVar1S651(0) <='0';
          end if;
        if(cVar1S0S90P020P039P010P003nsss(0)='1'  OR cVar2S1S90P041nsss(0)='1'  OR cVar1S2S90P020N039P025nsss(0)='1'  OR cVar2S3S90P050P024nsss(0)='1'  )then
          oVar1S652(0) <='1';
          else
          oVar1S652(0) <='0';
          end if;
        if(cVar2S4S90P050N024P051nsss(0)='1'  OR cVar1S5S90N020P040P021P002nsss(0)='1'  OR cVar2S6S90P018nsss(0)='1'  OR cVar2S7S90N018P004nsss(0)='1'  )then
          oVar1S653(0) <='1';
          else
          oVar1S653(0) <='0';
          end if;
        if(cVar2S8S90N018N004P003nsss(0)='1'  OR cVar1S9S90N020P040N021P057nsss(0)='1'  OR cVar2S10S90P003P009P042nsss(0)='1'  OR cVar2S11S90P043P065nsss(0)='1'  )then
          oVar1S654(0) <='1';
          else
          oVar1S654(0) <='0';
          end if;
        if(cVar2S12S90N043P048nsss(0)='1'  OR cVar2S13S90N043N048P060nsss(0)='1'  OR cVar2S14S90P015P013P025nsss(0)='1'  OR cVar2S15S90P015P013P059nsss(0)='1'  )then
          oVar1S655(0) <='1';
          else
          oVar1S655(0) <='0';
          end if;
        if(cVar2S16S90N015P057P055nsss(0)='1'  OR cVar2S17S90N015P057P010nsss(0)='1'  OR cVar1S18S90N020N040P039P005nsss(0)='1'  )then
          oVar1S656(0) <='1';
          else
          oVar1S656(0) <='0';
          end if;
        if(cVar1S0S91P020P039P010P003nsss(0)='1'  OR cVar2S1S91P041nsss(0)='1'  OR cVar1S2S91P020N039P025nsss(0)='1'  OR cVar1S3S91P020N039N025P024nsss(0)='1'  )then
          oVar1S657(0) <='1';
          else
          oVar1S657(0) <='0';
          end if;
        if(cVar2S4S91P053nsss(0)='1'  OR cVar2S5S91N053P069P032nsss(0)='1'  OR cVar1S6S91N020P045P004P018nsss(0)='1'  OR cVar2S7S91P022nsss(0)='1'  )then
          oVar1S658(0) <='1';
          else
          oVar1S658(0) <='0';
          end if;
        if(cVar2S8S91P024nsss(0)='1'  OR cVar2S9S91N024P022nsss(0)='1'  OR cVar2S10S91P007nsss(0)='1'  OR cVar2S11S91N007P051nsss(0)='1'  )then
          oVar1S659(0) <='1';
          else
          oVar1S659(0) <='0';
          end if;
        if(cVar2S12S91N007N051P014nsss(0)='1'  OR cVar1S13S91N020N045P040P021nsss(0)='1'  OR cVar2S14S91P054nsss(0)='1'  OR cVar2S15S91N054P003P014nsss(0)='1'  )then
          oVar1S660(0) <='1';
          else
          oVar1S660(0) <='0';
          end if;
        if(cVar2S16S91P010P028P012nsss(0)='1'  OR cVar2S17S91P010N028P030nsss(0)='1'  OR cVar2S18S91N010P067nsss(0)='1'  OR cVar2S19S91P057P043P065nsss(0)='1'  )then
          oVar1S661(0) <='1';
          else
          oVar1S661(0) <='0';
          end if;
        if(cVar2S20S91P057P059nsss(0)='1'  OR cVar2S21S91P057N059P068nsss(0)='1'  )then
          oVar1S662(0) <='1';
          else
          oVar1S662(0) <='0';
          end if;
        if(cVar1S0S92P020P039P010P003nsss(0)='1'  OR cVar2S1S92P002nsss(0)='1'  OR cVar2S2S92N002P019nsss(0)='1'  OR cVar1S3S92P020N039P025nsss(0)='1'  )then
          oVar1S663(0) <='1';
          else
          oVar1S663(0) <='0';
          end if;
        if(cVar2S4S92P035P029nsss(0)='1'  OR cVar2S5S92P035P014nsss(0)='1'  OR cVar1S6S92N020P045P004P018nsss(0)='1'  OR cVar2S7S92P022nsss(0)='1'  )then
          oVar1S664(0) <='1';
          else
          oVar1S664(0) <='0';
          end if;
        if(cVar2S8S92P024nsss(0)='1'  OR cVar2S9S92N024P022nsss(0)='1'  OR cVar2S10S92P007nsss(0)='1'  OR cVar2S11S92N007P051nsss(0)='1'  )then
          oVar1S665(0) <='1';
          else
          oVar1S665(0) <='0';
          end if;
        if(cVar2S12S92N007N051P014nsss(0)='1'  OR cVar1S13S92N020N045P040P021nsss(0)='1'  OR cVar2S14S92P003P052nsss(0)='1'  OR cVar2S15S92P003N052P023nsss(0)='1'  )then
          oVar1S666(0) <='1';
          else
          oVar1S666(0) <='0';
          end if;
        if(cVar2S16S92P006P048nsss(0)='1'  OR cVar2S17S92N006P002nsss(0)='1'  OR cVar2S18S92N006N002P007nsss(0)='1'  OR cVar2S19S92P042P023P002nsss(0)='1'  )then
          oVar1S667(0) <='1';
          else
          oVar1S667(0) <='0';
          end if;
        if(cVar2S20S92P042P023P041nsss(0)='1'  OR cVar2S21S92P042P064nsss(0)='1'  OR cVar2S22S92P042N064P035nsss(0)='1'  )then
          oVar1S668(0) <='1';
          else
          oVar1S668(0) <='0';
          end if;
        if(cVar1S0S93P040P002P021nsss(0)='1'  OR cVar1S1S93P040P002N021P041nsss(0)='1'  OR cVar2S2S93P038nsss(0)='1'  OR cVar1S3S93P040N002P004P022nsss(0)='1'  )then
          oVar1S669(0) <='1';
          else
          oVar1S669(0) <='0';
          end if;
        if(cVar2S4S93P023nsss(0)='1'  OR cVar2S5S93N023P038nsss(0)='1'  OR cVar1S6S93P040N002N004P000nsss(0)='1'  OR cVar2S7S93P057nsss(0)='1'  )then
          oVar1S670(0) <='1';
          else
          oVar1S670(0) <='0';
          end if;
        if(cVar2S8S93N057P050nsss(0)='1'  OR cVar2S9S93N057N050P005nsss(0)='1'  OR cVar1S10S93N040P045P022P019nsss(0)='1'  OR cVar2S11S93P014nsss(0)='1'  )then
          oVar1S671(0) <='1';
          else
          oVar1S671(0) <='0';
          end if;
        if(cVar2S12S93N014P007nsss(0)='1'  OR cVar2S13S93N014N007P004nsss(0)='1'  OR cVar2S14S93P017nsss(0)='1'  OR cVar2S15S93P027P006P024nsss(0)='1'  )then
          oVar1S672(0) <='1';
          else
          oVar1S672(0) <='0';
          end if;
        if(cVar2S16S93P027N006P003nsss(0)='1'  OR cVar2S17S93P003nsss(0)='1'  OR cVar2S18S93N003P002nsss(0)='1'  OR cVar2S19S93N003N002P005nsss(0)='1'  )then
          oVar1S673(0) <='1';
          else
          oVar1S673(0) <='0';
          end if;
        if(cVar2S20S93P004P010nsss(0)='1'  OR cVar2S21S93P004N010P048nsss(0)='1'  OR cVar2S22S93P006P048nsss(0)='1'  OR cVar2S23S93N006P004P042nsss(0)='1'  )then
          oVar1S674(0) <='1';
          else
          oVar1S674(0) <='0';
          end if;
        if(cVar2S24S93N006N004P005nsss(0)='1'  OR cVar2S25S93P042P004P028nsss(0)='1'  OR cVar2S26S93P042P004P005nsss(0)='1'  OR cVar2S27S93P042P064nsss(0)='1'  )then
          oVar1S675(0) <='1';
          else
          oVar1S675(0) <='0';
          end if;
        if(cVar2S28S93P042N064P035nsss(0)='1'  )then
          oVar1S676(0) <='1';
          else
          oVar1S676(0) <='0';
          end if;
        if(cVar1S0S94P040P002P021nsss(0)='1'  OR cVar1S1S94P040P002N021P041nsss(0)='1'  OR cVar2S2S94P038nsss(0)='1'  OR cVar1S3S94P040N002P004P022nsss(0)='1'  )then
          oVar1S677(0) <='1';
          else
          oVar1S677(0) <='0';
          end if;
        if(cVar2S4S94P023nsss(0)='1'  OR cVar2S5S94N023P038nsss(0)='1'  OR cVar1S6S94P040N002N004P020nsss(0)='1'  OR cVar2S7S94P042nsss(0)='1'  )then
          oVar1S678(0) <='1';
          else
          oVar1S678(0) <='0';
          end if;
        if(cVar2S8S94N042P025nsss(0)='1'  OR cVar2S9S94P005nsss(0)='1'  OR cVar2S10S94N005P004nsss(0)='1'  OR cVar2S11S94N005N004P007nsss(0)='1'  )then
          oVar1S679(0) <='1';
          else
          oVar1S679(0) <='0';
          end if;
        if(cVar2S12S94P051nsss(0)='1'  OR cVar2S13S94N051P002nsss(0)='1'  OR cVar2S14S94N051N002P043nsss(0)='1'  OR cVar2S15S94P039nsss(0)='1'  )then
          oVar1S680(0) <='1';
          else
          oVar1S680(0) <='0';
          end if;
        if(cVar2S16S94N039P004nsss(0)='1'  OR cVar2S17S94P045P006nsss(0)='1'  OR cVar2S18S94P045N006P022nsss(0)='1'  OR cVar2S19S94N045P004nsss(0)='1'  )then
          oVar1S681(0) <='1';
          else
          oVar1S681(0) <='0';
          end if;
        if(cVar2S20S94N045P004P019nsss(0)='1'  OR cVar1S21S94N040N044P042P058nsss(0)='1'  OR cVar2S22S94P069nsss(0)='1'  OR cVar2S23S94N069P043nsss(0)='1'  )then
          oVar1S682(0) <='1';
          else
          oVar1S682(0) <='0';
          end if;
        if(cVar1S0S95P044P023P005nsss(0)='1'  OR cVar1S1S95P044P023N005P004nsss(0)='1'  OR cVar2S2S95P007nsss(0)='1'  OR cVar2S3S95N007P006nsss(0)='1'  )then
          oVar1S684(0) <='1';
          else
          oVar1S684(0) <='0';
          end if;
        if(cVar1S4S95P044N023P051nsss(0)='1'  OR cVar1S5S95P044N023N051P057nsss(0)='1'  OR cVar2S6S95P006P022nsss(0)='1'  OR cVar2S7S95P006N022P024nsss(0)='1'  )then
          oVar1S685(0) <='1';
          else
          oVar1S685(0) <='0';
          end if;
        if(cVar2S8S95N006P060nsss(0)='1'  OR cVar2S9S95N006N060P054nsss(0)='1'  OR cVar1S10S95N044P040P002nsss(0)='1'  OR cVar2S11S95P023nsss(0)='1'  )then
          oVar1S686(0) <='1';
          else
          oVar1S686(0) <='0';
          end if;
        if(cVar2S12S95N023P022nsss(0)='1'  OR cVar2S13S95N023N022P038nsss(0)='1'  OR cVar2S14S95P000nsss(0)='1'  OR cVar2S15S95N000P039nsss(0)='1'  )then
          oVar1S687(0) <='1';
          else
          oVar1S687(0) <='0';
          end if;
        if(cVar2S16S95N000N039P012nsss(0)='1'  OR cVar1S17S95N044N040P045P022nsss(0)='1'  OR cVar2S18S95P023P017nsss(0)='1'  OR cVar2S19S95N023P006P024nsss(0)='1'  )then
          oVar1S688(0) <='1';
          else
          oVar1S688(0) <='0';
          end if;
        if(cVar2S20S95N023N006P067nsss(0)='1'  OR cVar2S21S95P039P003nsss(0)='1'  OR cVar2S22S95P039N003P002nsss(0)='1'  OR cVar2S23S95N039P048nsss(0)='1'  )then
          oVar1S689(0) <='1';
          else
          oVar1S689(0) <='0';
          end if;
        if(cVar2S24S95N039N048P004nsss(0)='1'  OR cVar2S25S95P042P016P033nsss(0)='1'  OR cVar2S26S95P042N016P033nsss(0)='1'  OR cVar2S27S95P042P064nsss(0)='1'  )then
          oVar1S690(0) <='1';
          else
          oVar1S690(0) <='0';
          end if;
        if(cVar2S28S95P042N064P035nsss(0)='1'  )then
          oVar1S691(0) <='1';
          else
          oVar1S691(0) <='0';
          end if;
        if(cVar1S0S96P044P004P023nsss(0)='1'  OR cVar2S1S96P019nsss(0)='1'  OR cVar1S2S96P044N004P021nsss(0)='1'  OR cVar2S3S96P023nsss(0)='1'  )then
          oVar1S692(0) <='1';
          else
          oVar1S692(0) <='0';
          end if;
        if(cVar2S4S96P006P024nsss(0)='1'  OR cVar2S5S96P006N024P025nsss(0)='1'  OR cVar2S6S96N006P007nsss(0)='1'  OR cVar2S7S96N006N007P050nsss(0)='1'  )then
          oVar1S693(0) <='1';
          else
          oVar1S693(0) <='0';
          end if;
        if(cVar2S8S96P030nsss(0)='1'  OR cVar2S9S96N030P065P031nsss(0)='1'  OR cVar2S10S96P067P065nsss(0)='1'  OR cVar2S11S96P067P065P009nsss(0)='1'  )then
          oVar1S694(0) <='1';
          else
          oVar1S694(0) <='0';
          end if;
        if(cVar2S12S96P067P034nsss(0)='1'  OR cVar2S13S96P067N034P062nsss(0)='1'  OR cVar2S14S96P028P015P018nsss(0)='1'  OR cVar2S15S96N028P066nsss(0)='1'  )then
          oVar1S695(0) <='1';
          else
          oVar1S695(0) <='0';
          end if;
        if(cVar2S16S96P030nsss(0)='1'  OR cVar2S17S96P030P031P010nsss(0)='1'  OR cVar2S18S96P047P053P003nsss(0)='1'  OR cVar2S19S96P047P066nsss(0)='1'  )then
          oVar1S696(0) <='1';
          else
          oVar1S696(0) <='0';
          end if;
        if(cVar2S20S96P047N066P026nsss(0)='1'  OR cVar2S21S96P062P060nsss(0)='1'  OR cVar2S22S96P062N060P034nsss(0)='1'  OR cVar2S23S96N062P058P018nsss(0)='1'  )then
          oVar1S697(0) <='1';
          else
          oVar1S697(0) <='0';
          end if;
        if(cVar1S24S96N044P016P052P065nsss(0)='1'  OR cVar2S25S96P007P010P050nsss(0)='1'  OR cVar2S26S96P007N010P008nsss(0)='1'  )then
          oVar1S698(0) <='1';
          else
          oVar1S698(0) <='0';
          end if;
        if(cVar1S0S97P044P004P023nsss(0)='1'  OR cVar2S1S97P019nsss(0)='1'  OR cVar1S2S97P044N004P021nsss(0)='1'  OR cVar2S3S97P023nsss(0)='1'  )then
          oVar1S699(0) <='1';
          else
          oVar1S699(0) <='0';
          end if;
        if(cVar2S4S97N023P025nsss(0)='1'  OR cVar2S5S97P057nsss(0)='1'  OR cVar2S6S97N057P006nsss(0)='1'  OR cVar2S7S97N057N006P066nsss(0)='1'  )then
          oVar1S700(0) <='1';
          else
          oVar1S700(0) <='0';
          end if;
        if(cVar2S8S97P047P053P028nsss(0)='1'  OR cVar2S9S97P047P066nsss(0)='1'  OR cVar2S10S97P047N066P026nsss(0)='1'  OR cVar2S11S97P065P058P014nsss(0)='1'  )then
          oVar1S701(0) <='1';
          else
          oVar1S701(0) <='0';
          end if;
        if(cVar2S12S97P065P058P018nsss(0)='1'  OR cVar2S13S97P065P063P064nsss(0)='1'  OR cVar1S14S97N044P016P052P065nsss(0)='1'  OR cVar2S15S97P007P010P050nsss(0)='1'  )then
          oVar1S702(0) <='1';
          else
          oVar1S702(0) <='0';
          end if;
        if(cVar2S16S97P030nsss(0)='1'  OR cVar2S17S97N030P065P031nsss(0)='1'  OR cVar2S18S97P032P014P066nsss(0)='1'  OR cVar2S19S97P032P014P019nsss(0)='1'  )then
          oVar1S703(0) <='1';
          else
          oVar1S703(0) <='0';
          end if;
        if(cVar2S20S97N032P054P030nsss(0)='1'  OR cVar2S21S97P028P011nsss(0)='1'  OR cVar2S22S97P028N011P015nsss(0)='1'  OR cVar2S23S97N028P066nsss(0)='1'  )then
          oVar1S704(0) <='1';
          else
          oVar1S704(0) <='0';
          end if;
        if(cVar2S24S97P032P041nsss(0)='1'  OR cVar2S25S97P032N041P040nsss(0)='1'  OR cVar2S26S97P032P014P060nsss(0)='1'  )then
          oVar1S705(0) <='1';
          else
          oVar1S705(0) <='0';
          end if;
        if(cVar1S0S98P016P044P004P023nsss(0)='1'  OR cVar2S1S98P019nsss(0)='1'  OR cVar1S2S98P016P044N004P047nsss(0)='1'  OR cVar2S3S98P021nsss(0)='1'  )then
          oVar1S706(0) <='1';
          else
          oVar1S706(0) <='0';
          end if;
        if(cVar2S4S98N021P025nsss(0)='1'  OR cVar2S5S98N021N025P023nsss(0)='1'  OR cVar2S6S98P030nsss(0)='1'  OR cVar2S7S98N030P065nsss(0)='1'  )then
          oVar1S707(0) <='1';
          else
          oVar1S707(0) <='0';
          end if;
        if(cVar2S8S98P041P032P014nsss(0)='1'  OR cVar2S9S98P041N032psss(0)='1'  OR cVar2S10S98P041P018P020nsss(0)='1'  OR cVar2S11S98P050nsss(0)='1'  )then
          oVar1S708(0) <='1';
          else
          oVar1S708(0) <='0';
          end if;
        if(cVar2S12S98P050P014P052nsss(0)='1'  OR cVar2S13S98P050P014P027nsss(0)='1'  OR cVar2S14S98P014P060nsss(0)='1'  OR cVar2S15S98P014N060P059nsss(0)='1'  )then
          oVar1S709(0) <='1';
          else
          oVar1S709(0) <='0';
          end if;
        if(cVar2S16S98N014P058P007nsss(0)='1'  OR cVar1S17S98P016P021P037P053nsss(0)='1'  OR cVar2S18S98P020P002nsss(0)='1'  OR cVar2S19S98P002P009nsss(0)='1'  )then
          oVar1S710(0) <='1';
          else
          oVar1S710(0) <='0';
          end if;
        if(cVar2S20S98P002N009P018nsss(0)='1'  OR cVar2S21S98N002P045P006nsss(0)='1'  OR cVar2S22S98P006nsss(0)='1'  OR cVar2S23S98N006P018P049nsss(0)='1'  )then
          oVar1S711(0) <='1';
          else
          oVar1S711(0) <='0';
          end if;
        if(cVar2S24S98N006N018P007nsss(0)='1'  OR cVar1S25S98P016P021P069P038nsss(0)='1'  OR cVar2S26S98P015P019nsss(0)='1'  OR cVar2S27S98P015N019P018nsss(0)='1'  )then
          oVar1S712(0) <='1';
          else
          oVar1S712(0) <='0';
          end if;
        if(cVar1S0S99P044P051nsss(0)='1'  OR cVar1S1S99P044N051P057nsss(0)='1'  OR cVar1S2S99P044N051N057P032nsss(0)='1'  OR cVar2S3S99P004P023nsss(0)='1'  )then
          oVar1S714(0) <='1';
          else
          oVar1S714(0) <='0';
          end if;
        if(cVar2S4S99P004N023P022nsss(0)='1'  OR cVar2S5S99N004P021nsss(0)='1'  OR cVar2S6S99N004N021P038nsss(0)='1'  OR cVar2S7S99P020nsss(0)='1'  )then
          oVar1S715(0) <='1';
          else
          oVar1S715(0) <='0';
          end if;
        if(cVar2S8S99N020P021nsss(0)='1'  OR cVar2S9S99P066P035P052nsss(0)='1'  OR cVar2S10S99P066P035P016nsss(0)='1'  OR cVar2S11S99P066P058P011nsss(0)='1'  )then
          oVar1S716(0) <='1';
          else
          oVar1S716(0) <='0';
          end if;
        if(cVar2S12S99P008P026nsss(0)='1'  OR cVar2S13S99P008N026P028nsss(0)='1'  OR cVar2S14S99N008P047P015nsss(0)='1'  OR cVar2S15S99N008P047P006nsss(0)='1'  )then
          oVar1S717(0) <='1';
          else
          oVar1S717(0) <='0';
          end if;
        if(cVar2S16S99P023nsss(0)='1'  OR cVar2S17S99N023P039nsss(0)='1'  OR cVar2S18S99N023N039P002nsss(0)='1'  OR cVar1S19S99N044P062P063P053nsss(0)='1'  )then
          oVar1S718(0) <='1';
          else
          oVar1S718(0) <='0';
          end if;
        if(cVar2S20S99P056P060nsss(0)='1'  OR cVar2S21S99P056N060P003nsss(0)='1'  OR cVar2S22S99P056P031nsss(0)='1'  OR cVar2S23S99P056N031P035nsss(0)='1'  )then
          oVar1S719(0) <='1';
          else
          oVar1S719(0) <='0';
          end if;
        if(cVar2S24S99N056P011P034nsss(0)='1'  OR cVar2S25S99N056P011P017nsss(0)='1'  OR cVar2S26S99P033P066P037nsss(0)='1'  OR cVar2S27S99P033N066P019nsss(0)='1'  )then
          oVar1S720(0) <='1';
          else
          oVar1S720(0) <='0';
          end if;
        if(cVar1S0S100P015P044P004nsss(0)='1'  OR cVar1S1S100P015P044N004P021nsss(0)='1'  OR cVar2S2S100P025P017nsss(0)='1'  OR cVar2S3S100N025P005nsss(0)='1'  )then
          oVar1S722(0) <='1';
          else
          oVar1S722(0) <='0';
          end if;
        if(cVar2S4S100N025N005P013nsss(0)='1'  OR cVar1S5S100P015N044P062P045nsss(0)='1'  OR cVar2S6S100P034P039nsss(0)='1'  OR cVar2S7S100P034N039P005nsss(0)='1'  )then
          oVar1S723(0) <='1';
          else
          oVar1S723(0) <='0';
          end if;
        if(cVar2S8S100P034P014P033nsss(0)='1'  OR cVar2S9S100P012P061nsss(0)='1'  OR cVar2S10S100P012N061P036nsss(0)='1'  OR cVar2S11S100P012P036nsss(0)='1'  )then
          oVar1S724(0) <='1';
          else
          oVar1S724(0) <='0';
          end if;
        if(cVar2S12S100P012N036P013nsss(0)='1'  OR cVar2S13S100P016P014P064nsss(0)='1'  OR cVar2S14S100P016P014P018nsss(0)='1'  OR cVar2S15S100N016P014P034nsss(0)='1'  )then
          oVar1S725(0) <='1';
          else
          oVar1S725(0) <='0';
          end if;
        if(cVar2S16S100N016N014P019nsss(0)='1'  OR cVar2S17S100P012P057nsss(0)='1'  OR cVar2S18S100P012N057P018nsss(0)='1'  OR cVar2S19S100P068P066P014nsss(0)='1'  )then
          oVar1S726(0) <='1';
          else
          oVar1S726(0) <='0';
          end if;
        if(cVar2S20S100P068P066P062nsss(0)='1'  OR cVar2S21S100P068P066P062nsss(0)='1'  OR cVar2S22S100P014nsss(0)='1'  OR cVar2S23S100P011P019nsss(0)='1'  )then
          oVar1S727(0) <='1';
          else
          oVar1S727(0) <='0';
          end if;
        if(cVar1S24S100P015P013P025nsss(0)='1'  OR cVar2S25S100P035P037nsss(0)='1'  OR cVar2S26S100P035N037P009nsss(0)='1'  OR cVar2S27S100P035P017nsss(0)='1'  )then
          oVar1S728(0) <='1';
          else
          oVar1S728(0) <='0';
          end if;
        if(cVar2S28S100P024P019nsss(0)='1'  OR cVar2S29S100N024P031P011nsss(0)='1'  OR cVar2S30S100N024N031P010nsss(0)='1'  )then
          oVar1S729(0) <='1';
          else
          oVar1S729(0) <='0';
          end if;
        if(cVar2S0S101P021P038nsss(0)='1'  OR cVar2S1S101P021P014nsss(0)='1'  OR cVar2S2S101P066P067nsss(0)='1'  OR cVar2S3S101P066N067P012nsss(0)='1'  )then
          oVar1S730(0) <='1';
          else
          oVar1S730(0) <='0';
          end if;
        if(cVar2S4S101P066P017P065nsss(0)='1'  OR cVar2S5S101P066N017P036nsss(0)='1'  OR cVar1S6S101P015P013P056P050nsss(0)='1'  OR cVar2S7S101P014P029nsss(0)='1'  )then
          oVar1S731(0) <='1';
          else
          oVar1S731(0) <='0';
          end if;
        if(cVar2S8S101P014N029P016nsss(0)='1'  OR cVar1S9S101P015P013P025nsss(0)='1'  OR cVar2S10S101P052nsss(0)='1'  OR cVar2S11S101N052P027nsss(0)='1'  )then
          oVar1S732(0) <='1';
          else
          oVar1S732(0) <='0';
          end if;
        if(cVar2S12S101N052N027P008nsss(0)='1'  OR cVar2S13S101P012nsss(0)='1'  OR cVar2S14S101P014nsss(0)='1'  OR cVar1S15S101N015P044P025P017psss(0)='1'  )then
          oVar1S733(0) <='1';
          else
          oVar1S733(0) <='0';
          end if;
        if(cVar2S16S101P023nsss(0)='1'  OR cVar2S17S101P004P042nsss(0)='1'  OR cVar2S18S101N004P021nsss(0)='1'  OR cVar2S19S101N004N021P065nsss(0)='1'  )then
          oVar1S734(0) <='1';
          else
          oVar1S734(0) <='0';
          end if;
        if(cVar2S20S101P019P047P007nsss(0)='1'  OR cVar2S21S101P019P047P007nsss(0)='1'  OR cVar2S22S101P019P010P004nsss(0)='1'  OR cVar2S23S101P019P010P037nsss(0)='1'  )then
          oVar1S735(0) <='1';
          else
          oVar1S735(0) <='0';
          end if;
        if(cVar2S24S101P065nsss(0)='1'  OR cVar2S25S101P056P030nsss(0)='1'  OR cVar2S26S101P056N030P019nsss(0)='1'  OR cVar2S27S101N056P032P035nsss(0)='1'  )then
          oVar1S736(0) <='1';
          else
          oVar1S736(0) <='0';
          end if;
        if(cVar2S28S101N056N032P033nsss(0)='1'  OR cVar2S29S101P002P009nsss(0)='1'  OR cVar2S30S101N002P032P014nsss(0)='1'  )then
          oVar1S737(0) <='1';
          else
          oVar1S737(0) <='0';
          end if;
        if(cVar1S0S102P016P015P044nsss(0)='1'  OR cVar2S1S102P031P056nsss(0)='1'  OR cVar2S2S102P031N056P061nsss(0)='1'  OR cVar2S3S102N031P054nsss(0)='1'  )then
          oVar1S738(0) <='1';
          else
          oVar1S738(0) <='0';
          end if;
        if(cVar2S4S102N031P054P029nsss(0)='1'  OR cVar2S5S102P012P014P035nsss(0)='1'  OR cVar2S6S102P012P014P059nsss(0)='1'  OR cVar2S7S102N012P050nsss(0)='1'  )then
          oVar1S739(0) <='1';
          else
          oVar1S739(0) <='0';
          end if;
        if(cVar2S8S102P035P002P062nsss(0)='1'  OR cVar2S9S102N035P063P048nsss(0)='1'  OR cVar2S10S102N035P063P034nsss(0)='1'  OR cVar2S11S102P036P013nsss(0)='1'  )then
          oVar1S740(0) <='1';
          else
          oVar1S740(0) <='0';
          end if;
        if(cVar2S12S102P036P013P018nsss(0)='1'  OR cVar2S13S102N036P068P035nsss(0)='1'  OR cVar2S14S102N036N068P028nsss(0)='1'  OR cVar1S15S102P016P015P043P005nsss(0)='1'  )then
          oVar1S741(0) <='1';
          else
          oVar1S741(0) <='0';
          end if;
        if(cVar2S16S102P004nsss(0)='1'  OR cVar2S17S102P019nsss(0)='1'  OR cVar2S18S102N019P011P054nsss(0)='1'  OR cVar2S19S102P005nsss(0)='1'  )then
          oVar1S742(0) <='1';
          else
          oVar1S742(0) <='0';
          end if;
        if(cVar2S20S102N005P013P054nsss(0)='1'  OR cVar1S21S102P016P021P012P040nsss(0)='1'  OR cVar2S22S102P000P010nsss(0)='1'  OR cVar2S23S102P000N010P018nsss(0)='1'  )then
          oVar1S743(0) <='1';
          else
          oVar1S743(0) <='0';
          end if;
        if(cVar2S24S102N000P032P013nsss(0)='1'  OR cVar1S25S102P016P021P069P038nsss(0)='1'  OR cVar2S26S102P008nsss(0)='1'  OR cVar2S27S102N008P015P019nsss(0)='1'  )then
          oVar1S744(0) <='1';
          else
          oVar1S744(0) <='0';
          end if;
        if(cVar2S0S103P036nsss(0)='1'  OR cVar2S1S103P036P011P019nsss(0)='1'  OR cVar2S2S103P036N011P069nsss(0)='1'  OR cVar2S3S103P059P016nsss(0)='1'  )then
          oVar1S746(0) <='1';
          else
          oVar1S746(0) <='0';
          end if;
        if(cVar2S4S103N059P019P016nsss(0)='1'  OR cVar2S5S103P065P034nsss(0)='1'  OR cVar2S6S103P069P014nsss(0)='1'  OR cVar2S7S103P069N014P018nsss(0)='1'  )then
          oVar1S747(0) <='1';
          else
          oVar1S747(0) <='0';
          end if;
        if(cVar2S8S103N069P034P014nsss(0)='1'  OR cVar2S9S103P001P027nsss(0)='1'  OR cVar2S10S103P065P034nsss(0)='1'  OR cVar2S11S103P065N034P024nsss(0)='1'  )then
          oVar1S748(0) <='1';
          else
          oVar1S748(0) <='0';
          end if;
        if(cVar2S12S103P065P011P034nsss(0)='1'  OR cVar2S13S103P037nsss(0)='1'  OR cVar1S14S103N015P044P004P023nsss(0)='1'  OR cVar2S15S103P022nsss(0)='1'  )then
          oVar1S749(0) <='1';
          else
          oVar1S749(0) <='0';
          end if;
        if(cVar2S16S103P023nsss(0)='1'  OR cVar2S17S103N023P025nsss(0)='1'  OR cVar2S18S103P059nsss(0)='1'  OR cVar2S19S103N059P014nsss(0)='1'  )then
          oVar1S750(0) <='1';
          else
          oVar1S750(0) <='0';
          end if;
        if(cVar2S20S103N059P014P046nsss(0)='1'  OR cVar2S21S103P054nsss(0)='1'  OR cVar2S22S103N054P011nsss(0)='1'  OR cVar2S23S103P011P057nsss(0)='1'  )then
          oVar1S751(0) <='1';
          else
          oVar1S751(0) <='0';
          end if;
        if(cVar2S24S103P011N057P017nsss(0)='1'  OR cVar2S25S103N011P055P012nsss(0)='1'  OR cVar2S26S103P060P010P036nsss(0)='1'  OR cVar2S27S103P060N010P012nsss(0)='1'  )then
          oVar1S752(0) <='1';
          else
          oVar1S752(0) <='0';
          end if;
        if(cVar2S28S103P060P066nsss(0)='1'  OR cVar2S29S103P060N066P017nsss(0)='1'  OR cVar2S30S103P057P010P053nsss(0)='1'  OR cVar2S31S103P057P060nsss(0)='1'  )then
          oVar1S753(0) <='1';
          else
          oVar1S753(0) <='0';
          end if;
        if(cVar2S32S103P057N060P043nsss(0)='1'  )then
          oVar1S754(0) <='1';
          else
          oVar1S754(0) <='0';
          end if;
        if(cVar2S0S104P065nsss(0)='1'  OR cVar2S1S104P065P018nsss(0)='1'  OR cVar2S2S104P010nsss(0)='1'  OR cVar1S3S104P015P005P060P017nsss(0)='1'  )then
          oVar1S755(0) <='1';
          else
          oVar1S755(0) <='0';
          end if;
        if(cVar2S4S104P065nsss(0)='1'  OR cVar2S5S104P026P035P017nsss(0)='1'  OR cVar2S6S104P026N035P027nsss(0)='1'  OR cVar2S7S104P026P034nsss(0)='1'  )then
          oVar1S756(0) <='1';
          else
          oVar1S756(0) <='0';
          end if;
        if(cVar2S8S104P013P031nsss(0)='1'  OR cVar2S9S104P013N031P002nsss(0)='1'  OR cVar2S10S104N013P061P034nsss(0)='1'  OR cVar2S11S104P008P047nsss(0)='1'  )then
          oVar1S757(0) <='1';
          else
          oVar1S757(0) <='0';
          end if;
        if(cVar2S12S104P008N047P060nsss(0)='1'  OR cVar2S13S104N008P047P011nsss(0)='1'  OR cVar2S14S104N008P047P046nsss(0)='1'  OR cVar2S15S104P019nsss(0)='1'  )then
          oVar1S758(0) <='1';
          else
          oVar1S758(0) <='0';
          end if;
        if(cVar2S16S104P019P012nsss(0)='1'  OR cVar2S17S104P019N012P011nsss(0)='1'  OR cVar2S18S104P054P066nsss(0)='1'  OR cVar2S19S104N054P026nsss(0)='1'  )then
          oVar1S759(0) <='1';
          else
          oVar1S759(0) <='0';
          end if;
        if(cVar2S20S104N054P026P052nsss(0)='1'  OR cVar2S21S104P054P049P019nsss(0)='1'  OR cVar2S22S104P054N049P058nsss(0)='1'  OR cVar2S23S104P014nsss(0)='1'  )then
          oVar1S760(0) <='1';
          else
          oVar1S760(0) <='0';
          end if;
        if(cVar2S24S104P068nsss(0)='1'  OR cVar2S25S104N068P012P030nsss(0)='1'  OR cVar2S26S104N068N012P033nsss(0)='1'  )then
          oVar1S761(0) <='1';
          else
          oVar1S761(0) <='0';
          end if;
        if(cVar2S0S105P005P037nsss(0)='1'  OR cVar2S1S105N005psss(0)='1'  OR cVar2S2S105P008nsss(0)='1'  OR cVar2S3S105N008P011P010nsss(0)='1'  )then
          oVar1S762(0) <='1';
          else
          oVar1S762(0) <='0';
          end if;
        if(cVar2S4S105N008N011P010nsss(0)='1'  OR cVar1S5S105P017P015P018P060nsss(0)='1'  OR cVar2S6S105P061P035nsss(0)='1'  OR cVar2S7S105P061N035P059nsss(0)='1'  )then
          oVar1S763(0) <='1';
          else
          oVar1S763(0) <='0';
          end if;
        if(cVar2S8S105P029P050nsss(0)='1'  OR cVar2S9S105P029N050P054nsss(0)='1'  OR cVar2S10S105N029P024P011nsss(0)='1'  OR cVar2S11S105N029N024P028nsss(0)='1'  )then
          oVar1S764(0) <='1';
          else
          oVar1S764(0) <='0';
          end if;
        if(cVar2S12S105P025nsss(0)='1'  OR cVar2S13S105N025P050nsss(0)='1'  OR cVar2S14S105P013P033nsss(0)='1'  OR cVar2S15S105N013P012P068nsss(0)='1'  )then
          oVar1S765(0) <='1';
          else
          oVar1S765(0) <='0';
          end if;
        if(cVar2S16S105P066P059nsss(0)='1'  OR cVar2S17S105P066N059P035nsss(0)='1'  OR cVar2S18S105P066P037nsss(0)='1'  OR cVar2S19S105P016P036nsss(0)='1'  )then
          oVar1S766(0) <='1';
          else
          oVar1S766(0) <='0';
          end if;
        if(cVar2S20S105P016P036P067nsss(0)='1'  OR cVar2S21S105N016P035nsss(0)='1'  OR cVar2S22S105N016N035P013nsss(0)='1'  OR cVar2S23S105P062P039nsss(0)='1'  )then
          oVar1S767(0) <='1';
          else
          oVar1S767(0) <='0';
          end if;
        if(cVar2S24S105P062N039P061nsss(0)='1'  OR cVar2S25S105P062N064P052nsss(0)='1'  OR cVar2S26S105P067P063nsss(0)='1'  OR cVar2S27S105P067P063P069nsss(0)='1'  )then
          oVar1S768(0) <='1';
          else
          oVar1S768(0) <='0';
          end if;
        if(cVar2S28S105N067P036P010nsss(0)='1'  OR cVar1S29S105N017P015P005P004nsss(0)='1'  OR cVar2S30S105P012P069P008nsss(0)='1'  OR cVar2S31S105P012P014nsss(0)='1'  )then
          oVar1S769(0) <='1';
          else
          oVar1S769(0) <='0';
          end if;
        if(cVar2S32S105P014P048P012nsss(0)='1'  OR cVar2S33S105P014N048P060nsss(0)='1'  OR cVar2S34S105P014P009P062nsss(0)='1'  OR cVar2S35S105P016nsss(0)='1'  )then
          oVar1S770(0) <='1';
          else
          oVar1S770(0) <='0';
          end if;
        if(cVar2S36S105N016P006nsss(0)='1'  OR cVar2S37S105N016N006P004nsss(0)='1'  )then
          oVar1S771(0) <='1';
          else
          oVar1S771(0) <='0';
          end if;
        if(cVar2S0S106P069nsss(0)='1'  OR cVar2S1S106P062nsss(0)='1'  OR cVar2S2S106P052nsss(0)='1'  OR cVar2S3S106P052P008P028nsss(0)='1'  )then
          oVar1S772(0) <='1';
          else
          oVar1S772(0) <='0';
          end if;
        if(cVar2S4S106P052N008P009nsss(0)='1'  OR cVar2S5S106P022nsss(0)='1'  OR cVar2S6S106N022P049nsss(0)='1'  OR cVar2S7S106N022N049P003nsss(0)='1'  )then
          oVar1S773(0) <='1';
          else
          oVar1S773(0) <='0';
          end if;
        if(cVar2S8S106P036P007nsss(0)='1'  OR cVar2S9S106P055P012P019nsss(0)='1'  OR cVar2S10S106N055P021nsss(0)='1'  OR cVar2S11S106N055P021P018nsss(0)='1'  )then
          oVar1S774(0) <='1';
          else
          oVar1S774(0) <='0';
          end if;
        if(cVar2S12S106P021P016nsss(0)='1'  OR cVar2S13S106N021P018P056nsss(0)='1'  OR cVar2S14S106N021P018P032nsss(0)='1'  OR cVar1S15S106P065P052nsss(0)='1'  )then
          oVar1S775(0) <='1';
          else
          oVar1S775(0) <='0';
          end if;
        if(cVar2S16S106P037P036nsss(0)='1'  OR cVar2S17S106P037P036P016nsss(0)='1'  OR cVar2S18S106P037P019nsss(0)='1'  OR cVar2S19S106P015P067nsss(0)='1'  )then
          oVar1S776(0) <='1';
          else
          oVar1S776(0) <='0';
          end if;
        if(cVar2S20S106P015N067P034nsss(0)='1'  OR cVar2S21S106N015P062P034nsss(0)='1'  OR cVar2S22S106P059P024P053nsss(0)='1'  OR cVar2S23S106P059P068P016nsss(0)='1'  )then
          oVar1S777(0) <='1';
          else
          oVar1S777(0) <='0';
          end if;
        if(cVar2S24S106P036P037nsss(0)='1'  OR cVar2S25S106N036P067P063nsss(0)='1'  OR cVar2S26S106N036N067P037nsss(0)='1'  )then
          oVar1S778(0) <='1';
          else
          oVar1S778(0) <='0';
          end if;
        if(cVar1S0S107P052P065nsss(0)='1'  OR cVar2S1S107P069nsss(0)='1'  OR cVar2S2S107N069P064nsss(0)='1'  OR cVar2S3S107P015nsss(0)='1'  )then
          oVar1S779(0) <='1';
          else
          oVar1S779(0) <='0';
          end if;
        if(cVar2S4S107N015P011nsss(0)='1'  OR cVar2S5S107P009P029nsss(0)='1'  OR cVar2S6S107P009N029P027nsss(0)='1'  OR cVar2S7S107N009P008P048nsss(0)='1'  )then
          oVar1S780(0) <='1';
          else
          oVar1S780(0) <='0';
          end if;
        if(cVar2S8S107N009N008P011nsss(0)='1'  OR cVar1S9S107N052P044P025P005nsss(0)='1'  OR cVar2S10S107P006nsss(0)='1'  OR cVar2S11S107N006P007nsss(0)='1'  )then
          oVar1S781(0) <='1';
          else
          oVar1S781(0) <='0';
          end if;
        if(cVar1S12S107N052P044N025P067nsss(0)='1'  OR cVar2S13S107P054nsss(0)='1'  OR cVar2S14S107N054P023P005nsss(0)='1'  OR cVar2S15S107N054N023P062nsss(0)='1'  )then
          oVar1S782(0) <='1';
          else
          oVar1S782(0) <='0';
          end if;
        if(cVar2S16S107P006P047P014nsss(0)='1'  OR cVar2S17S107P006N047P043nsss(0)='1'  OR cVar2S18S107N006P060P035nsss(0)='1'  OR cVar2S19S107P006P035P037nsss(0)='1'  )then
          oVar1S783(0) <='1';
          else
          oVar1S783(0) <='0';
          end if;
        if(cVar2S20S107P013P010P014nsss(0)='1'  OR cVar2S21S107N013P012P015nsss(0)='1'  OR cVar2S22S107N013N012P014nsss(0)='1'  OR cVar2S23S107P056P012nsss(0)='1'  )then
          oVar1S784(0) <='1';
          else
          oVar1S784(0) <='0';
          end if;
        if(cVar2S24S107P056N012P010nsss(0)='1'  OR cVar2S25S107N056P014P037nsss(0)='1'  OR cVar2S26S107N056N014P010nsss(0)='1'  )then
          oVar1S785(0) <='1';
          else
          oVar1S785(0) <='0';
          end if;
        if(cVar2S0S108P024P014nsss(0)='1'  OR cVar2S1S108P024P014P017nsss(0)='1'  OR cVar2S2S108N024psss(0)='1'  OR cVar2S3S108P029P011P014nsss(0)='1'  )then
          oVar1S786(0) <='1';
          else
          oVar1S786(0) <='0';
          end if;
        if(cVar2S4S108P029N011P026nsss(0)='1'  OR cVar2S5S108N029psss(0)='1'  OR cVar2S6S108P063nsss(0)='1'  OR cVar2S7S108N063P010P017nsss(0)='1'  )then
          oVar1S787(0) <='1';
          else
          oVar1S787(0) <='0';
          end if;
        if(cVar2S8S108P062P064P035nsss(0)='1'  OR cVar2S9S108P062P064P034nsss(0)='1'  OR cVar2S10S108N062P019P015nsss(0)='1'  OR cVar2S11S108P069P066P003nsss(0)='1'  )then
          oVar1S788(0) <='1';
          else
          oVar1S788(0) <='0';
          end if;
        if(cVar2S12S108P069N066P062nsss(0)='1'  OR cVar2S13S108P069P034nsss(0)='1'  OR cVar2S14S108P019nsss(0)='1'  OR cVar2S15S108P010P012P069nsss(0)='1'  )then
          oVar1S789(0) <='1';
          else
          oVar1S789(0) <='0';
          end if;
        if(cVar2S16S108P010P012psss(0)='1'  OR cVar2S17S108P031P011nsss(0)='1'  OR cVar2S18S108N031P064nsss(0)='1'  OR cVar2S19S108N031N064P067nsss(0)='1'  )then
          oVar1S790(0) <='1';
          else
          oVar1S790(0) <='0';
          end if;
        if(cVar2S20S108P009P015P060nsss(0)='1'  OR cVar2S21S108P009P015P037nsss(0)='1'  OR cVar2S22S108P012P015P061nsss(0)='1'  OR cVar2S23S108P012P015P018nsss(0)='1'  )then
          oVar1S791(0) <='1';
          else
          oVar1S791(0) <='0';
          end if;
        if(cVar2S24S108N012P015P035nsss(0)='1'  OR cVar1S25S108P058P006P017nsss(0)='1'  )then
          oVar1S792(0) <='1';
          else
          oVar1S792(0) <='0';
          end if;
        if(cVar1S0S109P045P004P016P018nsss(0)='1'  OR cVar1S1S109P045N004P006P024nsss(0)='1'  OR cVar2S2S109P022nsss(0)='1'  OR cVar1S3S109P045N004N006P023nsss(0)='1'  )then
          oVar1S793(0) <='1';
          else
          oVar1S793(0) <='0';
          end if;
        if(cVar2S4S109P050nsss(0)='1'  OR cVar2S5S109N050P007nsss(0)='1'  OR cVar2S6S109N050N007P051nsss(0)='1'  OR cVar2S7S109P057P050P009nsss(0)='1'  )then
          oVar1S794(0) <='1';
          else
          oVar1S794(0) <='0';
          end if;
        if(cVar2S8S109P057P050P056nsss(0)='1'  OR cVar2S9S109P053nsss(0)='1'  OR cVar2S10S109N053P055nsss(0)='1'  OR cVar2S11S109N053N055P052nsss(0)='1'  )then
          oVar1S795(0) <='1';
          else
          oVar1S795(0) <='0';
          end if;
        if(cVar2S12S109P052nsss(0)='1'  OR cVar2S13S109N052P054nsss(0)='1'  OR cVar2S14S109P009P050nsss(0)='1'  OR cVar2S15S109P009N050P051nsss(0)='1'  )then
          oVar1S796(0) <='1';
          else
          oVar1S796(0) <='0';
          end if;
        if(cVar2S16S109N009P015P019nsss(0)='1'  OR cVar2S17S109P025P046nsss(0)='1'  OR cVar2S18S109P025N046P047nsss(0)='1'  OR cVar2S19S109N025P028P027nsss(0)='1'  )then
          oVar1S797(0) <='1';
          else
          oVar1S797(0) <='0';
          end if;
        if(cVar2S20S109P047P009P051nsss(0)='1'  OR cVar2S21S109P047P006P014nsss(0)='1'  OR cVar2S22S109P047N006P008nsss(0)='1'  OR cVar2S23S109P031P054nsss(0)='1'  )then
          oVar1S798(0) <='1';
          else
          oVar1S798(0) <='0';
          end if;
        if(cVar2S24S109P031N054P013nsss(0)='1'  OR cVar2S25S109N031P013P037nsss(0)='1'  OR cVar2S26S109N031N013P028nsss(0)='1'  OR cVar2S27S109P037P064nsss(0)='1'  )then
          oVar1S799(0) <='1';
          else
          oVar1S799(0) <='0';
          end if;
        if(cVar2S28S109N037P055nsss(0)='1'  )then
          oVar1S800(0) <='1';
          else
          oVar1S800(0) <='0';
          end if;
        if(cVar2S0S110P046nsss(0)='1'  OR cVar2S1S110N046P047nsss(0)='1'  OR cVar2S2S110N046N047P042nsss(0)='1'  OR cVar2S3S110P028P009P010nsss(0)='1'  )then
          oVar1S801(0) <='1';
          else
          oVar1S801(0) <='0';
          end if;
        if(cVar2S4S110P028N009psss(0)='1'  OR cVar2S5S110P009P027nsss(0)='1'  OR cVar2S6S110P009P027P008nsss(0)='1'  OR cVar2S7S110P009P050P027nsss(0)='1'  )then
          oVar1S802(0) <='1';
          else
          oVar1S802(0) <='0';
          end if;
        if(cVar2S8S110P009N050P013nsss(0)='1'  OR cVar2S9S110P006P024nsss(0)='1'  OR cVar2S10S110P006N024P026nsss(0)='1'  OR cVar2S11S110N006P009P050nsss(0)='1'  )then
          oVar1S803(0) <='1';
          else
          oVar1S803(0) <='0';
          end if;
        if(cVar2S12S110N006N009P008nsss(0)='1'  OR cVar2S13S110P052nsss(0)='1'  OR cVar2S14S110N052P054nsss(0)='1'  OR cVar2S15S110P009nsss(0)='1'  )then
          oVar1S804(0) <='1';
          else
          oVar1S804(0) <='0';
          end if;
        if(cVar2S16S110N009P013P054nsss(0)='1'  OR cVar2S17S110N009N013P015nsss(0)='1'  OR cVar2S18S110P050P012nsss(0)='1'  OR cVar2S19S110P050P056nsss(0)='1'  )then
          oVar1S805(0) <='1';
          else
          oVar1S805(0) <='0';
          end if;
        if(cVar1S20S110P011P029N054P053nsss(0)='1'  OR cVar2S21S110P055nsss(0)='1'  OR cVar2S22S110N055P052P014nsss(0)='1'  OR cVar2S23S110P047P026nsss(0)='1'  )then
          oVar1S806(0) <='1';
          else
          oVar1S806(0) <='0';
          end if;
        if(cVar2S24S110P047N026P015nsss(0)='1'  OR cVar2S25S110N047P020P018nsss(0)='1'  OR cVar2S26S110N047N020P010nsss(0)='1'  OR cVar2S27S110P056nsss(0)='1'  )then
          oVar1S807(0) <='1';
          else
          oVar1S807(0) <='0';
          end if;
        if(cVar2S28S110N056P057P012nsss(0)='1'  OR cVar2S29S110P012nsss(0)='1'  OR cVar2S30S110N012P009P036nsss(0)='1'  OR cVar2S31S110P018P035P015nsss(0)='1'  )then
          oVar1S808(0) <='1';
          else
          oVar1S808(0) <='0';
          end if;
        if(cVar2S32S110N018P014P009nsss(0)='1'  )then
          oVar1S809(0) <='1';
          else
          oVar1S809(0) <='0';
          end if;
        if(cVar1S0S111P009P049P025nsss(0)='1'  OR cVar2S1S111P068P019nsss(0)='1'  OR cVar1S2S111P009N049P053P029nsss(0)='1'  OR cVar2S3S111P003P063P068nsss(0)='1'  )then
          oVar1S810(0) <='1';
          else
          oVar1S810(0) <='0';
          end if;
        if(cVar2S4S111P027P013nsss(0)='1'  OR cVar2S5S111N027P029P011nsss(0)='1'  OR cVar2S6S111N027N029P016nsss(0)='1'  OR cVar2S7S111P007P036P010nsss(0)='1'  )then
          oVar1S811(0) <='1';
          else
          oVar1S811(0) <='0';
          end if;
        if(cVar2S8S111N007P027P013nsss(0)='1'  OR cVar1S9S111N009P044P004nsss(0)='1'  OR cVar1S10S111N009P044N004P051nsss(0)='1'  OR cVar2S11S111P021nsss(0)='1'  )then
          oVar1S812(0) <='1';
          else
          oVar1S812(0) <='0';
          end if;
        if(cVar2S12S111N021P011nsss(0)='1'  OR cVar2S13S111N021N011P007nsss(0)='1'  OR cVar2S14S111P068P069nsss(0)='1'  OR cVar2S15S111N068P031P013nsss(0)='1'  )then
          oVar1S813(0) <='1';
          else
          oVar1S813(0) <='0';
          end if;
        if(cVar2S16S111P004P043nsss(0)='1'  OR cVar2S17S111P004N043P064nsss(0)='1'  OR cVar1S18S111N009N044P042P058nsss(0)='1'  OR cVar2S19S111P023nsss(0)='1'  )then
          oVar1S814(0) <='1';
          else
          oVar1S814(0) <='0';
          end if;
        if(cVar2S20S111N023P021P002nsss(0)='1'  )then
          oVar1S815(0) <='1';
          else
          oVar1S815(0) <='0';
          end if;
        if(cVar1S0S112P009P049P025nsss(0)='1'  OR cVar2S1S112P068P013nsss(0)='1'  OR cVar2S2S112P011nsss(0)='1'  OR cVar2S3S112P029P016nsss(0)='1'  )then
          oVar1S816(0) <='1';
          else
          oVar1S816(0) <='0';
          end if;
        if(cVar2S4S112N029P066nsss(0)='1'  OR cVar2S5S112N029N066P015nsss(0)='1'  OR cVar2S6S112P029nsss(0)='1'  OR cVar2S7S112N029P035nsss(0)='1'  )then
          oVar1S817(0) <='1';
          else
          oVar1S817(0) <='0';
          end if;
        if(cVar2S8S112N029N035P015nsss(0)='1'  OR cVar2S9S112P051P010P068nsss(0)='1'  OR cVar2S10S112P051P010P065nsss(0)='1'  OR cVar2S11S112P034P060P059nsss(0)='1'  )then
          oVar1S818(0) <='1';
          else
          oVar1S818(0) <='0';
          end if;
        if(cVar2S12S112P034P060P068nsss(0)='1'  OR cVar2S13S112P034P014P016nsss(0)='1'  OR cVar2S14S112P037P059P058nsss(0)='1'  OR cVar2S15S112P037N059psss(0)='1'  )then
          oVar1S819(0) <='1';
          else
          oVar1S819(0) <='0';
          end if;
        if(cVar2S16S112P042nsss(0)='1'  OR cVar2S17S112N042P005nsss(0)='1'  OR cVar2S18S112N042N005P020nsss(0)='1'  OR cVar2S19S112P019P015nsss(0)='1'  )then
          oVar1S820(0) <='1';
          else
          oVar1S820(0) <='0';
          end if;
        if(cVar2S20S112P017nsss(0)='1'  OR cVar2S21S112N017P014P050nsss(0)='1'  OR cVar2S22S112P053nsss(0)='1'  OR cVar2S23S112N053P055nsss(0)='1'  )then
          oVar1S821(0) <='1';
          else
          oVar1S821(0) <='0';
          end if;
        if(cVar2S24S112N053N055P052nsss(0)='1'  OR cVar2S25S112P026nsss(0)='1'  OR cVar2S26S112N026P066nsss(0)='1'  OR cVar2S27S112N026N066P024nsss(0)='1'  )then
          oVar1S822(0) <='1';
          else
          oVar1S822(0) <='0';
          end if;
        if(cVar2S28S112P020P041nsss(0)='1'  OR cVar2S29S112P020N041P018nsss(0)='1'  OR cVar2S30S112N020P039P013nsss(0)='1'  )then
          oVar1S823(0) <='1';
          else
          oVar1S823(0) <='0';
          end if;
        if(cVar1S0S113P037P066P027P047nsss(0)='1'  OR cVar2S1S113P048P042P023nsss(0)='1'  OR cVar2S2S113P048P017P046nsss(0)='1'  OR cVar2S3S113P018nsss(0)='1'  )then
          oVar1S824(0) <='1';
          else
          oVar1S824(0) <='0';
          end if;
        if(cVar2S4S113P060P064P035nsss(0)='1'  OR cVar2S5S113P060P064P036nsss(0)='1'  OR cVar2S6S113P062nsss(0)='1'  OR cVar2S7S113P062P064P015nsss(0)='1'  )then
          oVar1S825(0) <='1';
          else
          oVar1S825(0) <='0';
          end if;
        if(cVar2S8S113P021nsss(0)='1'  OR cVar2S9S113N021P018P061nsss(0)='1'  OR cVar2S10S113N021N018P058nsss(0)='1'  OR cVar1S11S113N037P059P043nsss(0)='1'  )then
          oVar1S826(0) <='1';
          else
          oVar1S826(0) <='0';
          end if;
        if(cVar2S12S113P000P055P065nsss(0)='1'  OR cVar2S13S113P067nsss(0)='1'  OR cVar2S14S113N067P060P057nsss(0)='1'  OR cVar2S15S113P025nsss(0)='1'  )then
          oVar1S827(0) <='1';
          else
          oVar1S827(0) <='0';
          end if;
        if(cVar2S16S113N025P019nsss(0)='1'  OR cVar2S17S113N025P019P027nsss(0)='1'  OR cVar2S18S113P057P028nsss(0)='1'  OR cVar2S19S113P057N028P055nsss(0)='1'  )then
          oVar1S828(0) <='1';
          else
          oVar1S828(0) <='0';
          end if;
        if(cVar2S20S113N057P027P018nsss(0)='1'  OR cVar2S21S113N057N027P065nsss(0)='1'  OR cVar2S22S113P010P019nsss(0)='1'  OR cVar2S23S113P010P019P016nsss(0)='1'  )then
          oVar1S829(0) <='1';
          else
          oVar1S829(0) <='0';
          end if;
        if(cVar2S24S113N010P011P029nsss(0)='1'  OR cVar2S25S113N010N011P013nsss(0)='1'  OR cVar2S26S113P031P016P017nsss(0)='1'  OR cVar2S27S113P031N016P064nsss(0)='1'  )then
          oVar1S830(0) <='1';
          else
          oVar1S830(0) <='0';
          end if;
        if(cVar2S28S113P031P058P019nsss(0)='1'  )then
          oVar1S831(0) <='1';
          else
          oVar1S831(0) <='0';
          end if;
        if(cVar2S0S114P013nsss(0)='1'  OR cVar2S1S114P007P009nsss(0)='1'  OR cVar2S2S114N007P069P068nsss(0)='1'  OR cVar2S3S114N007P069P012nsss(0)='1'  )then
          oVar1S832(0) <='1';
          else
          oVar1S832(0) <='0';
          end if;
        if(cVar2S4S114P053P012nsss(0)='1'  OR cVar2S5S114P053P012P010nsss(0)='1'  OR cVar2S6S114N053P012P055nsss(0)='1'  OR cVar2S7S114N053N012P057nsss(0)='1'  )then
          oVar1S833(0) <='1';
          else
          oVar1S833(0) <='0';
          end if;
        if(cVar2S8S114P029P054P057nsss(0)='1'  OR cVar2S9S114P029N054P033nsss(0)='1'  OR cVar2S10S114N029P026P069nsss(0)='1'  OR cVar2S11S114N029N026P049nsss(0)='1'  )then
          oVar1S834(0) <='1';
          else
          oVar1S834(0) <='0';
          end if;
        if(cVar2S12S114P013P016nsss(0)='1'  OR cVar2S13S114P013P016P066nsss(0)='1'  OR cVar2S14S114N013P056nsss(0)='1'  OR cVar2S15S114N013N056P006nsss(0)='1'  )then
          oVar1S835(0) <='1';
          else
          oVar1S835(0) <='0';
          end if;
        if(cVar2S16S114P068P000P054nsss(0)='1'  OR cVar2S17S114N068P069P036nsss(0)='1'  OR cVar1S18S114P064P037P061P062nsss(0)='1'  OR cVar2S19S114P069nsss(0)='1'  )then
          oVar1S836(0) <='1';
          else
          oVar1S836(0) <='0';
          end if;
        if(cVar2S20S114N069P016P059nsss(0)='1'  OR cVar1S21S114P064P046nsss(0)='1'  OR cVar1S22S114P064N046P042nsss(0)='1'  OR cVar2S23S114P036P066nsss(0)='1'  )then
          oVar1S837(0) <='1';
          else
          oVar1S837(0) <='0';
          end if;
        if(cVar2S24S114N036P011P054nsss(0)='1'  OR cVar2S25S114P007P036P017nsss(0)='1'  OR cVar2S26S114P007N036P010nsss(0)='1'  )then
          oVar1S838(0) <='1';
          else
          oVar1S838(0) <='0';
          end if;
        if(cVar1S0S115P049P026P033P007nsss(0)='1'  OR cVar2S1S115P011nsss(0)='1'  OR cVar2S2S115N011P024nsss(0)='1'  OR cVar1S3S115P049N026P024P004nsss(0)='1'  )then
          oVar1S839(0) <='1';
          else
          oVar1S839(0) <='0';
          end if;
        if(cVar2S4S115P006P014nsss(0)='1'  OR cVar2S5S115N006P005nsss(0)='1'  OR cVar2S6S115N006N005P007nsss(0)='1'  OR cVar2S7S115P048nsss(0)='1'  )then
          oVar1S840(0) <='1';
          else
          oVar1S840(0) <='0';
          end if;
        if(cVar2S8S115P048P047nsss(0)='1'  OR cVar2S9S115P048P047P050nsss(0)='1'  OR cVar2S10S115P047P033nsss(0)='1'  OR cVar2S11S115P047N033P034nsss(0)='1'  )then
          oVar1S841(0) <='1';
          else
          oVar1S841(0) <='0';
          end if;
        if(cVar2S12S115P047P025nsss(0)='1'  OR cVar1S13S115N049P064P050P065nsss(0)='1'  OR cVar2S14S115P018nsss(0)='1'  OR cVar2S15S115N018P016P017nsss(0)='1'  )then
          oVar1S842(0) <='1';
          else
          oVar1S842(0) <='0';
          end if;
        if(cVar2S16S115P005P059nsss(0)='1'  OR cVar2S17S115P005P059P058nsss(0)='1'  OR cVar2S18S115P005P019P037nsss(0)='1'  OR cVar2S19S115P010P019P037nsss(0)='1'  )then
          oVar1S843(0) <='1';
          else
          oVar1S843(0) <='0';
          end if;
        if(cVar2S20S115P010N019P034nsss(0)='1'  OR cVar2S21S115P053P063nsss(0)='1'  OR cVar2S22S115N053P057nsss(0)='1'  OR cVar2S23S115N053N057P054nsss(0)='1'  )then
          oVar1S844(0) <='1';
          else
          oVar1S844(0) <='0';
          end if;
        if(cVar2S24S115P029P063nsss(0)='1'  OR cVar2S25S115N029P005P065nsss(0)='1'  OR cVar2S26S115N029N005P060nsss(0)='1'  OR cVar1S27S115N049N064P047P069nsss(0)='1'  )then
          oVar1S845(0) <='1';
          else
          oVar1S845(0) <='0';
          end if;
        if(cVar2S28S115P045P004nsss(0)='1'  OR cVar2S29S115P045N004P019nsss(0)='1'  OR cVar2S30S115N045P014P008nsss(0)='1'  )then
          oVar1S846(0) <='1';
          else
          oVar1S846(0) <='0';
          end if;
        if(cVar2S0S116P004nsss(0)='1'  OR cVar2S1S116N004P006P014nsss(0)='1'  OR cVar2S2S116N004N006psss(0)='1'  OR cVar2S3S116P026nsss(0)='1'  )then
          oVar1S847(0) <='1';
          else
          oVar1S847(0) <='0';
          end if;
        if(cVar2S4S116N026P027nsss(0)='1'  OR cVar2S5S116P064P042nsss(0)='1'  OR cVar2S6S116P064P042P002nsss(0)='1'  OR cVar2S7S116P064P066P034nsss(0)='1'  )then
          oVar1S848(0) <='1';
          else
          oVar1S848(0) <='0';
          end if;
        if(cVar2S8S116P045P004nsss(0)='1'  OR cVar2S9S116P045N004P015nsss(0)='1'  OR cVar2S10S116N045P069nsss(0)='1'  OR cVar1S11S116P060P062P050P014nsss(0)='1'  )then
          oVar1S849(0) <='1';
          else
          oVar1S849(0) <='0';
          end if;
        if(cVar2S12S116P007P025P003nsss(0)='1'  OR cVar2S13S116P007P065nsss(0)='1'  OR cVar2S14S116P057nsss(0)='1'  OR cVar2S15S116N057P026nsss(0)='1'  )then
          oVar1S850(0) <='1';
          else
          oVar1S850(0) <='0';
          end if;
        if(cVar2S16S116N057N026P034nsss(0)='1'  OR cVar1S17S116P060P014P008P032nsss(0)='1'  OR cVar2S18S116P015P012P067nsss(0)='1'  OR cVar2S19S116P015P064nsss(0)='1'  )then
          oVar1S851(0) <='1';
          else
          oVar1S851(0) <='0';
          end if;
        if(cVar2S20S116P019P067nsss(0)='1'  OR cVar2S21S116P019P018nsss(0)='1'  OR cVar2S22S116P019N018P017nsss(0)='1'  OR cVar2S23S116P015P067nsss(0)='1'  )then
          oVar1S852(0) <='1';
          else
          oVar1S852(0) <='0';
          end if;
        if(cVar2S24S116P015N067P061nsss(0)='1'  OR cVar2S25S116N015P012nsss(0)='1'  OR cVar2S26S116P016nsss(0)='1'  OR cVar2S27S116N016P058P015nsss(0)='1'  )then
          oVar1S853(0) <='1';
          else
          oVar1S853(0) <='0';
          end if;
        if(cVar2S28S116P031P010nsss(0)='1'  OR cVar2S29S116P031N010P013nsss(0)='1'  OR cVar2S30S116N031P035P064nsss(0)='1'  OR cVar2S31S116N031N035P047nsss(0)='1'  )then
          oVar1S854(0) <='1';
          else
          oVar1S854(0) <='0';
          end if;
        if(cVar1S0S117P049P005nsss(0)='1'  OR cVar1S1S117P049N005P026P033nsss(0)='1'  OR cVar2S2S117P004nsss(0)='1'  OR cVar2S3S117N004P006P008nsss(0)='1'  )then
          oVar1S856(0) <='1';
          else
          oVar1S856(0) <='0';
          end if;
        if(cVar2S4S117N004N006P007nsss(0)='1'  OR cVar2S5S117P027nsss(0)='1'  OR cVar2S6S117N027P047P033nsss(0)='1'  OR cVar2S7S117N027P047P025nsss(0)='1'  )then
          oVar1S857(0) <='1';
          else
          oVar1S857(0) <='0';
          end if;
        if(cVar2S8S117P014nsss(0)='1'  OR cVar2S9S117P014P016nsss(0)='1'  OR cVar2S10S117P026P066P011nsss(0)='1'  OR cVar2S11S117N026P029nsss(0)='1'  )then
          oVar1S858(0) <='1';
          else
          oVar1S858(0) <='0';
          end if;
        if(cVar2S12S117N026N029P048nsss(0)='1'  OR cVar2S13S117P025P048P067nsss(0)='1'  OR cVar2S14S117P025N048P043nsss(0)='1'  OR cVar2S15S117N025P046P052nsss(0)='1'  )then
          oVar1S859(0) <='1';
          else
          oVar1S859(0) <='0';
          end if;
        if(cVar2S16S117N025P046P030nsss(0)='1'  OR cVar2S17S117P052P017nsss(0)='1'  OR cVar2S18S117P052N017P061nsss(0)='1'  OR cVar1S19S117N049P024P026P002nsss(0)='1'  )then
          oVar1S860(0) <='1';
          else
          oVar1S860(0) <='0';
          end if;
        if(cVar2S20S117P068P006nsss(0)='1'  )then
          oVar1S861(0) <='1';
          else
          oVar1S861(0) <='0';
          end if;
        if(cVar1S0S118P049P006P024nsss(0)='1'  OR cVar1S1S118P049P006N024P026nsss(0)='1'  OR cVar2S2S118P036nsss(0)='1'  OR cVar2S3S118P017nsss(0)='1'  )then
          oVar1S862(0) <='1';
          else
          oVar1S862(0) <='0';
          end if;
        if(cVar2S4S118P025nsss(0)='1'  OR cVar2S5S118N025P068P017nsss(0)='1'  OR cVar2S6S118P005nsss(0)='1'  OR cVar2S7S118N005P008P010nsss(0)='1'  )then
          oVar1S863(0) <='1';
          else
          oVar1S863(0) <='0';
          end if;
        if(cVar2S8S118N005N008P047nsss(0)='1'  OR cVar2S9S118P058nsss(0)='1'  OR cVar2S10S118N058P039nsss(0)='1'  OR cVar2S11S118N058N039P023nsss(0)='1'  )then
          oVar1S864(0) <='1';
          else
          oVar1S864(0) <='0';
          end if;
        if(cVar2S12S118P005P004P043nsss(0)='1'  OR cVar2S13S118P005P014nsss(0)='1'  OR cVar2S14S118P005N014P038nsss(0)='1'  OR cVar2S15S118P057P004nsss(0)='1'  )then
          oVar1S865(0) <='1';
          else
          oVar1S865(0) <='0';
          end if;
        if(cVar2S16S118P057N004P006nsss(0)='1'  OR cVar2S17S118P016P011nsss(0)='1'  OR cVar1S18S118N049P052P065P066nsss(0)='1'  OR cVar2S19S118P015nsss(0)='1'  )then
          oVar1S866(0) <='1';
          else
          oVar1S866(0) <='0';
          end if;
        if(cVar2S20S118N015P011nsss(0)='1'  OR cVar2S21S118P010P003P014nsss(0)='1'  OR cVar2S22S118N010P009P019nsss(0)='1'  OR cVar2S23S118N010N009P008nsss(0)='1'  )then
          oVar1S867(0) <='1';
          else
          oVar1S867(0) <='0';
          end if;
        if(cVar1S0S119P049P006P007P018nsss(0)='1'  OR cVar2S1S119P017nsss(0)='1'  OR cVar1S2S119P049N006P007P025nsss(0)='1'  OR cVar2S3S119P019nsss(0)='1'  )then
          oVar1S869(0) <='1';
          else
          oVar1S869(0) <='0';
          end if;
        if(cVar2S4S119P025nsss(0)='1'  OR cVar2S5S119N025P051P047nsss(0)='1'  OR cVar2S6S119N025P051P047nsss(0)='1'  OR cVar2S7S119P005nsss(0)='1'  )then
          oVar1S870(0) <='1';
          else
          oVar1S870(0) <='0';
          end if;
        if(cVar2S8S119N005P008P026nsss(0)='1'  OR cVar1S9S119N049P042P051nsss(0)='1'  OR cVar2S10S119P004nsss(0)='1'  OR cVar2S11S119N004P039nsss(0)='1'  )then
          oVar1S871(0) <='1';
          else
          oVar1S871(0) <='0';
          end if;
        if(cVar2S12S119N004N039P005nsss(0)='1'  OR cVar1S13S119N049N042P045P022nsss(0)='1'  OR cVar2S14S119P048nsss(0)='1'  OR cVar2S15S119N048P063nsss(0)='1'  )then
          oVar1S872(0) <='1';
          else
          oVar1S872(0) <='0';
          end if;
        if(cVar2S16S119N048N063P061nsss(0)='1'  OR cVar2S17S119P023P020P003nsss(0)='1'  OR cVar2S18S119P023P056nsss(0)='1'  OR cVar2S19S119P023N056P041nsss(0)='1'  )then
          oVar1S873(0) <='1';
          else
          oVar1S873(0) <='0';
          end if;
        if(cVar2S20S119P069nsss(0)='1'  )then
          oVar1S874(0) <='1';
          else
          oVar1S874(0) <='0';
          end if;
        if(cVar2S0S120P018nsss(0)='1'  OR cVar2S1S120P018P019nsss(0)='1'  OR cVar2S2S120P016P018nsss(0)='1'  OR cVar1S3S120P049N024P026P007nsss(0)='1'  )then
          oVar1S875(0) <='1';
          else
          oVar1S875(0) <='0';
          end if;
        if(cVar2S4S120P008P019nsss(0)='1'  OR cVar2S5S120N008P011nsss(0)='1'  OR cVar2S6S120N008N011P006nsss(0)='1'  OR cVar1S7S120P049N024N026P027nsss(0)='1'  )then
          oVar1S876(0) <='1';
          else
          oVar1S876(0) <='0';
          end if;
        if(cVar2S8S120P047P034nsss(0)='1'  OR cVar2S9S120P047N034P033nsss(0)='1'  OR cVar2S10S120P047P025nsss(0)='1'  OR cVar2S11S120P023nsss(0)='1'  )then
          oVar1S877(0) <='1';
          else
          oVar1S877(0) <='0';
          end if;
        if(cVar2S12S120N023P040nsss(0)='1'  OR cVar2S13S120N023N040P022nsss(0)='1'  OR cVar2S14S120P002nsss(0)='1'  OR cVar2S15S120N002P058nsss(0)='1'  )then
          oVar1S878(0) <='1';
          else
          oVar1S878(0) <='0';
          end if;
        if(cVar2S16S120N002N058P025nsss(0)='1'  OR cVar1S17S120N049N042P045P022nsss(0)='1'  OR cVar2S18S120P023P017nsss(0)='1'  OR cVar2S19S120N023P003P024nsss(0)='1'  )then
          oVar1S879(0) <='1';
          else
          oVar1S879(0) <='0';
          end if;
        if(cVar2S20S120P023nsss(0)='1'  OR cVar2S21S120P023P056nsss(0)='1'  OR cVar2S22S120P023N056P041nsss(0)='1'  OR cVar2S23S120P026P067nsss(0)='1'  )then
          oVar1S880(0) <='1';
          else
          oVar1S880(0) <='0';
          end if;
        if(cVar1S0S121P049P024P010P006nsss(0)='1'  OR cVar2S1S121P016P018nsss(0)='1'  OR cVar1S2S121P049N024P026P007nsss(0)='1'  OR cVar2S3S121P008P019nsss(0)='1'  )then
          oVar1S882(0) <='1';
          else
          oVar1S882(0) <='0';
          end if;
        if(cVar2S4S121N008P011nsss(0)='1'  OR cVar2S5S121N008N011P006nsss(0)='1'  OR cVar1S6S121P049N024N026P027nsss(0)='1'  OR cVar2S7S121P047P017nsss(0)='1'  )then
          oVar1S883(0) <='1';
          else
          oVar1S883(0) <='0';
          end if;
        if(cVar2S8S121P047N017P014nsss(0)='1'  OR cVar2S9S121P047P025nsss(0)='1'  OR cVar1S10S121N049P042P051nsss(0)='1'  OR cVar1S11S121N049P042N051P050nsss(0)='1'  )then
          oVar1S884(0) <='1';
          else
          oVar1S884(0) <='0';
          end if;
        if(cVar2S12S121P013P022nsss(0)='1'  OR cVar2S13S121P014P013nsss(0)='1'  OR cVar2S14S121N014P051nsss(0)='1'  OR cVar2S15S121N014N051P060nsss(0)='1'  )then
          oVar1S885(0) <='1';
          else
          oVar1S885(0) <='0';
          end if;
        if(cVar2S16S121P012P056P030nsss(0)='1'  OR cVar2S17S121N012P041nsss(0)='1'  OR cVar2S18S121P026P067nsss(0)='1'  )then
          oVar1S886(0) <='1';
          else
          oVar1S886(0) <='0';
          end if;
        if(cVar1S0S122P045P027P024P013nsss(0)='1'  OR cVar2S1S122P006nsss(0)='1'  OR cVar2S2S122N006P004nsss(0)='1'  OR cVar2S3S122N006N004P047nsss(0)='1'  )then
          oVar1S887(0) <='1';
          else
          oVar1S887(0) <='0';
          end if;
        if(cVar2S4S122P043nsss(0)='1'  OR cVar2S5S122N043P046nsss(0)='1'  OR cVar2S6S122P022nsss(0)='1'  OR cVar2S7S122N022P023P017nsss(0)='1'  )then
          oVar1S888(0) <='1';
          else
          oVar1S888(0) <='0';
          end if;
        if(cVar2S8S122N022N023P043nsss(0)='1'  OR cVar2S9S122P004nsss(0)='1'  OR cVar2S10S122N004P017nsss(0)='1'  OR cVar2S11S122N004P017P018nsss(0)='1'  )then
          oVar1S889(0) <='1';
          else
          oVar1S889(0) <='0';
          end if;
        if(cVar2S12S122P007nsss(0)='1'  OR cVar2S13S122N007P008P019nsss(0)='1'  OR cVar2S14S122N007N008P011nsss(0)='1'  OR cVar2S15S122P027nsss(0)='1'  )then
          oVar1S890(0) <='1';
          else
          oVar1S890(0) <='0';
          end if;
        if(cVar2S16S122N027P047nsss(0)='1'  OR cVar2S17S122N027P047P025nsss(0)='1'  OR cVar2S18S122P051nsss(0)='1'  OR cVar2S19S122N051P004nsss(0)='1'  )then
          oVar1S891(0) <='1';
          else
          oVar1S891(0) <='0';
          end if;
        if(cVar2S20S122N051N004P002nsss(0)='1'  OR cVar2S21S122P012P056nsss(0)='1'  OR cVar2S22S122P012N056P043nsss(0)='1'  OR cVar2S23S122N012P032P007nsss(0)='1'  )then
          oVar1S892(0) <='1';
          else
          oVar1S892(0) <='0';
          end if;
        if(cVar2S24S122N012P032P057nsss(0)='1'  OR cVar1S25S122N045N049P047P064nsss(0)='1'  OR cVar2S26S122P069nsss(0)='1'  OR cVar2S27S122N069P014P008nsss(0)='1'  )then
          oVar1S893(0) <='1';
          else
          oVar1S893(0) <='0';
          end if;
        if(cVar1S0S123P042P051nsss(0)='1'  OR cVar1S1S123P042N051P050P039nsss(0)='1'  OR cVar2S2S123P004nsss(0)='1'  OR cVar2S3S123N004P025nsss(0)='1'  )then
          oVar1S895(0) <='1';
          else
          oVar1S895(0) <='0';
          end if;
        if(cVar2S4S123N004N025P058nsss(0)='1'  OR cVar1S5S123N042P049P024P004nsss(0)='1'  OR cVar2S6S123P006P008nsss(0)='1'  OR cVar2S7S123N006P005nsss(0)='1'  )then
          oVar1S896(0) <='1';
          else
          oVar1S896(0) <='0';
          end if;
        if(cVar2S8S123N006N005P026nsss(0)='1'  OR cVar2S9S123P007nsss(0)='1'  OR cVar2S10S123N007P011nsss(0)='1'  OR cVar2S11S123N007N011P008nsss(0)='1'  )then
          oVar1S897(0) <='1';
          else
          oVar1S897(0) <='0';
          end if;
        if(cVar2S12S123P027nsss(0)='1'  OR cVar2S13S123N027P047P017nsss(0)='1'  OR cVar2S14S123N027P047P025nsss(0)='1'  OR cVar2S15S123P022nsss(0)='1'  )then
          oVar1S898(0) <='1';
          else
          oVar1S898(0) <='0';
          end if;
        if(cVar2S16S123N022P015nsss(0)='1'  OR cVar2S17S123P004P013P022nsss(0)='1'  OR cVar2S18S123N004P006nsss(0)='1'  OR cVar2S19S123N004N006P057nsss(0)='1'  )then
          oVar1S899(0) <='1';
          else
          oVar1S899(0) <='0';
          end if;
        if(cVar2S20S123P009P050P027nsss(0)='1'  OR cVar2S21S123P009N050P008nsss(0)='1'  OR cVar2S22S123P026P014P012nsss(0)='1'  )then
          oVar1S900(0) <='1';
          else
          oVar1S900(0) <='0';
          end if;
        if(cVar1S0S124P042P050P021nsss(0)='1'  OR cVar1S1S124P042P050N021P051nsss(0)='1'  OR cVar2S2S124P025nsss(0)='1'  OR cVar2S3S124N025P058nsss(0)='1'  )then
          oVar1S901(0) <='1';
          else
          oVar1S901(0) <='0';
          end if;
        if(cVar2S4S124N025N058P039nsss(0)='1'  OR cVar2S5S124P006nsss(0)='1'  OR cVar2S6S124N006P004nsss(0)='1'  OR cVar2S7S124N006N004P007nsss(0)='1'  )then
          oVar1S902(0) <='1';
          else
          oVar1S902(0) <='0';
          end if;
        if(cVar2S8S124P025P043nsss(0)='1'  OR cVar2S9S124P025N043P046nsss(0)='1'  OR cVar2S10S124N025P001nsss(0)='1'  OR cVar2S11S124N025N001P022nsss(0)='1'  )then
          oVar1S903(0) <='1';
          else
          oVar1S903(0) <='0';
          end if;
        if(cVar2S12S124P004nsss(0)='1'  OR cVar2S13S124N004P006P008nsss(0)='1'  OR cVar2S14S124N004N006P026nsss(0)='1'  OR cVar2S15S124P026nsss(0)='1'  )then
          oVar1S904(0) <='1';
          else
          oVar1S904(0) <='0';
          end if;
        if(cVar2S16S124N026P027nsss(0)='1'  OR cVar2S17S124N026N027P047nsss(0)='1'  OR cVar2S18S124P019P046nsss(0)='1'  OR cVar2S19S124P019P046P064nsss(0)='1'  )then
          oVar1S905(0) <='1';
          else
          oVar1S905(0) <='0';
          end if;
        if(cVar2S20S124N019P016P021nsss(0)='1'  OR cVar2S21S124N019N016psss(0)='1'  OR cVar2S22S124P026P014P066nsss(0)='1'  )then
          oVar1S906(0) <='1';
          else
          oVar1S906(0) <='0';
          end if;
        if(cVar1S0S125P042P050nsss(0)='1'  OR cVar2S1S125P006nsss(0)='1'  OR cVar2S2S125N006P004nsss(0)='1'  OR cVar2S3S125N006N004P007nsss(0)='1'  )then
          oVar1S907(0) <='1';
          else
          oVar1S907(0) <='0';
          end if;
        if(cVar1S4S125N042P045P027N024psss(0)='1'  OR cVar2S5S125P004nsss(0)='1'  OR cVar2S6S125N004P006P008nsss(0)='1'  OR cVar2S7S125N004N006P005nsss(0)='1'  )then
          oVar1S908(0) <='1';
          else
          oVar1S908(0) <='0';
          end if;
        if(cVar2S8S125P026nsss(0)='1'  OR cVar2S9S125N026P027nsss(0)='1'  OR cVar2S10S125P030P057nsss(0)='1'  OR cVar2S11S125P030N057P056nsss(0)='1'  )then
          oVar1S909(0) <='1';
          else
          oVar1S909(0) <='0';
          end if;
        if(cVar2S12S125P059P038P021nsss(0)='1'  OR cVar2S13S125P059N038P028nsss(0)='1'  )then
          oVar1S910(0) <='1';
          else
          oVar1S910(0) <='0';
          end if;
        if(cVar1S0S126P042P051nsss(0)='1'  OR cVar1S1S126P042N051P023P005nsss(0)='1'  OR cVar2S2S126P004nsss(0)='1'  OR cVar2S3S126N004P007nsss(0)='1'  )then
          oVar1S911(0) <='1';
          else
          oVar1S911(0) <='0';
          end if;
        if(cVar2S4S126N004N007P006nsss(0)='1'  OR cVar1S5S126P042N051N023P000nsss(0)='1'  OR cVar2S6S126P050P039nsss(0)='1'  OR cVar2S7S126P050N039P021nsss(0)='1'  )then
          oVar1S912(0) <='1';
          else
          oVar1S912(0) <='0';
          end if;
        if(cVar2S8S126P006nsss(0)='1'  OR cVar2S9S126N006P004nsss(0)='1'  OR cVar2S10S126N006N004P047nsss(0)='1'  OR cVar2S11S126P025P043nsss(0)='1'  )then
          oVar1S913(0) <='1';
          else
          oVar1S913(0) <='0';
          end if;
        if(cVar2S12S126P025N043P046nsss(0)='1'  OR cVar2S13S126N025P036nsss(0)='1'  OR cVar2S14S126N025N036P061nsss(0)='1'  OR cVar2S15S126P006P019nsss(0)='1'  )then
          oVar1S914(0) <='1';
          else
          oVar1S914(0) <='0';
          end if;
        if(cVar2S16S126P009P051nsss(0)='1'  OR cVar2S17S126P009P051P047nsss(0)='1'  OR cVar2S18S126N009P006P014nsss(0)='1'  OR cVar2S19S126N009N006P005nsss(0)='1'  )then
          oVar1S915(0) <='1';
          else
          oVar1S915(0) <='0';
          end if;
        if(cVar2S20S126P043nsss(0)='1'  OR cVar2S21S126P043P003nsss(0)='1'  OR cVar2S22S126P043N003P067nsss(0)='1'  OR cVar2S23S126P043nsss(0)='1'  )then
          oVar1S916(0) <='1';
          else
          oVar1S916(0) <='0';
          end if;
        if(cVar2S24S126N043P067nsss(0)='1'  )then
          oVar1S917(0) <='1';
          else
          oVar1S917(0) <='0';
          end if;
        if(cVar1S0S127P042P050P004P040nsss(0)='1'  OR cVar2S1S127P044nsss(0)='1'  OR cVar1S2S127P042P050N004P005nsss(0)='1'  OR cVar2S3S127P053nsss(0)='1'  )then
          oVar1S918(0) <='1';
          else
          oVar1S918(0) <='0';
          end if;
        if(cVar2S4S127N053P002nsss(0)='1'  OR cVar2S5S127N053N002P058nsss(0)='1'  OR cVar1S6S127N042P049P024P004nsss(0)='1'  OR cVar2S7S127P006P014nsss(0)='1'  )then
          oVar1S919(0) <='1';
          else
          oVar1S919(0) <='0';
          end if;
        if(cVar2S8S127N006P005nsss(0)='1'  OR cVar2S9S127N006N005P026nsss(0)='1'  OR cVar2S10S127P007nsss(0)='1'  OR cVar2S11S127N007P011nsss(0)='1'  )then
          oVar1S920(0) <='1';
          else
          oVar1S920(0) <='0';
          end if;
        if(cVar2S12S127N007N011P008nsss(0)='1'  OR cVar2S13S127P027nsss(0)='1'  OR cVar2S14S127N027P047P043nsss(0)='1'  OR cVar2S15S127N027P047P025nsss(0)='1'  )then
          oVar1S921(0) <='1';
          else
          oVar1S921(0) <='0';
          end if;
        if(cVar2S16S127P006nsss(0)='1'  OR cVar2S17S127N006P004nsss(0)='1'  OR cVar2S18S127N006N004P007nsss(0)='1'  OR cVar2S19S127P025P043nsss(0)='1'  )then
          oVar1S922(0) <='1';
          else
          oVar1S922(0) <='0';
          end if;
        if(cVar2S20S127P025N043P046nsss(0)='1'  OR cVar2S21S127N025P011nsss(0)='1'  OR cVar2S22S127N025N011P013nsss(0)='1'  OR cVar2S23S127P003nsss(0)='1'  )then
          oVar1S923(0) <='1';
          else
          oVar1S923(0) <='0';
          end if;
        if(cVar2S24S127N003P048nsss(0)='1'  OR cVar2S25S127N003N048P002nsss(0)='1'  OR cVar2S26S127P039P047P034nsss(0)='1'  OR cVar2S27S127P039P021nsss(0)='1'  )then
          oVar1S924(0) <='1';
          else
          oVar1S924(0) <='0';
          end if;
        if(cVar2S28S127P039N021P016nsss(0)='1'  )then
          oVar1S925(0) <='1';
          else
          oVar1S925(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV4 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar1S0(0)='1'  OR oVar1S1(0)='1'  OR oVar1S2(0)='1'  OR oVar1S3(0)='1'  )then
          oVar2S0(0) <='1';
          else
          oVar2S0(0) <='0';
          end if;
        if(oVar1S4(0)='1'  OR oVar1S5(0)='1'  )then
          oVar2S1(0) <='1';
          else
          oVar2S1(0) <='0';
          end if;
        if(oVar1S7(0)='1'  OR oVar1S8(0)='1'  OR oVar1S9(0)='1'  OR oVar1S10(0)='1'  )then
          oVar2S2(0) <='1';
          else
          oVar2S2(0) <='0';
          end if;
        if(oVar1S11(0)='1'  OR oVar1S12(0)='1'  OR oVar1S13(0)='1'  )then
          oVar2S3(0) <='1';
          else
          oVar2S3(0) <='0';
          end if;
        if(oVar1S14(0)='1'  OR oVar1S15(0)='1'  OR oVar1S16(0)='1'  OR oVar1S17(0)='1'  )then
          oVar2S4(0) <='1';
          else
          oVar2S4(0) <='0';
          end if;
        if(oVar1S18(0)='1'  OR oVar1S19(0)='1'  OR oVar1S20(0)='1'  )then
          oVar2S5(0) <='1';
          else
          oVar2S5(0) <='0';
          end if;
        if(oVar1S21(0)='1'  OR oVar1S22(0)='1'  OR oVar1S23(0)='1'  OR oVar1S24(0)='1'  )then
          oVar2S6(0) <='1';
          else
          oVar2S6(0) <='0';
          end if;
        if(oVar1S25(0)='1'  OR oVar1S26(0)='1'  OR oVar1S27(0)='1'  OR oVar1S28(0)='1'  )then
          oVar2S7(0) <='1';
          else
          oVar2S7(0) <='0';
          end if;
        if(oVar1S29(0)='1'  OR oVar1S30(0)='1'  OR oVar1S31(0)='1'  OR oVar1S32(0)='1'  )then
          oVar2S9(0) <='1';
          else
          oVar2S9(0) <='0';
          end if;
        if(oVar1S33(0)='1'  )then
          oVar2S10(0) <='1';
          else
          oVar2S10(0) <='0';
          end if;
        if(oVar1S34(0)='1'  OR oVar1S35(0)='1'  OR oVar1S36(0)='1'  OR oVar1S37(0)='1'  )then
          oVar2S11(0) <='1';
          else
          oVar2S11(0) <='0';
          end if;
        if(oVar1S38(0)='1'  OR oVar1S39(0)='1'  )then
          oVar2S12(0) <='1';
          else
          oVar2S12(0) <='0';
          end if;
        if(oVar1S40(0)='1'  OR oVar1S41(0)='1'  OR oVar1S42(0)='1'  OR oVar1S43(0)='1'  )then
          oVar2S13(0) <='1';
          else
          oVar2S13(0) <='0';
          end if;
        if(oVar1S44(0)='1'  OR oVar1S45(0)='1'  OR oVar1S46(0)='1'  )then
          oVar2S14(0) <='1';
          else
          oVar2S14(0) <='0';
          end if;
        if(oVar1S47(0)='1'  OR oVar1S48(0)='1'  OR oVar1S49(0)='1'  OR oVar1S50(0)='1'  )then
          oVar2S15(0) <='1';
          else
          oVar2S15(0) <='0';
          end if;
        if(oVar1S51(0)='1'  OR oVar1S52(0)='1'  OR oVar1S53(0)='1'  )then
          oVar2S16(0) <='1';
          else
          oVar2S16(0) <='0';
          end if;
        if(oVar1S54(0)='1'  OR oVar1S55(0)='1'  OR oVar1S56(0)='1'  OR oVar1S57(0)='1'  )then
          oVar2S17(0) <='1';
          else
          oVar2S17(0) <='0';
          end if;
        if(oVar1S58(0)='1'  OR oVar1S59(0)='1'  OR oVar1S60(0)='1'  OR oVar1S61(0)='1'  )then
          oVar2S18(0) <='1';
          else
          oVar2S18(0) <='0';
          end if;
        if(oVar1S62(0)='1'  OR oVar1S63(0)='1'  OR oVar1S64(0)='1'  OR oVar1S65(0)='1'  )then
          oVar2S20(0) <='1';
          else
          oVar2S20(0) <='0';
          end if;
        if(oVar1S66(0)='1'  OR oVar1S67(0)='1'  )then
          oVar2S21(0) <='1';
          else
          oVar2S21(0) <='0';
          end if;
        if(oVar1S68(0)='1'  OR oVar1S69(0)='1'  OR oVar1S70(0)='1'  OR oVar1S71(0)='1'  )then
          oVar2S22(0) <='1';
          else
          oVar2S22(0) <='0';
          end if;
        if(oVar1S72(0)='1'  OR oVar1S73(0)='1'  OR oVar1S74(0)='1'  OR oVar1S75(0)='1'  )then
          oVar2S23(0) <='1';
          else
          oVar2S23(0) <='0';
          end if;
        if(oVar1S76(0)='1'  )then
          oVar2S24(0) <='1';
          else
          oVar2S24(0) <='0';
          end if;
        if(oVar1S77(0)='1'  OR oVar1S78(0)='1'  OR oVar1S79(0)='1'  OR oVar1S80(0)='1'  )then
          oVar2S25(0) <='1';
          else
          oVar2S25(0) <='0';
          end if;
        if(oVar1S81(0)='1'  OR oVar1S82(0)='1'  OR oVar1S83(0)='1'  OR oVar1S84(0)='1'  )then
          oVar2S26(0) <='1';
          else
          oVar2S26(0) <='0';
          end if;
        if(oVar1S85(0)='1'  OR oVar1S86(0)='1'  OR oVar1S87(0)='1'  OR oVar1S88(0)='1'  )then
          oVar2S28(0) <='1';
          else
          oVar2S28(0) <='0';
          end if;
        if(oVar1S89(0)='1'  OR oVar1S90(0)='1'  )then
          oVar2S29(0) <='1';
          else
          oVar2S29(0) <='0';
          end if;
        if(oVar1S91(0)='1'  OR oVar1S92(0)='1'  OR oVar1S93(0)='1'  OR oVar1S94(0)='1'  )then
          oVar2S30(0) <='1';
          else
          oVar2S30(0) <='0';
          end if;
        if(oVar1S95(0)='1'  OR oVar1S96(0)='1'  OR oVar1S97(0)='1'  )then
          oVar2S31(0) <='1';
          else
          oVar2S31(0) <='0';
          end if;
        if(oVar1S99(0)='1'  OR oVar1S100(0)='1'  OR oVar1S101(0)='1'  OR oVar1S102(0)='1'  )then
          oVar2S33(0) <='1';
          else
          oVar2S33(0) <='0';
          end if;
        if(oVar1S103(0)='1'  OR oVar1S104(0)='1'  OR oVar1S105(0)='1'  OR oVar1S106(0)='1'  )then
          oVar2S34(0) <='1';
          else
          oVar2S34(0) <='0';
          end if;
        if(oVar1S107(0)='1'  OR oVar1S108(0)='1'  OR oVar1S109(0)='1'  OR oVar1S110(0)='1'  )then
          oVar2S36(0) <='1';
          else
          oVar2S36(0) <='0';
          end if;
        if(oVar1S111(0)='1'  OR oVar1S112(0)='1'  OR oVar1S113(0)='1'  OR oVar1S114(0)='1'  )then
          oVar2S37(0) <='1';
          else
          oVar2S37(0) <='0';
          end if;
        if(oVar1S115(0)='1'  OR oVar1S116(0)='1'  OR oVar1S117(0)='1'  OR oVar1S118(0)='1'  )then
          oVar2S39(0) <='1';
          else
          oVar2S39(0) <='0';
          end if;
        if(oVar1S119(0)='1'  OR oVar1S120(0)='1'  OR oVar1S121(0)='1'  OR oVar1S122(0)='1'  )then
          oVar2S40(0) <='1';
          else
          oVar2S40(0) <='0';
          end if;
        if(oVar1S123(0)='1'  OR oVar1S124(0)='1'  OR oVar1S125(0)='1'  OR oVar1S126(0)='1'  )then
          oVar2S42(0) <='1';
          else
          oVar2S42(0) <='0';
          end if;
        if(oVar1S127(0)='1'  OR oVar1S128(0)='1'  OR oVar1S129(0)='1'  )then
          oVar2S43(0) <='1';
          else
          oVar2S43(0) <='0';
          end if;
        if(oVar1S130(0)='1'  OR oVar1S131(0)='1'  OR oVar1S132(0)='1'  OR oVar1S133(0)='1'  )then
          oVar2S44(0) <='1';
          else
          oVar2S44(0) <='0';
          end if;
        if(oVar1S134(0)='1'  )then
          oVar2S45(0) <='1';
          else
          oVar2S45(0) <='0';
          end if;
        if(oVar1S135(0)='1'  OR oVar1S136(0)='1'  OR oVar1S137(0)='1'  OR oVar1S138(0)='1'  )then
          oVar2S46(0) <='1';
          else
          oVar2S46(0) <='0';
          end if;
        if(oVar1S139(0)='1'  OR oVar1S140(0)='1'  )then
          oVar2S47(0) <='1';
          else
          oVar2S47(0) <='0';
          end if;
        if(oVar1S141(0)='1'  OR oVar1S142(0)='1'  OR oVar1S143(0)='1'  OR oVar1S144(0)='1'  )then
          oVar2S48(0) <='1';
          else
          oVar2S48(0) <='0';
          end if;
        if(oVar1S145(0)='1'  OR oVar1S146(0)='1'  OR oVar1S147(0)='1'  OR oVar1S148(0)='1'  )then
          oVar2S49(0) <='1';
          else
          oVar2S49(0) <='0';
          end if;
        if(oVar1S149(0)='1'  OR oVar1S150(0)='1'  OR oVar1S151(0)='1'  OR oVar1S152(0)='1'  )then
          oVar2S51(0) <='1';
          else
          oVar2S51(0) <='0';
          end if;
        if(oVar1S153(0)='1'  )then
          oVar2S52(0) <='1';
          else
          oVar2S52(0) <='0';
          end if;
        if(oVar1S154(0)='1'  OR oVar1S155(0)='1'  OR oVar1S156(0)='1'  OR oVar1S157(0)='1'  )then
          oVar2S53(0) <='1';
          else
          oVar2S53(0) <='0';
          end if;
        if(oVar1S158(0)='1'  )then
          oVar2S54(0) <='1';
          else
          oVar2S54(0) <='0';
          end if;
        if(oVar1S160(0)='1'  OR oVar1S161(0)='1'  OR oVar1S162(0)='1'  OR oVar1S163(0)='1'  )then
          oVar2S55(0) <='1';
          else
          oVar2S55(0) <='0';
          end if;
        if(oVar1S164(0)='1'  )then
          oVar2S56(0) <='1';
          else
          oVar2S56(0) <='0';
          end if;
        if(oVar1S166(0)='1'  OR oVar1S167(0)='1'  OR oVar1S168(0)='1'  OR oVar1S169(0)='1'  )then
          oVar2S57(0) <='1';
          else
          oVar2S57(0) <='0';
          end if;
        if(oVar1S170(0)='1'  OR oVar1S171(0)='1'  )then
          oVar2S58(0) <='1';
          else
          oVar2S58(0) <='0';
          end if;
        if(oVar1S172(0)='1'  OR oVar1S173(0)='1'  OR oVar1S174(0)='1'  OR oVar1S175(0)='1'  )then
          oVar2S59(0) <='1';
          else
          oVar2S59(0) <='0';
          end if;
        if(oVar1S176(0)='1'  OR oVar1S177(0)='1'  )then
          oVar2S60(0) <='1';
          else
          oVar2S60(0) <='0';
          end if;
        if(oVar1S178(0)='1'  OR oVar1S179(0)='1'  OR oVar1S180(0)='1'  OR oVar1S181(0)='1'  )then
          oVar2S61(0) <='1';
          else
          oVar2S61(0) <='0';
          end if;
        if(oVar1S182(0)='1'  OR oVar1S183(0)='1'  OR oVar1S184(0)='1'  OR oVar1S185(0)='1'  )then
          oVar2S62(0) <='1';
          else
          oVar2S62(0) <='0';
          end if;
        if(oVar1S187(0)='1'  OR oVar1S188(0)='1'  OR oVar1S189(0)='1'  OR oVar1S190(0)='1'  )then
          oVar2S64(0) <='1';
          else
          oVar2S64(0) <='0';
          end if;
        if(oVar1S191(0)='1'  OR oVar1S192(0)='1'  OR oVar1S193(0)='1'  OR oVar1S194(0)='1'  )then
          oVar2S65(0) <='1';
          else
          oVar2S65(0) <='0';
          end if;
        if(oVar1S195(0)='1'  OR oVar1S196(0)='1'  OR oVar1S197(0)='1'  OR oVar1S198(0)='1'  )then
          oVar2S67(0) <='1';
          else
          oVar2S67(0) <='0';
          end if;
        if(oVar1S199(0)='1'  OR oVar1S200(0)='1'  )then
          oVar2S68(0) <='1';
          else
          oVar2S68(0) <='0';
          end if;
        if(oVar1S201(0)='1'  OR oVar1S202(0)='1'  OR oVar1S203(0)='1'  OR oVar1S204(0)='1'  )then
          oVar2S69(0) <='1';
          else
          oVar2S69(0) <='0';
          end if;
        if(oVar1S205(0)='1'  OR oVar1S206(0)='1'  )then
          oVar2S70(0) <='1';
          else
          oVar2S70(0) <='0';
          end if;
        if(oVar1S208(0)='1'  OR oVar1S209(0)='1'  OR oVar1S210(0)='1'  OR oVar1S211(0)='1'  )then
          oVar2S71(0) <='1';
          else
          oVar2S71(0) <='0';
          end if;
        if(oVar1S212(0)='1'  OR oVar1S213(0)='1'  OR oVar1S214(0)='1'  OR oVar1S215(0)='1'  )then
          oVar2S72(0) <='1';
          else
          oVar2S72(0) <='0';
          end if;
        if(oVar1S216(0)='1'  )then
          oVar2S73(0) <='1';
          else
          oVar2S73(0) <='0';
          end if;
        if(oVar1S217(0)='1'  OR oVar1S218(0)='1'  OR oVar1S219(0)='1'  OR oVar1S220(0)='1'  )then
          oVar2S74(0) <='1';
          else
          oVar2S74(0) <='0';
          end if;
        if(oVar1S221(0)='1'  OR oVar1S222(0)='1'  OR oVar1S223(0)='1'  )then
          oVar2S75(0) <='1';
          else
          oVar2S75(0) <='0';
          end if;
        if(oVar1S224(0)='1'  OR oVar1S225(0)='1'  OR oVar1S226(0)='1'  OR oVar1S227(0)='1'  )then
          oVar2S76(0) <='1';
          else
          oVar2S76(0) <='0';
          end if;
        if(oVar1S228(0)='1'  OR oVar1S229(0)='1'  OR oVar1S230(0)='1'  OR oVar1S231(0)='1'  )then
          oVar2S77(0) <='1';
          else
          oVar2S77(0) <='0';
          end if;
        if(oVar1S232(0)='1'  OR oVar1S233(0)='1'  )then
          oVar2S78(0) <='1';
          else
          oVar2S78(0) <='0';
          end if;
        if(oVar1S234(0)='1'  OR oVar1S235(0)='1'  OR oVar1S236(0)='1'  OR oVar1S237(0)='1'  )then
          oVar2S79(0) <='1';
          else
          oVar2S79(0) <='0';
          end if;
        if(oVar1S238(0)='1'  OR oVar1S239(0)='1'  OR oVar1S240(0)='1'  OR oVar1S241(0)='1'  )then
          oVar2S80(0) <='1';
          else
          oVar2S80(0) <='0';
          end if;
        if(oVar1S243(0)='1'  OR oVar1S244(0)='1'  OR oVar1S245(0)='1'  OR oVar1S246(0)='1'  )then
          oVar2S82(0) <='1';
          else
          oVar2S82(0) <='0';
          end if;
        if(oVar1S247(0)='1'  OR oVar1S248(0)='1'  OR oVar1S249(0)='1'  OR oVar1S250(0)='1'  )then
          oVar2S83(0) <='1';
          else
          oVar2S83(0) <='0';
          end if;
        if(oVar1S251(0)='1'  OR oVar1S252(0)='1'  OR oVar1S253(0)='1'  OR oVar1S254(0)='1'  )then
          oVar2S85(0) <='1';
          else
          oVar2S85(0) <='0';
          end if;
        if(oVar1S255(0)='1'  OR oVar1S256(0)='1'  OR oVar1S257(0)='1'  )then
          oVar2S86(0) <='1';
          else
          oVar2S86(0) <='0';
          end if;
        if(oVar1S258(0)='1'  OR oVar1S259(0)='1'  OR oVar1S260(0)='1'  OR oVar1S261(0)='1'  )then
          oVar2S87(0) <='1';
          else
          oVar2S87(0) <='0';
          end if;
        if(oVar1S262(0)='1'  OR oVar1S263(0)='1'  OR oVar1S264(0)='1'  )then
          oVar2S88(0) <='1';
          else
          oVar2S88(0) <='0';
          end if;
        if(oVar1S265(0)='1'  OR oVar1S266(0)='1'  OR oVar1S267(0)='1'  OR oVar1S268(0)='1'  )then
          oVar2S89(0) <='1';
          else
          oVar2S89(0) <='0';
          end if;
        if(oVar1S269(0)='1'  OR oVar1S270(0)='1'  OR oVar1S271(0)='1'  )then
          oVar2S90(0) <='1';
          else
          oVar2S90(0) <='0';
          end if;
        if(oVar1S272(0)='1'  OR oVar1S273(0)='1'  OR oVar1S274(0)='1'  OR oVar1S275(0)='1'  )then
          oVar2S91(0) <='1';
          else
          oVar2S91(0) <='0';
          end if;
        if(oVar1S276(0)='1'  OR oVar1S277(0)='1'  OR oVar1S278(0)='1'  )then
          oVar2S92(0) <='1';
          else
          oVar2S92(0) <='0';
          end if;
        if(oVar1S280(0)='1'  OR oVar1S281(0)='1'  OR oVar1S282(0)='1'  OR oVar1S283(0)='1'  )then
          oVar2S94(0) <='1';
          else
          oVar2S94(0) <='0';
          end if;
        if(oVar1S284(0)='1'  OR oVar1S285(0)='1'  OR oVar1S286(0)='1'  OR oVar1S287(0)='1'  )then
          oVar2S95(0) <='1';
          else
          oVar2S95(0) <='0';
          end if;
        if(oVar1S288(0)='1'  OR oVar1S289(0)='1'  OR oVar1S290(0)='1'  OR oVar1S291(0)='1'  )then
          oVar2S97(0) <='1';
          else
          oVar2S97(0) <='0';
          end if;
        if(oVar1S292(0)='1'  OR oVar1S293(0)='1'  OR oVar1S294(0)='1'  OR oVar1S295(0)='1'  )then
          oVar2S98(0) <='1';
          else
          oVar2S98(0) <='0';
          end if;
        if(oVar1S296(0)='1'  OR oVar1S297(0)='1'  OR oVar1S298(0)='1'  OR oVar1S299(0)='1'  )then
          oVar2S100(0) <='1';
          else
          oVar2S100(0) <='0';
          end if;
        if(oVar1S300(0)='1'  OR oVar1S301(0)='1'  OR oVar1S302(0)='1'  OR oVar1S303(0)='1'  )then
          oVar2S101(0) <='1';
          else
          oVar2S101(0) <='0';
          end if;
        if(oVar1S304(0)='1'  OR oVar1S305(0)='1'  OR oVar1S306(0)='1'  OR oVar1S307(0)='1'  )then
          oVar2S103(0) <='1';
          else
          oVar2S103(0) <='0';
          end if;
        if(oVar1S308(0)='1'  OR oVar1S309(0)='1'  OR oVar1S310(0)='1'  )then
          oVar2S104(0) <='1';
          else
          oVar2S104(0) <='0';
          end if;
        if(oVar1S312(0)='1'  OR oVar1S313(0)='1'  OR oVar1S314(0)='1'  OR oVar1S315(0)='1'  )then
          oVar2S106(0) <='1';
          else
          oVar2S106(0) <='0';
          end if;
        if(oVar1S316(0)='1'  OR oVar1S317(0)='1'  OR oVar1S318(0)='1'  )then
          oVar2S107(0) <='1';
          else
          oVar2S107(0) <='0';
          end if;
        if(oVar1S319(0)='1'  OR oVar1S320(0)='1'  OR oVar1S321(0)='1'  OR oVar1S322(0)='1'  )then
          oVar2S108(0) <='1';
          else
          oVar2S108(0) <='0';
          end if;
        if(oVar1S323(0)='1'  OR oVar1S324(0)='1'  )then
          oVar2S109(0) <='1';
          else
          oVar2S109(0) <='0';
          end if;
        if(oVar1S325(0)='1'  OR oVar1S326(0)='1'  OR oVar1S327(0)='1'  OR oVar1S328(0)='1'  )then
          oVar2S110(0) <='1';
          else
          oVar2S110(0) <='0';
          end if;
        if(oVar1S329(0)='1'  OR oVar1S330(0)='1'  OR oVar1S331(0)='1'  )then
          oVar2S111(0) <='1';
          else
          oVar2S111(0) <='0';
          end if;
        if(oVar1S332(0)='1'  OR oVar1S333(0)='1'  OR oVar1S334(0)='1'  OR oVar1S335(0)='1'  )then
          oVar2S112(0) <='1';
          else
          oVar2S112(0) <='0';
          end if;
        if(oVar1S336(0)='1'  OR oVar1S337(0)='1'  )then
          oVar2S113(0) <='1';
          else
          oVar2S113(0) <='0';
          end if;
        if(oVar1S338(0)='1'  OR oVar1S339(0)='1'  OR oVar1S340(0)='1'  OR oVar1S341(0)='1'  )then
          oVar2S114(0) <='1';
          else
          oVar2S114(0) <='0';
          end if;
        if(oVar1S342(0)='1'  OR oVar1S343(0)='1'  )then
          oVar2S115(0) <='1';
          else
          oVar2S115(0) <='0';
          end if;
        if(oVar1S345(0)='1'  OR oVar1S346(0)='1'  OR oVar1S347(0)='1'  OR oVar1S348(0)='1'  )then
          oVar2S116(0) <='1';
          else
          oVar2S116(0) <='0';
          end if;
        if(oVar1S349(0)='1'  OR oVar1S350(0)='1'  OR oVar1S351(0)='1'  OR oVar1S352(0)='1'  )then
          oVar2S117(0) <='1';
          else
          oVar2S117(0) <='0';
          end if;
        if(oVar1S354(0)='1'  OR oVar1S355(0)='1'  OR oVar1S356(0)='1'  OR oVar1S357(0)='1'  )then
          oVar2S119(0) <='1';
          else
          oVar2S119(0) <='0';
          end if;
        if(oVar1S358(0)='1'  OR oVar1S359(0)='1'  OR oVar1S360(0)='1'  )then
          oVar2S120(0) <='1';
          else
          oVar2S120(0) <='0';
          end if;
        if(oVar1S361(0)='1'  OR oVar1S362(0)='1'  OR oVar1S363(0)='1'  OR oVar1S364(0)='1'  )then
          oVar2S121(0) <='1';
          else
          oVar2S121(0) <='0';
          end if;
        if(oVar1S365(0)='1'  )then
          oVar2S122(0) <='1';
          else
          oVar2S122(0) <='0';
          end if;
        if(oVar1S367(0)='1'  OR oVar1S368(0)='1'  OR oVar1S369(0)='1'  OR oVar1S370(0)='1'  )then
          oVar2S123(0) <='1';
          else
          oVar2S123(0) <='0';
          end if;
        if(oVar1S371(0)='1'  )then
          oVar2S124(0) <='1';
          else
          oVar2S124(0) <='0';
          end if;
        if(oVar1S372(0)='1'  OR oVar1S373(0)='1'  OR oVar1S374(0)='1'  OR oVar1S375(0)='1'  )then
          oVar2S125(0) <='1';
          else
          oVar2S125(0) <='0';
          end if;
        if(oVar1S376(0)='1'  OR oVar1S377(0)='1'  OR oVar1S378(0)='1'  OR oVar1S379(0)='1'  )then
          oVar2S126(0) <='1';
          else
          oVar2S126(0) <='0';
          end if;
        if(oVar1S380(0)='1'  OR oVar1S381(0)='1'  OR oVar1S382(0)='1'  OR oVar1S383(0)='1'  )then
          oVar2S128(0) <='1';
          else
          oVar2S128(0) <='0';
          end if;
        if(oVar1S384(0)='1'  OR oVar1S385(0)='1'  )then
          oVar2S129(0) <='1';
          else
          oVar2S129(0) <='0';
          end if;
        if(oVar1S387(0)='1'  OR oVar1S388(0)='1'  OR oVar1S389(0)='1'  OR oVar1S390(0)='1'  )then
          oVar2S130(0) <='1';
          else
          oVar2S130(0) <='0';
          end if;
        if(oVar1S391(0)='1'  OR oVar1S392(0)='1'  OR oVar1S393(0)='1'  )then
          oVar2S131(0) <='1';
          else
          oVar2S131(0) <='0';
          end if;
        if(oVar1S394(0)='1'  OR oVar1S395(0)='1'  OR oVar1S396(0)='1'  OR oVar1S397(0)='1'  )then
          oVar2S132(0) <='1';
          else
          oVar2S132(0) <='0';
          end if;
        if(oVar1S398(0)='1'  OR oVar1S399(0)='1'  OR oVar1S400(0)='1'  )then
          oVar2S133(0) <='1';
          else
          oVar2S133(0) <='0';
          end if;
        if(oVar1S401(0)='1'  OR oVar1S402(0)='1'  OR oVar1S403(0)='1'  OR oVar1S404(0)='1'  )then
          oVar2S134(0) <='1';
          else
          oVar2S134(0) <='0';
          end if;
        if(oVar1S405(0)='1'  OR oVar1S406(0)='1'  )then
          oVar2S135(0) <='1';
          else
          oVar2S135(0) <='0';
          end if;
        if(oVar1S407(0)='1'  OR oVar1S408(0)='1'  OR oVar1S409(0)='1'  OR oVar1S410(0)='1'  )then
          oVar2S136(0) <='1';
          else
          oVar2S136(0) <='0';
          end if;
        if(oVar1S411(0)='1'  OR oVar1S412(0)='1'  OR oVar1S413(0)='1'  )then
          oVar2S137(0) <='1';
          else
          oVar2S137(0) <='0';
          end if;
        if(oVar1S414(0)='1'  OR oVar1S415(0)='1'  OR oVar1S416(0)='1'  OR oVar1S417(0)='1'  )then
          oVar2S138(0) <='1';
          else
          oVar2S138(0) <='0';
          end if;
        if(oVar1S418(0)='1'  OR oVar1S419(0)='1'  OR oVar1S420(0)='1'  )then
          oVar2S139(0) <='1';
          else
          oVar2S139(0) <='0';
          end if;
        if(oVar1S421(0)='1'  OR oVar1S422(0)='1'  OR oVar1S423(0)='1'  OR oVar1S424(0)='1'  )then
          oVar2S140(0) <='1';
          else
          oVar2S140(0) <='0';
          end if;
        if(oVar1S425(0)='1'  OR oVar1S426(0)='1'  )then
          oVar2S141(0) <='1';
          else
          oVar2S141(0) <='0';
          end if;
        if(oVar1S427(0)='1'  OR oVar1S428(0)='1'  OR oVar1S429(0)='1'  OR oVar1S430(0)='1'  )then
          oVar2S142(0) <='1';
          else
          oVar2S142(0) <='0';
          end if;
        if(oVar1S431(0)='1'  OR oVar1S432(0)='1'  OR oVar1S433(0)='1'  )then
          oVar2S143(0) <='1';
          else
          oVar2S143(0) <='0';
          end if;
        if(oVar1S434(0)='1'  OR oVar1S435(0)='1'  OR oVar1S436(0)='1'  OR oVar1S437(0)='1'  )then
          oVar2S144(0) <='1';
          else
          oVar2S144(0) <='0';
          end if;
        if(oVar1S438(0)='1'  OR oVar1S439(0)='1'  )then
          oVar2S145(0) <='1';
          else
          oVar2S145(0) <='0';
          end if;
        if(oVar1S440(0)='1'  OR oVar1S441(0)='1'  OR oVar1S442(0)='1'  OR oVar1S443(0)='1'  )then
          oVar2S146(0) <='1';
          else
          oVar2S146(0) <='0';
          end if;
        if(oVar1S444(0)='1'  OR oVar1S445(0)='1'  OR oVar1S446(0)='1'  )then
          oVar2S147(0) <='1';
          else
          oVar2S147(0) <='0';
          end if;
        if(oVar1S447(0)='1'  OR oVar1S448(0)='1'  OR oVar1S449(0)='1'  OR oVar1S450(0)='1'  )then
          oVar2S148(0) <='1';
          else
          oVar2S148(0) <='0';
          end if;
        if(oVar1S451(0)='1'  OR oVar1S452(0)='1'  OR oVar1S453(0)='1'  )then
          oVar2S149(0) <='1';
          else
          oVar2S149(0) <='0';
          end if;
        if(oVar1S454(0)='1'  OR oVar1S455(0)='1'  OR oVar1S456(0)='1'  OR oVar1S457(0)='1'  )then
          oVar2S150(0) <='1';
          else
          oVar2S150(0) <='0';
          end if;
        if(oVar1S458(0)='1'  OR oVar1S459(0)='1'  OR oVar1S460(0)='1'  OR oVar1S461(0)='1'  )then
          oVar2S151(0) <='1';
          else
          oVar2S151(0) <='0';
          end if;
        if(oVar1S462(0)='1'  )then
          oVar2S152(0) <='1';
          else
          oVar2S152(0) <='0';
          end if;
        if(oVar1S463(0)='1'  OR oVar1S464(0)='1'  OR oVar1S465(0)='1'  OR oVar1S466(0)='1'  )then
          oVar2S153(0) <='1';
          else
          oVar2S153(0) <='0';
          end if;
        if(oVar1S467(0)='1'  OR oVar1S468(0)='1'  OR oVar1S469(0)='1'  )then
          oVar2S154(0) <='1';
          else
          oVar2S154(0) <='0';
          end if;
        if(oVar1S470(0)='1'  OR oVar1S471(0)='1'  OR oVar1S472(0)='1'  OR oVar1S473(0)='1'  )then
          oVar2S155(0) <='1';
          else
          oVar2S155(0) <='0';
          end if;
        if(oVar1S474(0)='1'  OR oVar1S475(0)='1'  OR oVar1S476(0)='1'  )then
          oVar2S156(0) <='1';
          else
          oVar2S156(0) <='0';
          end if;
        if(oVar1S477(0)='1'  OR oVar1S478(0)='1'  OR oVar1S479(0)='1'  OR oVar1S480(0)='1'  )then
          oVar2S157(0) <='1';
          else
          oVar2S157(0) <='0';
          end if;
        if(oVar1S481(0)='1'  OR oVar1S482(0)='1'  OR oVar1S483(0)='1'  )then
          oVar2S158(0) <='1';
          else
          oVar2S158(0) <='0';
          end if;
        if(oVar1S484(0)='1'  OR oVar1S485(0)='1'  OR oVar1S486(0)='1'  OR oVar1S487(0)='1'  )then
          oVar2S159(0) <='1';
          else
          oVar2S159(0) <='0';
          end if;
        if(oVar1S488(0)='1'  OR oVar1S489(0)='1'  OR oVar1S490(0)='1'  OR oVar1S491(0)='1'  )then
          oVar2S160(0) <='1';
          else
          oVar2S160(0) <='0';
          end if;
        if(oVar1S493(0)='1'  OR oVar1S494(0)='1'  OR oVar1S495(0)='1'  OR oVar1S496(0)='1'  )then
          oVar2S162(0) <='1';
          else
          oVar2S162(0) <='0';
          end if;
        if(oVar1S497(0)='1'  OR oVar1S498(0)='1'  OR oVar1S499(0)='1'  OR oVar1S500(0)='1'  )then
          oVar2S163(0) <='1';
          else
          oVar2S163(0) <='0';
          end if;
        if(oVar1S502(0)='1'  OR oVar1S503(0)='1'  OR oVar1S504(0)='1'  OR oVar1S505(0)='1'  )then
          oVar2S165(0) <='1';
          else
          oVar2S165(0) <='0';
          end if;
        if(oVar1S506(0)='1'  OR oVar1S507(0)='1'  OR oVar1S508(0)='1'  )then
          oVar2S166(0) <='1';
          else
          oVar2S166(0) <='0';
          end if;
        if(oVar1S510(0)='1'  OR oVar1S511(0)='1'  OR oVar1S512(0)='1'  OR oVar1S513(0)='1'  )then
          oVar2S168(0) <='1';
          else
          oVar2S168(0) <='0';
          end if;
        if(oVar1S514(0)='1'  OR oVar1S515(0)='1'  OR oVar1S516(0)='1'  )then
          oVar2S169(0) <='1';
          else
          oVar2S169(0) <='0';
          end if;
        if(oVar1S517(0)='1'  OR oVar1S518(0)='1'  OR oVar1S519(0)='1'  OR oVar1S520(0)='1'  )then
          oVar2S170(0) <='1';
          else
          oVar2S170(0) <='0';
          end if;
        if(oVar1S521(0)='1'  OR oVar1S522(0)='1'  OR oVar1S523(0)='1'  OR oVar1S524(0)='1'  )then
          oVar2S171(0) <='1';
          else
          oVar2S171(0) <='0';
          end if;
        if(oVar1S525(0)='1'  OR oVar1S526(0)='1'  OR oVar1S527(0)='1'  OR oVar1S528(0)='1'  )then
          oVar2S173(0) <='1';
          else
          oVar2S173(0) <='0';
          end if;
        if(oVar1S529(0)='1'  OR oVar1S530(0)='1'  OR oVar1S531(0)='1'  OR oVar1S532(0)='1'  )then
          oVar2S174(0) <='1';
          else
          oVar2S174(0) <='0';
          end if;
        if(oVar1S533(0)='1'  OR oVar1S534(0)='1'  OR oVar1S535(0)='1'  OR oVar1S536(0)='1'  )then
          oVar2S176(0) <='1';
          else
          oVar2S176(0) <='0';
          end if;
        if(oVar1S537(0)='1'  OR oVar1S538(0)='1'  OR oVar1S539(0)='1'  OR oVar1S540(0)='1'  )then
          oVar2S177(0) <='1';
          else
          oVar2S177(0) <='0';
          end if;
        if(oVar1S541(0)='1'  OR oVar1S542(0)='1'  OR oVar1S543(0)='1'  OR oVar1S544(0)='1'  )then
          oVar2S179(0) <='1';
          else
          oVar2S179(0) <='0';
          end if;
        if(oVar1S545(0)='1'  OR oVar1S546(0)='1'  OR oVar1S547(0)='1'  )then
          oVar2S180(0) <='1';
          else
          oVar2S180(0) <='0';
          end if;
        if(oVar1S549(0)='1'  OR oVar1S550(0)='1'  OR oVar1S551(0)='1'  OR oVar1S552(0)='1'  )then
          oVar2S182(0) <='1';
          else
          oVar2S182(0) <='0';
          end if;
        if(oVar1S553(0)='1'  OR oVar1S554(0)='1'  OR oVar1S555(0)='1'  )then
          oVar2S183(0) <='1';
          else
          oVar2S183(0) <='0';
          end if;
        if(oVar1S556(0)='1'  OR oVar1S557(0)='1'  OR oVar1S558(0)='1'  OR oVar1S559(0)='1'  )then
          oVar2S184(0) <='1';
          else
          oVar2S184(0) <='0';
          end if;
        if(oVar1S560(0)='1'  OR oVar1S561(0)='1'  OR oVar1S562(0)='1'  OR oVar1S563(0)='1'  )then
          oVar2S185(0) <='1';
          else
          oVar2S185(0) <='0';
          end if;
        if(oVar1S564(0)='1'  OR oVar1S565(0)='1'  OR oVar1S566(0)='1'  OR oVar1S567(0)='1'  )then
          oVar2S187(0) <='1';
          else
          oVar2S187(0) <='0';
          end if;
        if(oVar1S568(0)='1'  OR oVar1S569(0)='1'  OR oVar1S570(0)='1'  OR oVar1S571(0)='1'  )then
          oVar2S188(0) <='1';
          else
          oVar2S188(0) <='0';
          end if;
        if(oVar1S572(0)='1'  OR oVar1S573(0)='1'  OR oVar1S574(0)='1'  OR oVar1S575(0)='1'  )then
          oVar2S190(0) <='1';
          else
          oVar2S190(0) <='0';
          end if;
        if(oVar1S576(0)='1'  OR oVar1S577(0)='1'  OR oVar1S578(0)='1'  OR oVar1S579(0)='1'  )then
          oVar2S191(0) <='1';
          else
          oVar2S191(0) <='0';
          end if;
        if(oVar1S580(0)='1'  OR oVar1S581(0)='1'  OR oVar1S582(0)='1'  OR oVar1S583(0)='1'  )then
          oVar2S193(0) <='1';
          else
          oVar2S193(0) <='0';
          end if;
        if(oVar1S584(0)='1'  OR oVar1S585(0)='1'  OR oVar1S586(0)='1'  )then
          oVar2S194(0) <='1';
          else
          oVar2S194(0) <='0';
          end if;
        if(oVar1S587(0)='1'  OR oVar1S588(0)='1'  OR oVar1S589(0)='1'  OR oVar1S590(0)='1'  )then
          oVar2S195(0) <='1';
          else
          oVar2S195(0) <='0';
          end if;
        if(oVar1S591(0)='1'  OR oVar1S592(0)='1'  )then
          oVar2S196(0) <='1';
          else
          oVar2S196(0) <='0';
          end if;
        if(oVar1S593(0)='1'  OR oVar1S594(0)='1'  OR oVar1S595(0)='1'  OR oVar1S596(0)='1'  )then
          oVar2S197(0) <='1';
          else
          oVar2S197(0) <='0';
          end if;
        if(oVar1S597(0)='1'  OR oVar1S598(0)='1'  OR oVar1S599(0)='1'  )then
          oVar2S198(0) <='1';
          else
          oVar2S198(0) <='0';
          end if;
        if(oVar1S600(0)='1'  OR oVar1S601(0)='1'  OR oVar1S602(0)='1'  OR oVar1S603(0)='1'  )then
          oVar2S199(0) <='1';
          else
          oVar2S199(0) <='0';
          end if;
        if(oVar1S604(0)='1'  OR oVar1S605(0)='1'  )then
          oVar2S200(0) <='1';
          else
          oVar2S200(0) <='0';
          end if;
        if(oVar1S607(0)='1'  OR oVar1S608(0)='1'  OR oVar1S609(0)='1'  OR oVar1S610(0)='1'  )then
          oVar2S201(0) <='1';
          else
          oVar2S201(0) <='0';
          end if;
        if(oVar1S611(0)='1'  OR oVar1S612(0)='1'  OR oVar1S613(0)='1'  OR oVar1S614(0)='1'  )then
          oVar2S202(0) <='1';
          else
          oVar2S202(0) <='0';
          end if;
        if(oVar1S615(0)='1'  OR oVar1S616(0)='1'  OR oVar1S617(0)='1'  OR oVar1S618(0)='1'  )then
          oVar2S204(0) <='1';
          else
          oVar2S204(0) <='0';
          end if;
        if(oVar1S619(0)='1'  OR oVar1S620(0)='1'  )then
          oVar2S205(0) <='1';
          else
          oVar2S205(0) <='0';
          end if;
        if(oVar1S622(0)='1'  OR oVar1S623(0)='1'  OR oVar1S624(0)='1'  OR oVar1S625(0)='1'  )then
          oVar2S206(0) <='1';
          else
          oVar2S206(0) <='0';
          end if;
        if(oVar1S626(0)='1'  OR oVar1S627(0)='1'  OR oVar1S628(0)='1'  )then
          oVar2S207(0) <='1';
          else
          oVar2S207(0) <='0';
          end if;
        if(oVar1S629(0)='1'  OR oVar1S630(0)='1'  OR oVar1S631(0)='1'  OR oVar1S632(0)='1'  )then
          oVar2S208(0) <='1';
          else
          oVar2S208(0) <='0';
          end if;
        if(oVar1S633(0)='1'  OR oVar1S634(0)='1'  OR oVar1S635(0)='1'  )then
          oVar2S209(0) <='1';
          else
          oVar2S209(0) <='0';
          end if;
        if(oVar1S637(0)='1'  OR oVar1S638(0)='1'  OR oVar1S639(0)='1'  OR oVar1S640(0)='1'  )then
          oVar2S211(0) <='1';
          else
          oVar2S211(0) <='0';
          end if;
        if(oVar1S641(0)='1'  OR oVar1S642(0)='1'  OR oVar1S643(0)='1'  )then
          oVar2S212(0) <='1';
          else
          oVar2S212(0) <='0';
          end if;
        if(oVar1S644(0)='1'  OR oVar1S645(0)='1'  OR oVar1S646(0)='1'  OR oVar1S647(0)='1'  )then
          oVar2S213(0) <='1';
          else
          oVar2S213(0) <='0';
          end if;
        if(oVar1S648(0)='1'  OR oVar1S649(0)='1'  OR oVar1S650(0)='1'  OR oVar1S651(0)='1'  )then
          oVar2S214(0) <='1';
          else
          oVar2S214(0) <='0';
          end if;
        if(oVar1S652(0)='1'  OR oVar1S653(0)='1'  OR oVar1S654(0)='1'  OR oVar1S655(0)='1'  )then
          oVar2S216(0) <='1';
          else
          oVar2S216(0) <='0';
          end if;
        if(oVar1S656(0)='1'  )then
          oVar2S217(0) <='1';
          else
          oVar2S217(0) <='0';
          end if;
        if(oVar1S657(0)='1'  OR oVar1S658(0)='1'  OR oVar1S659(0)='1'  OR oVar1S660(0)='1'  )then
          oVar2S218(0) <='1';
          else
          oVar2S218(0) <='0';
          end if;
        if(oVar1S661(0)='1'  OR oVar1S662(0)='1'  )then
          oVar2S219(0) <='1';
          else
          oVar2S219(0) <='0';
          end if;
        if(oVar1S663(0)='1'  OR oVar1S664(0)='1'  OR oVar1S665(0)='1'  OR oVar1S666(0)='1'  )then
          oVar2S220(0) <='1';
          else
          oVar2S220(0) <='0';
          end if;
        if(oVar1S667(0)='1'  OR oVar1S668(0)='1'  )then
          oVar2S221(0) <='1';
          else
          oVar2S221(0) <='0';
          end if;
        if(oVar1S669(0)='1'  OR oVar1S670(0)='1'  OR oVar1S671(0)='1'  OR oVar1S672(0)='1'  )then
          oVar2S222(0) <='1';
          else
          oVar2S222(0) <='0';
          end if;
        if(oVar1S673(0)='1'  OR oVar1S674(0)='1'  OR oVar1S675(0)='1'  OR oVar1S676(0)='1'  )then
          oVar2S223(0) <='1';
          else
          oVar2S223(0) <='0';
          end if;
        if(oVar1S677(0)='1'  OR oVar1S678(0)='1'  OR oVar1S679(0)='1'  OR oVar1S680(0)='1'  )then
          oVar2S225(0) <='1';
          else
          oVar2S225(0) <='0';
          end if;
        if(oVar1S681(0)='1'  OR oVar1S682(0)='1'  )then
          oVar2S226(0) <='1';
          else
          oVar2S226(0) <='0';
          end if;
        if(oVar1S684(0)='1'  OR oVar1S685(0)='1'  OR oVar1S686(0)='1'  OR oVar1S687(0)='1'  )then
          oVar2S227(0) <='1';
          else
          oVar2S227(0) <='0';
          end if;
        if(oVar1S688(0)='1'  OR oVar1S689(0)='1'  OR oVar1S690(0)='1'  OR oVar1S691(0)='1'  )then
          oVar2S228(0) <='1';
          else
          oVar2S228(0) <='0';
          end if;
        if(oVar1S692(0)='1'  OR oVar1S693(0)='1'  OR oVar1S694(0)='1'  OR oVar1S695(0)='1'  )then
          oVar2S230(0) <='1';
          else
          oVar2S230(0) <='0';
          end if;
        if(oVar1S696(0)='1'  OR oVar1S697(0)='1'  OR oVar1S698(0)='1'  )then
          oVar2S231(0) <='1';
          else
          oVar2S231(0) <='0';
          end if;
        if(oVar1S699(0)='1'  OR oVar1S700(0)='1'  OR oVar1S701(0)='1'  OR oVar1S702(0)='1'  )then
          oVar2S232(0) <='1';
          else
          oVar2S232(0) <='0';
          end if;
        if(oVar1S703(0)='1'  OR oVar1S704(0)='1'  OR oVar1S705(0)='1'  )then
          oVar2S233(0) <='1';
          else
          oVar2S233(0) <='0';
          end if;
        if(oVar1S706(0)='1'  OR oVar1S707(0)='1'  OR oVar1S708(0)='1'  OR oVar1S709(0)='1'  )then
          oVar2S234(0) <='1';
          else
          oVar2S234(0) <='0';
          end if;
        if(oVar1S710(0)='1'  OR oVar1S711(0)='1'  OR oVar1S712(0)='1'  )then
          oVar2S235(0) <='1';
          else
          oVar2S235(0) <='0';
          end if;
        if(oVar1S714(0)='1'  OR oVar1S715(0)='1'  OR oVar1S716(0)='1'  OR oVar1S717(0)='1'  )then
          oVar2S237(0) <='1';
          else
          oVar2S237(0) <='0';
          end if;
        if(oVar1S718(0)='1'  OR oVar1S719(0)='1'  OR oVar1S720(0)='1'  )then
          oVar2S238(0) <='1';
          else
          oVar2S238(0) <='0';
          end if;
        if(oVar1S722(0)='1'  OR oVar1S723(0)='1'  OR oVar1S724(0)='1'  OR oVar1S725(0)='1'  )then
          oVar2S240(0) <='1';
          else
          oVar2S240(0) <='0';
          end if;
        if(oVar1S726(0)='1'  OR oVar1S727(0)='1'  OR oVar1S728(0)='1'  OR oVar1S729(0)='1'  )then
          oVar2S241(0) <='1';
          else
          oVar2S241(0) <='0';
          end if;
        if(oVar1S730(0)='1'  OR oVar1S731(0)='1'  OR oVar1S732(0)='1'  OR oVar1S733(0)='1'  )then
          oVar2S243(0) <='1';
          else
          oVar2S243(0) <='0';
          end if;
        if(oVar1S734(0)='1'  OR oVar1S735(0)='1'  OR oVar1S736(0)='1'  OR oVar1S737(0)='1'  )then
          oVar2S244(0) <='1';
          else
          oVar2S244(0) <='0';
          end if;
        if(oVar1S738(0)='1'  OR oVar1S739(0)='1'  OR oVar1S740(0)='1'  OR oVar1S741(0)='1'  )then
          oVar2S246(0) <='1';
          else
          oVar2S246(0) <='0';
          end if;
        if(oVar1S742(0)='1'  OR oVar1S743(0)='1'  OR oVar1S744(0)='1'  )then
          oVar2S247(0) <='1';
          else
          oVar2S247(0) <='0';
          end if;
        if(oVar1S746(0)='1'  OR oVar1S747(0)='1'  OR oVar1S748(0)='1'  OR oVar1S749(0)='1'  )then
          oVar2S249(0) <='1';
          else
          oVar2S249(0) <='0';
          end if;
        if(oVar1S750(0)='1'  OR oVar1S751(0)='1'  OR oVar1S752(0)='1'  OR oVar1S753(0)='1'  )then
          oVar2S250(0) <='1';
          else
          oVar2S250(0) <='0';
          end if;
        if(oVar1S754(0)='1'  )then
          oVar2S251(0) <='1';
          else
          oVar2S251(0) <='0';
          end if;
        if(oVar1S755(0)='1'  OR oVar1S756(0)='1'  OR oVar1S757(0)='1'  OR oVar1S758(0)='1'  )then
          oVar2S252(0) <='1';
          else
          oVar2S252(0) <='0';
          end if;
        if(oVar1S759(0)='1'  OR oVar1S760(0)='1'  OR oVar1S761(0)='1'  )then
          oVar2S253(0) <='1';
          else
          oVar2S253(0) <='0';
          end if;
        if(oVar1S762(0)='1'  OR oVar1S763(0)='1'  OR oVar1S764(0)='1'  OR oVar1S765(0)='1'  )then
          oVar2S254(0) <='1';
          else
          oVar2S254(0) <='0';
          end if;
        if(oVar1S766(0)='1'  OR oVar1S767(0)='1'  OR oVar1S768(0)='1'  OR oVar1S769(0)='1'  )then
          oVar2S255(0) <='1';
          else
          oVar2S255(0) <='0';
          end if;
        if(oVar1S770(0)='1'  OR oVar1S771(0)='1'  )then
          oVar2S256(0) <='1';
          else
          oVar2S256(0) <='0';
          end if;
        if(oVar1S772(0)='1'  OR oVar1S773(0)='1'  OR oVar1S774(0)='1'  OR oVar1S775(0)='1'  )then
          oVar2S257(0) <='1';
          else
          oVar2S257(0) <='0';
          end if;
        if(oVar1S776(0)='1'  OR oVar1S777(0)='1'  OR oVar1S778(0)='1'  )then
          oVar2S258(0) <='1';
          else
          oVar2S258(0) <='0';
          end if;
        if(oVar1S779(0)='1'  OR oVar1S780(0)='1'  OR oVar1S781(0)='1'  OR oVar1S782(0)='1'  )then
          oVar2S259(0) <='1';
          else
          oVar2S259(0) <='0';
          end if;
        if(oVar1S783(0)='1'  OR oVar1S784(0)='1'  OR oVar1S785(0)='1'  )then
          oVar2S260(0) <='1';
          else
          oVar2S260(0) <='0';
          end if;
        if(oVar1S786(0)='1'  OR oVar1S787(0)='1'  OR oVar1S788(0)='1'  OR oVar1S789(0)='1'  )then
          oVar2S261(0) <='1';
          else
          oVar2S261(0) <='0';
          end if;
        if(oVar1S790(0)='1'  OR oVar1S791(0)='1'  OR oVar1S792(0)='1'  )then
          oVar2S262(0) <='1';
          else
          oVar2S262(0) <='0';
          end if;
        if(oVar1S793(0)='1'  OR oVar1S794(0)='1'  OR oVar1S795(0)='1'  OR oVar1S796(0)='1'  )then
          oVar2S263(0) <='1';
          else
          oVar2S263(0) <='0';
          end if;
        if(oVar1S797(0)='1'  OR oVar1S798(0)='1'  OR oVar1S799(0)='1'  OR oVar1S800(0)='1'  )then
          oVar2S264(0) <='1';
          else
          oVar2S264(0) <='0';
          end if;
        if(oVar1S801(0)='1'  OR oVar1S802(0)='1'  OR oVar1S803(0)='1'  OR oVar1S804(0)='1'  )then
          oVar2S266(0) <='1';
          else
          oVar2S266(0) <='0';
          end if;
        if(oVar1S805(0)='1'  OR oVar1S806(0)='1'  OR oVar1S807(0)='1'  OR oVar1S808(0)='1'  )then
          oVar2S267(0) <='1';
          else
          oVar2S267(0) <='0';
          end if;
        if(oVar1S809(0)='1'  )then
          oVar2S268(0) <='1';
          else
          oVar2S268(0) <='0';
          end if;
        if(oVar1S810(0)='1'  OR oVar1S811(0)='1'  OR oVar1S812(0)='1'  OR oVar1S813(0)='1'  )then
          oVar2S269(0) <='1';
          else
          oVar2S269(0) <='0';
          end if;
        if(oVar1S814(0)='1'  OR oVar1S815(0)='1'  )then
          oVar2S270(0) <='1';
          else
          oVar2S270(0) <='0';
          end if;
        if(oVar1S816(0)='1'  OR oVar1S817(0)='1'  OR oVar1S818(0)='1'  OR oVar1S819(0)='1'  )then
          oVar2S271(0) <='1';
          else
          oVar2S271(0) <='0';
          end if;
        if(oVar1S820(0)='1'  OR oVar1S821(0)='1'  OR oVar1S822(0)='1'  OR oVar1S823(0)='1'  )then
          oVar2S272(0) <='1';
          else
          oVar2S272(0) <='0';
          end if;
        if(oVar1S824(0)='1'  OR oVar1S825(0)='1'  OR oVar1S826(0)='1'  OR oVar1S827(0)='1'  )then
          oVar2S274(0) <='1';
          else
          oVar2S274(0) <='0';
          end if;
        if(oVar1S828(0)='1'  OR oVar1S829(0)='1'  OR oVar1S830(0)='1'  OR oVar1S831(0)='1'  )then
          oVar2S275(0) <='1';
          else
          oVar2S275(0) <='0';
          end if;
        if(oVar1S832(0)='1'  OR oVar1S833(0)='1'  OR oVar1S834(0)='1'  OR oVar1S835(0)='1'  )then
          oVar2S277(0) <='1';
          else
          oVar2S277(0) <='0';
          end if;
        if(oVar1S836(0)='1'  OR oVar1S837(0)='1'  OR oVar1S838(0)='1'  )then
          oVar2S278(0) <='1';
          else
          oVar2S278(0) <='0';
          end if;
        if(oVar1S839(0)='1'  OR oVar1S840(0)='1'  OR oVar1S841(0)='1'  OR oVar1S842(0)='1'  )then
          oVar2S279(0) <='1';
          else
          oVar2S279(0) <='0';
          end if;
        if(oVar1S843(0)='1'  OR oVar1S844(0)='1'  OR oVar1S845(0)='1'  OR oVar1S846(0)='1'  )then
          oVar2S280(0) <='1';
          else
          oVar2S280(0) <='0';
          end if;
        if(oVar1S847(0)='1'  OR oVar1S848(0)='1'  OR oVar1S849(0)='1'  OR oVar1S850(0)='1'  )then
          oVar2S282(0) <='1';
          else
          oVar2S282(0) <='0';
          end if;
        if(oVar1S851(0)='1'  OR oVar1S852(0)='1'  OR oVar1S853(0)='1'  OR oVar1S854(0)='1'  )then
          oVar2S283(0) <='1';
          else
          oVar2S283(0) <='0';
          end if;
        if(oVar1S856(0)='1'  OR oVar1S857(0)='1'  OR oVar1S858(0)='1'  OR oVar1S859(0)='1'  )then
          oVar2S285(0) <='1';
          else
          oVar2S285(0) <='0';
          end if;
        if(oVar1S860(0)='1'  OR oVar1S861(0)='1'  )then
          oVar2S286(0) <='1';
          else
          oVar2S286(0) <='0';
          end if;
        if(oVar1S862(0)='1'  OR oVar1S863(0)='1'  OR oVar1S864(0)='1'  OR oVar1S865(0)='1'  )then
          oVar2S287(0) <='1';
          else
          oVar2S287(0) <='0';
          end if;
        if(oVar1S866(0)='1'  OR oVar1S867(0)='1'  )then
          oVar2S288(0) <='1';
          else
          oVar2S288(0) <='0';
          end if;
        if(oVar1S869(0)='1'  OR oVar1S870(0)='1'  OR oVar1S871(0)='1'  OR oVar1S872(0)='1'  )then
          oVar2S289(0) <='1';
          else
          oVar2S289(0) <='0';
          end if;
        if(oVar1S873(0)='1'  OR oVar1S874(0)='1'  )then
          oVar2S290(0) <='1';
          else
          oVar2S290(0) <='0';
          end if;
        if(oVar1S875(0)='1'  OR oVar1S876(0)='1'  OR oVar1S877(0)='1'  OR oVar1S878(0)='1'  )then
          oVar2S291(0) <='1';
          else
          oVar2S291(0) <='0';
          end if;
        if(oVar1S879(0)='1'  OR oVar1S880(0)='1'  )then
          oVar2S292(0) <='1';
          else
          oVar2S292(0) <='0';
          end if;
        if(oVar1S882(0)='1'  OR oVar1S883(0)='1'  OR oVar1S884(0)='1'  OR oVar1S885(0)='1'  )then
          oVar2S293(0) <='1';
          else
          oVar2S293(0) <='0';
          end if;
        if(oVar1S886(0)='1'  )then
          oVar2S294(0) <='1';
          else
          oVar2S294(0) <='0';
          end if;
        if(oVar1S887(0)='1'  OR oVar1S888(0)='1'  OR oVar1S889(0)='1'  OR oVar1S890(0)='1'  )then
          oVar2S295(0) <='1';
          else
          oVar2S295(0) <='0';
          end if;
        if(oVar1S891(0)='1'  OR oVar1S892(0)='1'  OR oVar1S893(0)='1'  )then
          oVar2S296(0) <='1';
          else
          oVar2S296(0) <='0';
          end if;
        if(oVar1S895(0)='1'  OR oVar1S896(0)='1'  OR oVar1S897(0)='1'  OR oVar1S898(0)='1'  )then
          oVar2S298(0) <='1';
          else
          oVar2S298(0) <='0';
          end if;
        if(oVar1S899(0)='1'  OR oVar1S900(0)='1'  )then
          oVar2S299(0) <='1';
          else
          oVar2S299(0) <='0';
          end if;
        if(oVar1S901(0)='1'  OR oVar1S902(0)='1'  OR oVar1S903(0)='1'  OR oVar1S904(0)='1'  )then
          oVar2S300(0) <='1';
          else
          oVar2S300(0) <='0';
          end if;
        if(oVar1S905(0)='1'  OR oVar1S906(0)='1'  )then
          oVar2S301(0) <='1';
          else
          oVar2S301(0) <='0';
          end if;
        if(oVar1S907(0)='1'  OR oVar1S908(0)='1'  OR oVar1S909(0)='1'  OR oVar1S910(0)='1'  )then
          oVar2S302(0) <='1';
          else
          oVar2S302(0) <='0';
          end if;
        if(oVar1S911(0)='1'  OR oVar1S912(0)='1'  OR oVar1S913(0)='1'  OR oVar1S914(0)='1'  )then
          oVar2S304(0) <='1';
          else
          oVar2S304(0) <='0';
          end if;
        if(oVar1S915(0)='1'  OR oVar1S916(0)='1'  OR oVar1S917(0)='1'  )then
          oVar2S305(0) <='1';
          else
          oVar2S305(0) <='0';
          end if;
        if(oVar1S918(0)='1'  OR oVar1S919(0)='1'  OR oVar1S920(0)='1'  OR oVar1S921(0)='1'  )then
          oVar2S306(0) <='1';
          else
          oVar2S306(0) <='0';
          end if;
        if(oVar1S922(0)='1'  OR oVar1S923(0)='1'  OR oVar1S924(0)='1'  OR oVar1S925(0)='1'  )then
          oVar2S307(0) <='1';
          else
          oVar2S307(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV5 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar2S254(0)='1' OR oVar2S255(0)='1' OR oVar2S256(0)='1' )then
          ADDM4K3S8(0)<='1';
          else
          ADDM4K3S8(0)<='0';
          end if;
        if(oVar2S257(0)='1' OR oVar2S258(0)='1' )then
          ADDM4K3S8(1)<='1';
          else
          ADDM4K3S8(1)<='0';
          end if;
        if(oVar2S261(0)='1' OR oVar2S262(0)='1' )then
          ADDM4K3S8(2)<='1';
          else
          ADDM4K3S8(2)<='0';
          end if;
        if(oVar2S153(0)='1' OR oVar2S154(0)='1' )then
          ADDM4K3S8(3)<='1';
          else
          ADDM4K3S8(3)<='0';
          end if;
        if(oVar2S182(0)='1' OR oVar2S183(0)='1' )then
          ADDM4K3S8(4)<='1';
          else
          ADDM4K3S8(4)<='0';
          end if;
        if(oVar2S184(0)='1' OR oVar2S185(0)='1' )then
          ADDM4K3S8(5)<='1';
          else
          ADDM4K3S8(5)<='0';
          end if;
        if(oVar2S103(0)='1' OR oVar2S104(0)='1' )then
          ADDM4K3S8(6)<='1';
          else
          ADDM4K3S8(6)<='0';
          end if;
        if(oVar2S123(0)='1' OR oVar2S124(0)='1' )then
          ADDM4K3S8(7)<='1';
          else
          ADDM4K3S8(7)<='0';
          end if;
        if(oVar2S282(0)='1' OR oVar2S283(0)='1' )then
          ADDM4K3S9(0)<='1';
          else
          ADDM4K3S9(0)<='0';
          end if;
        if(oVar2S69(0)='1' OR oVar2S70(0)='1' )then
          ADDM4K3S9(1)<='1';
          else
          ADDM4K3S9(1)<='0';
          end if;
        if(oVar2S146(0)='1' OR oVar2S147(0)='1' )then
          ADDM4K3S9(2)<='1';
          else
          ADDM4K3S9(2)<='0';
          end if;
        if(oVar2S91(0)='1' OR oVar2S92(0)='1' )then
          ADDM4K3S9(3)<='1';
          else
          ADDM4K3S9(3)<='0';
          end if;
        if(oVar2S274(0)='1' OR oVar2S275(0)='1' )then
          ADDM4K3S9(4)<='1';
          else
          ADDM4K3S9(4)<='0';
          end if;
        if(oVar2S190(0)='1' OR oVar2S191(0)='1' )then
          ADDM4K3S9(5)<='1';
          else
          ADDM4K3S9(5)<='0';
          end if;
        if(oVar2S110(0)='1' OR oVar2S111(0)='1' )then
          ADDM4K3S9(6)<='1';
          else
          ADDM4K3S9(6)<='0';
          end if;
        if(oVar2S67(0)='1' OR oVar2S68(0)='1' )then
          ADDM4K3S9(7)<='1';
          else
          ADDM4K3S9(7)<='0';
          end if;
        if(oVar2S44(0)='1' OR oVar2S45(0)='1' )then
          ADDM4K3S12(0)<='1';
          else
          ADDM4K3S12(0)<='0';
          end if;
        if(oVar2S36(0)='1' OR oVar2S37(0)='1' )then
          ADDM4K3S12(1)<='1';
          else
          ADDM4K3S12(1)<='0';
          end if;
        if(oVar2S64(0)='1' OR oVar2S65(0)='1' )then
          ADDM4K3S12(2)<='1';
          else
          ADDM4K3S12(2)<='0';
          end if;
        if(oVar2S46(0)='1' OR oVar2S47(0)='1' )then
          ADDM4K3S12(3)<='1';
          else
          ADDM4K3S12(3)<='0';
          end if;
        if(oVar2S55(0)='1' OR oVar2S56(0)='1' )then
          ADDM4K3S12(4)<='1';
          else
          ADDM4K3S12(4)<='0';
          end if;
        if(oVar2S82(0)='1' OR oVar2S83(0)='1' )then
          ADDM4K3S12(5)<='1';
          else
          ADDM4K3S12(5)<='0';
          end if;
        if(oVar2S53(0)='1' OR oVar2S54(0)='1' )then
          ADDM4K3S12(6)<='1';
          else
          ADDM4K3S12(6)<='0';
          end if;
        if(oVar2S79(0)='1' OR oVar2S80(0)='1' )then
          ADDM4K3S12(7)<='1';
          else
          ADDM4K3S12(7)<='0';
          end if;
        if(oVar2S85(0)='1' OR oVar2S86(0)='1' )then
          ADDM4K3S13(0)<='1';
          else
          ADDM4K3S13(0)<='0';
          end if;
        if(oVar2S74(0)='1' OR oVar2S75(0)='1' )then
          ADDM4K3S13(1)<='1';
          else
          ADDM4K3S13(1)<='0';
          end if;
        if(oVar2S61(0)='1' OR oVar2S62(0)='1' )then
          ADDM4K3S13(2)<='1';
          else
          ADDM4K3S13(2)<='0';
          end if;
        if(oVar2S39(0)='1' OR oVar2S40(0)='1' )then
          ADDM4K3S13(3)<='1';
          else
          ADDM4K3S13(3)<='0';
          end if;
        if(oVar2S57(0)='1' OR oVar2S58(0)='1' )then
          ADDM4K3S13(4)<='1';
          else
          ADDM4K3S13(4)<='0';
          end if;
        if(oVar2S48(0)='1' OR oVar2S49(0)='1' )then
          ADDM4K3S13(5)<='1';
          else
          ADDM4K3S13(5)<='0';
          end if;
        if(oVar2S42(0)='1' OR oVar2S43(0)='1' )then
          ADDM4K3S13(6)<='1';
          else
          ADDM4K3S13(6)<='0';
          end if;
        if(oVar2S59(0)='1' OR oVar2S60(0)='1' )then
          ADDM4K3S13(7)<='1';
          else
          ADDM4K3S13(7)<='0';
          end if;
        if(oVar2S162(0)='1' OR oVar2S163(0)='1' )then
          ADDM4K3S10(0)<='1';
          else
          ADDM4K3S10(0)<='0';
          end if;
        if(oVar2S94(0)='1' OR oVar2S95(0)='1' )then
          ADDM4K3S10(1)<='1';
          else
          ADDM4K3S10(1)<='0';
          end if;
        if(oVar2S176(0)='1' OR oVar2S177(0)='1' )then
          ADDM4K3S10(2)<='1';
          else
          ADDM4K3S10(2)<='0';
          end if;
        if(oVar2S121(0)='1' OR oVar2S122(0)='1' )then
          ADDM4K3S10(3)<='1';
          else
          ADDM4K3S10(3)<='0';
          end if;
        if(oVar2S148(0)='1' OR oVar2S149(0)='1' )then
          ADDM4K3S10(4)<='1';
          else
          ADDM4K3S10(4)<='0';
          end if;
        if(oVar2S108(0)='1' OR oVar2S109(0)='1' )then
          ADDM4K3S10(5)<='1';
          else
          ADDM4K3S10(5)<='0';
          end if;
        if(oVar2S187(0)='1' OR oVar2S188(0)='1' )then
          ADDM4K3S10(6)<='1';
          else
          ADDM4K3S10(6)<='0';
          end if;
        if(oVar2S150(0)='1' OR oVar2S151(0)='1' OR oVar2S152(0)='1' )then
          ADDM4K3S10(7)<='1';
          else
          ADDM4K3S10(7)<='0';
          end if;
        if(oVar2S173(0)='1' OR oVar2S174(0)='1' )then
          ADDM4K3S11(0)<='1';
          else
          ADDM4K3S11(0)<='0';
          end if;
        if(oVar2S116(0)='1' OR oVar2S117(0)='1' )then
          ADDM4K3S11(1)<='1';
          else
          ADDM4K3S11(1)<='0';
          end if;
        if(oVar2S97(0)='1' OR oVar2S98(0)='1' )then
          ADDM4K3S11(2)<='1';
          else
          ADDM4K3S11(2)<='0';
          end if;
        if(oVar2S87(0)='1' OR oVar2S88(0)='1' )then
          ADDM4K3S11(3)<='1';
          else
          ADDM4K3S11(3)<='0';
          end if;
        if(oVar2S100(0)='1' OR oVar2S101(0)='1' )then
          ADDM4K3S11(4)<='1';
          else
          ADDM4K3S11(4)<='0';
          end if;
        if(oVar2S119(0)='1' OR oVar2S120(0)='1' )then
          ADDM4K3S11(5)<='1';
          else
          ADDM4K3S11(5)<='0';
          end if;
        if(oVar2S71(0)='1' OR oVar2S72(0)='1' OR oVar2S73(0)='1' )then
          ADDM4K3S11(6)<='1';
          else
          ADDM4K3S11(6)<='0';
          end if;
        if(oVar2S51(0)='1' OR oVar2S52(0)='1' )then
          ADDM4K3S11(7)<='1';
          else
          ADDM4K3S11(7)<='0';
          end if;
        if(oVar2S76(0)='1' OR oVar2S77(0)='1' OR oVar2S78(0)='1' )then
          ADDM4K3S14(0)<='1';
          else
          ADDM4K3S14(0)<='0';
          end if;
        if(oVar2S33(0)='1' OR oVar2S34(0)='1' )then
          ADDM4K3S14(1)<='1';
          else
          ADDM4K3S14(1)<='0';
          end if;
        if(oVar2S28(0)='1' OR oVar2S29(0)='1' )then
          ADDM4K3S14(2)<='1';
          else
          ADDM4K3S14(2)<='0';
          end if;
        if(oVar2S25(0)='1' OR oVar2S26(0)='1' )then
          ADDM4K3S14(3)<='1';
          else
          ADDM4K3S14(3)<='0';
          end if;
        if(oVar2S30(0)='1' OR oVar2S31(0)='1' )then
          ADDM4K3S14(4)<='1';
          else
          ADDM4K3S14(4)<='0';
          end if;
        if(oVar2S20(0)='1' OR oVar2S21(0)='1' )then
          ADDM4K3S14(5)<='1';
          else
          ADDM4K3S14(5)<='0';
          end if;
        if(oVar2S17(0)='1' OR oVar2S18(0)='1' )then
          ADDM4K3S14(6)<='1';
          else
          ADDM4K3S14(6)<='0';
          end if;
        if(oVar2S9(0)='1' OR oVar2S10(0)='1' )then
          ADDM4K3S14(7)<='1';
          else
          ADDM4K3S14(7)<='0';
          end if;
        if(oVar2S22(0)='1' OR oVar2S23(0)='1' OR oVar2S24(0)='1' )then
          ADDM4K3S15(0)<='1';
          else
          ADDM4K3S15(0)<='0';
          end if;
        if(oVar2S15(0)='1' OR oVar2S16(0)='1' )then
          ADDM4K3S15(1)<='1';
          else
          ADDM4K3S15(1)<='0';
          end if;
        if(oVar2S13(0)='1' OR oVar2S14(0)='1' )then
          ADDM4K3S15(2)<='1';
          else
          ADDM4K3S15(2)<='0';
          end if;
        if(oVar2S11(0)='1' OR oVar2S12(0)='1' )then
          ADDM4K3S15(3)<='1';
          else
          ADDM4K3S15(3)<='0';
          end if;
        if(oVar2S4(0)='1' OR oVar2S5(0)='1' )then
          ADDM4K3S15(4)<='1';
          else
          ADDM4K3S15(4)<='0';
          end if;
        if(oVar2S6(0)='1' OR oVar2S7(0)='1' )then
          ADDM4K3S15(5)<='1';
          else
          ADDM4K3S15(5)<='0';
          end if;
        if(oVar2S2(0)='1' OR oVar2S3(0)='1' )then
          ADDM4K3S15(6)<='1';
          else
          ADDM4K3S15(6)<='0';
          end if;
        if(oVar2S0(0)='1' OR oVar2S1(0)='1' )then
          ADDM4K3S15(7)<='1';
          else
          ADDM4K3S15(7)<='0';
          end if;
        if(oVar2S216(0)='1' OR oVar2S217(0)='1' )then
          ADDM4K3S2(0)<='1';
          else
          ADDM4K3S2(0)<='0';
          end if;
        if(oVar2S237(0)='1' OR oVar2S238(0)='1' )then
          ADDM4K3S2(1)<='1';
          else
          ADDM4K3S2(1)<='0';
          end if;
        if(oVar2S287(0)='1' OR oVar2S288(0)='1' )then
          ADDM4K3S2(2)<='1';
          else
          ADDM4K3S2(2)<='0';
          end if;
        if(oVar2S206(0)='1' OR oVar2S207(0)='1' )then
          ADDM4K3S2(3)<='1';
          else
          ADDM4K3S2(3)<='0';
          end if;
        if(oVar2S193(0)='1' OR oVar2S194(0)='1' )then
          ADDM4K3S2(4)<='1';
          else
          ADDM4K3S2(4)<='0';
          end if;
        if(oVar2S134(0)='1' OR oVar2S135(0)='1' )then
          ADDM4K3S2(5)<='1';
          else
          ADDM4K3S2(5)<='0';
          end if;
        if(oVar2S140(0)='1' OR oVar2S141(0)='1' )then
          ADDM4K3S2(6)<='1';
          else
          ADDM4K3S2(6)<='0';
          end if;
        if(oVar2S208(0)='1' OR oVar2S209(0)='1' )then
          ADDM4K3S2(7)<='1';
          else
          ADDM4K3S2(7)<='0';
          end if;
        if(oVar2S234(0)='1' OR oVar2S235(0)='1' )then
          ADDM4K3S3(0)<='1';
          else
          ADDM4K3S3(0)<='0';
          end if;
        if(oVar2S271(0)='1' OR oVar2S272(0)='1' )then
          ADDM4K3S3(1)<='1';
          else
          ADDM4K3S3(1)<='0';
          end if;
        if(oVar2S138(0)='1' OR oVar2S139(0)='1' )then
          ADDM4K3S3(2)<='1';
          else
          ADDM4K3S3(2)<='0';
          end if;
        if(oVar2S269(0)='1' OR oVar2S270(0)='1' )then
          ADDM4K3S3(3)<='1';
          else
          ADDM4K3S3(3)<='0';
          end if;
        if(oVar2S195(0)='1' OR oVar2S196(0)='1' )then
          ADDM4K3S3(4)<='1';
          else
          ADDM4K3S3(4)<='0';
          end if;
        if(oVar2S232(0)='1' OR oVar2S233(0)='1' )then
          ADDM4K3S3(5)<='1';
          else
          ADDM4K3S3(5)<='0';
          end if;
        if(oVar2S89(0)='1' OR oVar2S90(0)='1' )then
          ADDM4K3S3(6)<='1';
          else
          ADDM4K3S3(6)<='0';
          end if;
        if(oVar2S204(0)='1' OR oVar2S205(0)='1' )then
          ADDM4K3S3(7)<='1';
          else
          ADDM4K3S3(7)<='0';
          end if;
        if(oVar2S252(0)='1' OR oVar2S253(0)='1' )then
          ADDM4K3S4(0)<='1';
          else
          ADDM4K3S4(0)<='0';
          end if;
        if(oVar2S142(0)='1' OR oVar2S143(0)='1' )then
          ADDM4K3S4(1)<='1';
          else
          ADDM4K3S4(1)<='0';
          end if;
        if(oVar2S136(0)='1' OR oVar2S137(0)='1' )then
          ADDM4K3S4(2)<='1';
          else
          ADDM4K3S4(2)<='0';
          end if;
        if(oVar2S114(0)='1' OR oVar2S115(0)='1' )then
          ADDM4K3S4(3)<='1';
          else
          ADDM4K3S4(3)<='0';
          end if;
        if(oVar2S199(0)='1' OR oVar2S200(0)='1' )then
          ADDM4K3S4(4)<='1';
          else
          ADDM4K3S4(4)<='0';
          end if;
        if(oVar2S279(0)='1' OR oVar2S280(0)='1' )then
          ADDM4K3S4(5)<='1';
          else
          ADDM4K3S4(5)<='0';
          end if;
        if(oVar2S259(0)='1' OR oVar2S260(0)='1' )then
          ADDM4K3S4(6)<='1';
          else
          ADDM4K3S4(6)<='0';
          end if;
        if(oVar2S201(0)='1' OR oVar2S202(0)='1' )then
          ADDM4K3S4(7)<='1';
          else
          ADDM4K3S4(7)<='0';
          end if;
        if(oVar2S144(0)='1' OR oVar2S145(0)='1' )then
          ADDM4K3S5(0)<='1';
          else
          ADDM4K3S5(0)<='0';
          end if;
        if(oVar2S263(0)='1' OR oVar2S264(0)='1' )then
          ADDM4K3S5(1)<='1';
          else
          ADDM4K3S5(1)<='0';
          end if;
        if(oVar2S249(0)='1' OR oVar2S250(0)='1' OR oVar2S251(0)='1' )then
          ADDM4K3S5(2)<='1';
          else
          ADDM4K3S5(2)<='0';
          end if;
        if(oVar2S246(0)='1' OR oVar2S247(0)='1' )then
          ADDM4K3S5(3)<='1';
          else
          ADDM4K3S5(3)<='0';
          end if;
        if(oVar2S155(0)='1' OR oVar2S156(0)='1' )then
          ADDM4K3S5(4)<='1';
          else
          ADDM4K3S5(4)<='0';
          end if;
        if(oVar2S240(0)='1' OR oVar2S241(0)='1' )then
          ADDM4K3S5(5)<='1';
          else
          ADDM4K3S5(5)<='0';
          end if;
        if(oVar2S168(0)='1' OR oVar2S169(0)='1' )then
          ADDM4K3S5(6)<='1';
          else
          ADDM4K3S5(6)<='0';
          end if;
        if(oVar2S170(0)='1' OR oVar2S171(0)='1' )then
          ADDM4K3S5(7)<='1';
          else
          ADDM4K3S5(7)<='0';
          end if;
        if(oVar2S213(0)='1' OR oVar2S214(0)='1' )then
          ADDM4K3S6(0)<='1';
          else
          ADDM4K3S6(0)<='0';
          end if;
        if(oVar2S266(0)='1' OR oVar2S267(0)='1' OR oVar2S268(0)='1' )then
          ADDM4K3S6(1)<='1';
          else
          ADDM4K3S6(1)<='0';
          end if;
        if(oVar2S157(0)='1' OR oVar2S158(0)='1' )then
          ADDM4K3S6(2)<='1';
          else
          ADDM4K3S6(2)<='0';
          end if;
        if(oVar2S106(0)='1' OR oVar2S107(0)='1' )then
          ADDM4K3S6(3)<='1';
          else
          ADDM4K3S6(3)<='0';
          end if;
        if(oVar2S285(0)='1' OR oVar2S286(0)='1' )then
          ADDM4K3S6(4)<='1';
          else
          ADDM4K3S6(4)<='0';
          end if;
        if(oVar2S130(0)='1' OR oVar2S131(0)='1' )then
          ADDM4K3S6(5)<='1';
          else
          ADDM4K3S6(5)<='0';
          end if;
        if(oVar2S179(0)='1' OR oVar2S180(0)='1' )then
          ADDM4K3S6(6)<='1';
          else
          ADDM4K3S6(6)<='0';
          end if;
        if(oVar2S112(0)='1' OR oVar2S113(0)='1' )then
          ADDM4K3S6(7)<='1';
          else
          ADDM4K3S6(7)<='0';
          end if;
        if(oVar2S277(0)='1' OR oVar2S278(0)='1' )then
          ADDM4K3S7(0)<='1';
          else
          ADDM4K3S7(0)<='0';
          end if;
        if(oVar2S243(0)='1' OR oVar2S244(0)='1' )then
          ADDM4K3S7(1)<='1';
          else
          ADDM4K3S7(1)<='0';
          end if;
        if(oVar2S211(0)='1' OR oVar2S212(0)='1' )then
          ADDM4K3S7(2)<='1';
          else
          ADDM4K3S7(2)<='0';
          end if;
        if(oVar2S197(0)='1' OR oVar2S198(0)='1' )then
          ADDM4K3S7(3)<='1';
          else
          ADDM4K3S7(3)<='0';
          end if;
        if(oVar2S165(0)='1' OR oVar2S166(0)='1' )then
          ADDM4K3S7(4)<='1';
          else
          ADDM4K3S7(4)<='0';
          end if;
        if(oVar2S128(0)='1' OR oVar2S129(0)='1' )then
          ADDM4K3S7(5)<='1';
          else
          ADDM4K3S7(5)<='0';
          end if;
        if(oVar2S132(0)='1' OR oVar2S133(0)='1' )then
          ADDM4K3S7(6)<='1';
          else
          ADDM4K3S7(6)<='0';
          end if;
        if(oVar2S125(0)='1' OR oVar2S126(0)='1' )then
          ADDM4K3S7(7)<='1';
          else
          ADDM4K3S7(7)<='0';
          end if;
        if(oVar2S300(0)='1' OR oVar2S301(0)='1' )then
          ADDM4K3S0(0)<='1';
          else
          ADDM4K3S0(0)<='0';
          end if;
        if(oVar2S306(0)='1' OR oVar2S307(0)='1' )then
          ADDM4K3S0(1)<='1';
          else
          ADDM4K3S0(1)<='0';
          end if;
        if(oVar2S302(0)='1' )then
          ADDM4K3S0(2)<='1';
          else
          ADDM4K3S0(2)<='0';
          end if;
        if(oVar2S304(0)='1' OR oVar2S305(0)='1' )then
          ADDM4K3S0(3)<='1';
          else
          ADDM4K3S0(3)<='0';
          end if;
        if(oVar2S225(0)='1' OR oVar2S226(0)='1' )then
          ADDM4K3S0(4)<='1';
          else
          ADDM4K3S0(4)<='0';
          end if;
        if(oVar2S298(0)='1' OR oVar2S299(0)='1' )then
          ADDM4K3S0(5)<='1';
          else
          ADDM4K3S0(5)<='0';
          end if;
        if(oVar2S291(0)='1' OR oVar2S292(0)='1' )then
          ADDM4K3S0(6)<='1';
          else
          ADDM4K3S0(6)<='0';
          end if;
        if(oVar2S222(0)='1' OR oVar2S223(0)='1' )then
          ADDM4K3S0(7)<='1';
          else
          ADDM4K3S0(7)<='0';
          end if;
        if(oVar2S293(0)='1' OR oVar2S294(0)='1' )then
          ADDM4K3S1(0)<='1';
          else
          ADDM4K3S1(0)<='0';
          end if;
        if(oVar2S227(0)='1' OR oVar2S228(0)='1' )then
          ADDM4K3S1(1)<='1';
          else
          ADDM4K3S1(1)<='0';
          end if;
        if(oVar2S295(0)='1' OR oVar2S296(0)='1' )then
          ADDM4K3S1(2)<='1';
          else
          ADDM4K3S1(2)<='0';
          end if;
        if(oVar2S220(0)='1' OR oVar2S221(0)='1' )then
          ADDM4K3S1(3)<='1';
          else
          ADDM4K3S1(3)<='0';
          end if;
        if(oVar2S218(0)='1' OR oVar2S219(0)='1' )then
          ADDM4K3S1(4)<='1';
          else
          ADDM4K3S1(4)<='0';
          end if;
        if(oVar2S230(0)='1' OR oVar2S231(0)='1' )then
          ADDM4K3S1(5)<='1';
          else
          ADDM4K3S1(5)<='0';
          end if;
        if(oVar2S289(0)='1' OR oVar2S290(0)='1' )then
          ADDM4K3S1(6)<='1';
          else
          ADDM4K3S1(6)<='0';
          end if;
        if(oVar2S159(0)='1' OR oVar2S160(0)='1' )then
          ADDM4K3S1(7)<='1';
          else
          ADDM4K3S1(7)<='0';
          end if;
 end if;
end process;
ADDM4K3S8c : ADDM4K3S8RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S8,
                q    => aVar3S8
    );
ADDM4K3S9c : ADDM4K3S9RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S9,
                q    => aVar3S9
    );
ADDM4K3S12c : ADDM4K3S12RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S12,
                q    => aVar3S12
    );
ADDM4K3S13c : ADDM4K3S13RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S13,
                q    => aVar3S13
    );
ADDM4K3S10c : ADDM4K3S10RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S10,
                q    => aVar3S10
    );
ADDM4K3S11c : ADDM4K3S11RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S11,
                q    => aVar3S11
    );
ADDM4K3S14c : ADDM4K3S14RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S14,
                q    => aVar3S14
    );
ADDM4K3S15c : ADDM4K3S15RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S15,
                q    => aVar3S15
    );
ADDM4K3S2c : ADDM4K3S2RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S2,
                q    => aVar3S2
    );
ADDM4K3S3c : ADDM4K3S3RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S3,
                q    => aVar3S3
    );
ADDM4K3S4c : ADDM4K3S4RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S4,
                q    => aVar3S4
    );
ADDM4K3S5c : ADDM4K3S5RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S5,
                q    => aVar3S5
    );
ADDM4K3S6c : ADDM4K3S6RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S6,
                q    => aVar3S6
    );
ADDM4K3S7c : ADDM4K3S7RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S7,
                q    => aVar3S7
    );
ADDM4K3S0c : ADDM4K3S0RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S0,
                q    => aVar3S0
    );
ADDM4K3S1c : ADDM4K3S1RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S1,
                q    => aVar3S1
    );
Adder_1: Adder_type
port map(
dataa => aVar3S0, 
datab => aVar3S1, 
result => aVar4S0
);

Adder_2: Adder_type
port map(
dataa => aVar3S2, 
datab => aVar3S3, 
result => aVar4S1
);

Adder_3: Adder_type
port map(
dataa => aVar3S4, 
datab => aVar3S5, 
result => aVar4S2
);

Adder_4: Adder_type
port map(
dataa => aVar3S6, 
datab => aVar3S7, 
result => aVar4S3
);

Adder_5: Adder_type
port map(
dataa => aVar3S8, 
datab => aVar3S9, 
result => aVar4S4
);

Adder_6: Adder_type
port map(
dataa => aVar3S10, 
datab => aVar3S11, 
result => aVar4S5
);

Adder_7: Adder_type
port map(
dataa => aVar3S12, 
datab => aVar3S13, 
result => aVar4S6
);

Adder_8: Adder_type
port map(
dataa => aVar3S14, 
datab => aVar3S15, 
result => aVar4S7
);

Adder_9: Adder_type
port map(
dataa => aVar4S0, 
datab => aVar4S1, 
result => aVar5S0
);

Adder_10: Adder_type
port map(
dataa => aVar4S2, 
datab => aVar4S3, 
result => aVar5S1
);

Adder_11: Adder_type
port map(
dataa => aVar4S4, 
datab => aVar4S5, 
result => aVar5S2
);

Adder_12: Adder_type
port map(
dataa => aVar4S6, 
datab => aVar4S7, 
result => aVar5S3
);

Adder_13: Adder_type
port map(
dataa => aVar5S0, 
datab => aVar5S1, 
result => aVar6S0
);

Adder_14: Adder_type
port map(
dataa => aVar5S2, 
datab => aVar5S3, 
result => aVar6S1
);

Adder_15: Adder_type
port map(
dataa => aVar6S0, 
datab => aVar6S1, 
result => aVar7S0
);

end rtl;
