LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY code_450 IS
   PORT(
      --*************************************************
      -- V1495 Front Panel Ports (PORT A,B,C,G)
      --*************************************************
      A_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In A (32 x LVDS/ECL)
      B_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In B (32 x LVDS/ECL)
      D_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In D (32 x LVDS/ECL)
      E_DIN_L       : IN     std_logic_vector (31 DOWNTO 0);  -- In E (32 x LVDS/ECL)
      F_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- OUT F (32 x LVDS/ECL)
      C_DOUT_L      : OUT    std_logic_vector (31 DOWNTO 0);  -- Out C (32 x LVDS)
      c1            : IN STD_LOGIC                            -- the PLL1 output
   );
END code_450 ;
ARCHITECTURE rtl OF code_450 IS
	signal A     : std_logic_vector(31 downto 0);
	signal B     : std_logic_vector(31 downto 0);
	signal C     : std_logic_vector(31 downto 0);
	signal D     : std_logic_vector(31 downto 0);
	signal E     : std_logic_vector(31 downto 0);
	signal F     : std_logic_vector(31 downto 0);
	signal G     : std_logic_vector(1 downto 0);
	signal output	: std_logic_vector(15 downto 0);
component Adder_type
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
end component;
component  ADDM4K3S8RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S9RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S12RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S13RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S10RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S11RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S14RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S15RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S2RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S3RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S4RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S5RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S6RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S7RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S0RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

component  ADDM4K3S1RAM 
    PORT
    (
        clock        : IN STD_LOGIC ;
        address        : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
        q        : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
end component;

        signal cVar1S0S0P068P069P012P008: std_logic_vector(   0 downto 0);
        signal cVar1S1S0P068P069P012P008: std_logic_vector(   0 downto 0);
        signal cVar1S2S0P068N069P065P012: std_logic_vector(   0 downto 0);
        signal cVar1S3S0P068N069N065P055: std_logic_vector(   0 downto 0);
        signal cVar1S4S0P068N069N065P055: std_logic_vector(   0 downto 0);
        signal cVar1S5S0P068N069N065N055: std_logic_vector(   0 downto 0);
        signal cVar1S6S0N068P064P063P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S0N068P064N063P035: std_logic_vector(   0 downto 0);
        signal cVar1S8S0N068P064N063P035: std_logic_vector(   0 downto 0);
        signal cVar1S9S0N068P064N063P035: std_logic_vector(   0 downto 0);
        signal cVar1S10S0N068P064N063N035: std_logic_vector(   0 downto 0);
        signal cVar1S11S0N068P064N063N035: std_logic_vector(   0 downto 0);
        signal cVar1S12S0N068N064P067P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S0N068N064P067P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S0N068N064N067P059: std_logic_vector(   0 downto 0);
        signal cVar1S15S0N068N064N067P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S0N068N064N067N059: std_logic_vector(   0 downto 0);
        signal cVar1S17S0N068N064N067N059: std_logic_vector(   0 downto 0);
        signal cVar1S0S1P067P010P068P069: std_logic_vector(   0 downto 0);
        signal cVar1S1S1P067P010P068P069: std_logic_vector(   0 downto 0);
        signal cVar1S2S1P067P010P068N069: std_logic_vector(   0 downto 0);
        signal cVar1S3S1P067P010P068N069: std_logic_vector(   0 downto 0);
        signal cVar1S4S1P067P010P068P012: std_logic_vector(   0 downto 0);
        signal cVar1S5S1P067P010P068N012: std_logic_vector(   0 downto 0);
        signal cVar1S6S1P067P010P068N012: std_logic_vector(   0 downto 0);
        signal cVar1S7S1P067P010P024P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S1P067P010P024N028: std_logic_vector(   0 downto 0);
        signal cVar1S9S1N067P068P014P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S1N067P068P014P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S1N067P068P014P063: std_logic_vector(   0 downto 0);
        signal cVar1S12S1N067P068P014P063: std_logic_vector(   0 downto 0);
        signal cVar1S13S1N067P068P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S14S1N067P068P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S15S1N067P068P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S16S1N067P068P014N066: std_logic_vector(   0 downto 0);
        signal cVar1S17S1N067N068P055P030nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S1N067N068P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S19S1N067N068P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S20S1N067N068P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S21S1N067N068N055P052: std_logic_vector(   0 downto 0);
        signal cVar1S22S1N067N068N055P052: std_logic_vector(   0 downto 0);
        signal cVar1S23S1N067N068N055P052: std_logic_vector(   0 downto 0);
        signal cVar1S24S1N067N068N055N052: std_logic_vector(   0 downto 0);
        signal cVar1S25S1N067N068N055N052: std_logic_vector(   0 downto 0);
        signal cVar1S26S1N067N068N055N052: std_logic_vector(   0 downto 0);
        signal cVar1S0S2P016P047P000P049nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S2P016P047P000N049: std_logic_vector(   0 downto 0);
        signal cVar1S2S2P016P047P000N049: std_logic_vector(   0 downto 0);
        signal cVar1S3S2P016N047P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S2P016N047P052N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S2P016N047N052P060: std_logic_vector(   0 downto 0);
        signal cVar1S6S2P016N047N052P060: std_logic_vector(   0 downto 0);
        signal cVar1S7S2P016N047N052P060: std_logic_vector(   0 downto 0);
        signal cVar1S8S2P016N047N052N060: std_logic_vector(   0 downto 0);
        signal cVar1S9S2P016N047N052N060: std_logic_vector(   0 downto 0);
        signal cVar1S10S2P016N047N052N060: std_logic_vector(   0 downto 0);
        signal cVar1S11S2P016P014P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S12S2P016P014P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S2P016P014P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S14S2P016P014P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S15S2P016P014P063P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S2P016P014N063P060: std_logic_vector(   0 downto 0);
        signal cVar1S17S2P016P014N063P060: std_logic_vector(   0 downto 0);
        signal cVar1S18S2P016P014N063N060: std_logic_vector(   0 downto 0);
        signal cVar1S19S2P016P014N063N060: std_logic_vector(   0 downto 0);
        signal cVar1S20S2P016P014P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S21S2P016P014P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S22S2P016P014P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S23S2P016P014P008P010: std_logic_vector(   0 downto 0);
        signal cVar1S24S2P016P014P008P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S3P047P049P064P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S3P047P049P064P014: std_logic_vector(   0 downto 0);
        signal cVar1S2S3P047P049P064psss: std_logic_vector(   0 downto 0);
        signal cVar1S3S3P047N049P034P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S3N047P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S3N047P052N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S3N047P052N029N027: std_logic_vector(   0 downto 0);
        signal cVar1S7S3N047P052N029N027: std_logic_vector(   0 downto 0);
        signal cVar1S8S3N047P052N029N027: std_logic_vector(   0 downto 0);
        signal cVar1S9S3N047N052P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S10S3N047N052P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S11S3N047N052P060P065: std_logic_vector(   0 downto 0);
        signal cVar1S12S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S16S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S18S3N047N052N060P014: std_logic_vector(   0 downto 0);
        signal cVar1S0S4P014P069P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S4P014P069P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S4P014P069P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S3S4P014P069P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S4S4P014P069P006P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S4P014N069P053P051: std_logic_vector(   0 downto 0);
        signal cVar1S6S4P014N069P053P051: std_logic_vector(   0 downto 0);
        signal cVar1S7S4P014N069P053N051: std_logic_vector(   0 downto 0);
        signal cVar1S8S4P014N069N053P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S4P014N069N053P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S4P014N069N053P045: std_logic_vector(   0 downto 0);
        signal cVar1S11S4P014N069N053N045: std_logic_vector(   0 downto 0);
        signal cVar1S12S4P014N069N053N045: std_logic_vector(   0 downto 0);
        signal cVar1S13S4P014N069N053N045: std_logic_vector(   0 downto 0);
        signal cVar1S14S4P014P024P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S15S4P014P024P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S16S4P014P024P060P010: std_logic_vector(   0 downto 0);
        signal cVar1S17S4P014P024N060P029: std_logic_vector(   0 downto 0);
        signal cVar1S18S4P014P024N060P029: std_logic_vector(   0 downto 0);
        signal cVar1S19S4P014P024N060P029: std_logic_vector(   0 downto 0);
        signal cVar1S20S4P014P024N060N029: std_logic_vector(   0 downto 0);
        signal cVar1S21S4P014P024N060N029: std_logic_vector(   0 downto 0);
        signal cVar1S22S4P014P024N060N029: std_logic_vector(   0 downto 0);
        signal cVar1S23S4P014P024P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S24S4P014P024N047P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S5P053P051P024P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S5P053P051P024N028: std_logic_vector(   0 downto 0);
        signal cVar1S2S5P053P051P024N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S5P053P051P024N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S5P053N051P010P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S5P053N051P010N047: std_logic_vector(   0 downto 0);
        signal cVar1S6S5P053N051P010N047: std_logic_vector(   0 downto 0);
        signal cVar1S7S5P053N051P010N047: std_logic_vector(   0 downto 0);
        signal cVar1S8S5P053N051P010P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S5N053P051P069P010: std_logic_vector(   0 downto 0);
        signal cVar1S10S5N053P051P069P010: std_logic_vector(   0 downto 0);
        signal cVar1S11S5N053P051P069P010: std_logic_vector(   0 downto 0);
        signal cVar1S12S5N053P051P069P010: std_logic_vector(   0 downto 0);
        signal cVar1S13S5N053P051P069P010: std_logic_vector(   0 downto 0);
        signal cVar1S14S5N053P051N069P045: std_logic_vector(   0 downto 0);
        signal cVar1S15S5N053P051N069P045: std_logic_vector(   0 downto 0);
        signal cVar1S16S5N053P051N069N045: std_logic_vector(   0 downto 0);
        signal cVar1S17S5N053P051N069N045: std_logic_vector(   0 downto 0);
        signal cVar1S18S5N053P051N069N045: std_logic_vector(   0 downto 0);
        signal cVar1S19S5N053P051P049P061: std_logic_vector(   0 downto 0);
        signal cVar1S20S5N053P051N049P015: std_logic_vector(   0 downto 0);
        signal cVar1S0S6P047P049P064P012nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S6P047P049P064P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S6P047N049P034P035: std_logic_vector(   0 downto 0);
        signal cVar1S3S6P047N049P034P035: std_logic_vector(   0 downto 0);
        signal cVar1S4S6N047P024P055P030: std_logic_vector(   0 downto 0);
        signal cVar1S5S6N047P024P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S6S6N047P024P055N030: std_logic_vector(   0 downto 0);
        signal cVar1S7S6N047P024N055P053: std_logic_vector(   0 downto 0);
        signal cVar1S8S6N047P024N055P053: std_logic_vector(   0 downto 0);
        signal cVar1S9S6N047P024N055N053: std_logic_vector(   0 downto 0);
        signal cVar1S10S6N047P024P032P045: std_logic_vector(   0 downto 0);
        signal cVar1S11S6N047P024P032N045: std_logic_vector(   0 downto 0);
        signal cVar1S12S6N047P024P032N045: std_logic_vector(   0 downto 0);
        signal cVar1S0S7P053P006P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S7P053P006N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S7P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S3S7P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S4S7P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S7P053P006P063P017: std_logic_vector(   0 downto 0);
        signal cVar1S6S7N053P055P030P057: std_logic_vector(   0 downto 0);
        signal cVar1S7S7N053P055P030P057: std_logic_vector(   0 downto 0);
        signal cVar1S8S7N053P055N030P068: std_logic_vector(   0 downto 0);
        signal cVar1S9S7N053P055N030P068: std_logic_vector(   0 downto 0);
        signal cVar1S10S7N053P055N030P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S7N053N055P047P049nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S7N053N055P047N049: std_logic_vector(   0 downto 0);
        signal cVar1S13S7N053N055P047N049: std_logic_vector(   0 downto 0);
        signal cVar1S14S7N053N055N047P033: std_logic_vector(   0 downto 0);
        signal cVar1S15S7N053N055N047P033: std_logic_vector(   0 downto 0);
        signal cVar1S16S7N053N055N047P033: std_logic_vector(   0 downto 0);
        signal cVar1S17S7N053N055N047N033: std_logic_vector(   0 downto 0);
        signal cVar1S18S7N053N055N047N033: std_logic_vector(   0 downto 0);
        signal cVar1S19S7N053N055N047N033: std_logic_vector(   0 downto 0);
        signal cVar1S0S8P036P053P000P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S8P036P053P000N028: std_logic_vector(   0 downto 0);
        signal cVar1S2S8P036P053P000N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S8P036P053P000N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S8P036N053P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S8P036N053P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S6S8P036N053P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S7S8P036N053P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S8S8P036N053N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S9S8P036N053N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S10S8P036N053N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S11S8P036N053N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S12S8P036N053N046P051: std_logic_vector(   0 downto 0);
        signal cVar1S13S8P036P010P016P008: std_logic_vector(   0 downto 0);
        signal cVar1S14S8P036P010P016P008: std_logic_vector(   0 downto 0);
        signal cVar1S15S8P036P010N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S16S8P036P010N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S8P036P010N016P018: std_logic_vector(   0 downto 0);
        signal cVar1S18S8P036P010N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S19S8P036P010N016N018: std_logic_vector(   0 downto 0);
        signal cVar1S20S8P036P010P024P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S9P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S9P052N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S9P052N029N027P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S9P052N029N027N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S9P052N029N027N028: std_logic_vector(   0 downto 0);
        signal cVar1S5S9N052P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S9N052P046N025P014: std_logic_vector(   0 downto 0);
        signal cVar1S7S9N052P046N025P014: std_logic_vector(   0 downto 0);
        signal cVar1S8S9N052P046N025P014: std_logic_vector(   0 downto 0);
        signal cVar1S9S9N052N046P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S10S9N052N046P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S11S9N052N046P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S12S9N052N046P041N039: std_logic_vector(   0 downto 0);
        signal cVar1S13S9N052N046N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S14S9N052N046N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S9N052N046N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S9N052N046N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S9N052N046N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S0S10P012P053P063P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S10P012P053P063N028: std_logic_vector(   0 downto 0);
        signal cVar1S2S10P012P053P063N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S10P012P053P063N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S10P012P053P063P062: std_logic_vector(   0 downto 0);
        signal cVar1S5S10P012N053P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S6S10P012N053P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S7S10P012N053P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S8S10P012N053P041N039: std_logic_vector(   0 downto 0);
        signal cVar1S9S10P012N053N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S10S10P012N053N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S11S10P012N053N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S12S10P012N053N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S13S10P012P030P006P014: std_logic_vector(   0 downto 0);
        signal cVar1S14S10P012P030P006P014: std_logic_vector(   0 downto 0);
        signal cVar1S15S10P012P030P006P014: std_logic_vector(   0 downto 0);
        signal cVar1S16S10P012P030P006P014: std_logic_vector(   0 downto 0);
        signal cVar1S17S10P012N030P008P031: std_logic_vector(   0 downto 0);
        signal cVar1S18S10P012N030P008P031: std_logic_vector(   0 downto 0);
        signal cVar1S19S10P012N030P008P031: std_logic_vector(   0 downto 0);
        signal cVar1S20S10P012N030P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S21S10P012N030P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S22S10P012N030P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S23S10P012N030P008P011: std_logic_vector(   0 downto 0);
        signal cVar1S0S11P053P006P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S11P053P006N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S11P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S3S11P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S4S11P053P006N028N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S11P053P006P063P017: std_logic_vector(   0 downto 0);
        signal cVar1S6S11N053P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S11N053P041N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S11N053P041N020N021: std_logic_vector(   0 downto 0);
        signal cVar1S9S11N053N041P039P046: std_logic_vector(   0 downto 0);
        signal cVar1S10S11N053N041P039P046: std_logic_vector(   0 downto 0);
        signal cVar1S11S11N053N041P039P046: std_logic_vector(   0 downto 0);
        signal cVar1S12S11N053N041P039N046: std_logic_vector(   0 downto 0);
        signal cVar1S13S11N053N041P039N046: std_logic_vector(   0 downto 0);
        signal cVar1S14S11N053N041P039N046: std_logic_vector(   0 downto 0);
        signal cVar1S15S11N053N041P039N046: std_logic_vector(   0 downto 0);
        signal cVar1S16S11N053N041P039P008: std_logic_vector(   0 downto 0);
        signal cVar1S0S12P015P016P037P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S12P015P016P037P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S12P015P016P037P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S12P015P016N037P063: std_logic_vector(   0 downto 0);
        signal cVar1S4S12P015P016N037P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S12P015P016N037N063: std_logic_vector(   0 downto 0);
        signal cVar1S6S12P015P016N037N063: std_logic_vector(   0 downto 0);
        signal cVar1S7S12P015N016P065P041: std_logic_vector(   0 downto 0);
        signal cVar1S8S12P015N016P065P041: std_logic_vector(   0 downto 0);
        signal cVar1S9S12P015N016P065N041: std_logic_vector(   0 downto 0);
        signal cVar1S10S12P015N016P065N041: std_logic_vector(   0 downto 0);
        signal cVar1S11S12P015N016P065N041: std_logic_vector(   0 downto 0);
        signal cVar1S12S12P015N016P065P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S12P015N016P065P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S12P015N016P065P004: std_logic_vector(   0 downto 0);
        signal cVar1S15S12P015P016P033P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S12P015P016P033P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S12P015P016N033P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S12P015P016N033P035: std_logic_vector(   0 downto 0);
        signal cVar1S19S12P015P016N033N035: std_logic_vector(   0 downto 0);
        signal cVar1S20S12P015P016N033N035: std_logic_vector(   0 downto 0);
        signal cVar1S21S12P015P016P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S12P015P016P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S12P015P016P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S0S13P001P066P011P068: std_logic_vector(   0 downto 0);
        signal cVar1S1S13P001P066P011P068: std_logic_vector(   0 downto 0);
        signal cVar1S2S13P001P066P011P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S13P001P066P011N068: std_logic_vector(   0 downto 0);
        signal cVar1S4S13P001P066P011P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S13P001P066P011P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S13P001P066P011P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S13P001N066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S8S13P001N066P027P009: std_logic_vector(   0 downto 0);
        signal cVar1S9S13P001N066P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S10S13P001N066P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S11S13P001N066N027P053: std_logic_vector(   0 downto 0);
        signal cVar1S12S13P001N066N027P053: std_logic_vector(   0 downto 0);
        signal cVar1S13S13P001N066N027P053: std_logic_vector(   0 downto 0);
        signal cVar1S14S13P001N066N027N053: std_logic_vector(   0 downto 0);
        signal cVar1S15S13P001N066N027N053: std_logic_vector(   0 downto 0);
        signal cVar1S16S13P001N066N027N053: std_logic_vector(   0 downto 0);
        signal cVar1S17S13P001N066N027N053: std_logic_vector(   0 downto 0);
        signal cVar1S18S13P001P006P051P004: std_logic_vector(   0 downto 0);
        signal cVar1S19S13P001P006P051P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S14P015P016P034P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S14P015P016P034N063: std_logic_vector(   0 downto 0);
        signal cVar1S2S14P015P016N034P037: std_logic_vector(   0 downto 0);
        signal cVar1S3S14P015P016N034P037: std_logic_vector(   0 downto 0);
        signal cVar1S4S14P015P016N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S5S14P015P016N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S6S14P015P016N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S7S14P015N016P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S14P015N016P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S9S14P015N016P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S10S14P015N016N046P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S14P015N016N046P022: std_logic_vector(   0 downto 0);
        signal cVar1S12S14P015N016N046P022: std_logic_vector(   0 downto 0);
        signal cVar1S13S14P015N016N046N022: std_logic_vector(   0 downto 0);
        signal cVar1S14S14P015N016N046N022: std_logic_vector(   0 downto 0);
        signal cVar1S15S14P015N016N046N022: std_logic_vector(   0 downto 0);
        signal cVar1S16S14P015N016N046N022: std_logic_vector(   0 downto 0);
        signal cVar1S17S14P015P009P016P033: std_logic_vector(   0 downto 0);
        signal cVar1S18S14P015P009P016P033: std_logic_vector(   0 downto 0);
        signal cVar1S19S14P015P009P016N033: std_logic_vector(   0 downto 0);
        signal cVar1S20S14P015P009P016N033: std_logic_vector(   0 downto 0);
        signal cVar1S21S14P015P009P016P019: std_logic_vector(   0 downto 0);
        signal cVar1S22S14P015P009P016P019: std_logic_vector(   0 downto 0);
        signal cVar1S23S14P015P009P016P019: std_logic_vector(   0 downto 0);
        signal cVar1S24S14P015P009P016P019: std_logic_vector(   0 downto 0);
        signal cVar1S25S14P015P009P016P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S14P015P009P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S15P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S15P046N025P032P014: std_logic_vector(   0 downto 0);
        signal cVar1S2S15P046N025P032P014: std_logic_vector(   0 downto 0);
        signal cVar1S3S15P046N025P032P014: std_logic_vector(   0 downto 0);
        signal cVar1S4S15P046N025P032P014: std_logic_vector(   0 downto 0);
        signal cVar1S5S15N046P016P018P034: std_logic_vector(   0 downto 0);
        signal cVar1S6S15N046P016P018P034: std_logic_vector(   0 downto 0);
        signal cVar1S7S15N046P016P018N034: std_logic_vector(   0 downto 0);
        signal cVar1S8S15N046P016P018N034: std_logic_vector(   0 downto 0);
        signal cVar1S9S15N046P016P018N034: std_logic_vector(   0 downto 0);
        signal cVar1S10S15N046P016P018P019: std_logic_vector(   0 downto 0);
        signal cVar1S11S15N046P016P018P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S15N046P016P018P019: std_logic_vector(   0 downto 0);
        signal cVar1S13S15N046N016P056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S15N046N016P056N057: std_logic_vector(   0 downto 0);
        signal cVar1S15S15N046N016P056N057: std_logic_vector(   0 downto 0);
        signal cVar1S16S15N046N016N056P054: std_logic_vector(   0 downto 0);
        signal cVar1S17S15N046N016N056P054: std_logic_vector(   0 downto 0);
        signal cVar1S18S15N046N016N056P054: std_logic_vector(   0 downto 0);
        signal cVar1S19S15N046N016N056P054: std_logic_vector(   0 downto 0);
        signal cVar1S0S16P016P000P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S16P016P000P023N042: std_logic_vector(   0 downto 0);
        signal cVar1S2S16P016P000N023P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S16P016P000N023P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S16P016P000N023N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S16P016P000N023N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S16P016P000P053P062: std_logic_vector(   0 downto 0);
        signal cVar1S7S16P016P015P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S16P016P015P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S16P016P015P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S16P016P015P034N063: std_logic_vector(   0 downto 0);
        signal cVar1S11S16P016P015N034P037: std_logic_vector(   0 downto 0);
        signal cVar1S12S16P016P015N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S13S16P016P015N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S14S16P016P015N034N037: std_logic_vector(   0 downto 0);
        signal cVar1S15S16P016P015P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S16S16P016P015P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S17S16P016P015P006P019: std_logic_vector(   0 downto 0);
        signal cVar1S18S16P016P015P006P011: std_logic_vector(   0 downto 0);
        signal cVar1S0S17P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S17P023N042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S17P023N042N005P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S17N023P005P053P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S17N023P005P053P006: std_logic_vector(   0 downto 0);
        signal cVar1S5S17N023P005P053P006: std_logic_vector(   0 downto 0);
        signal cVar1S6S17N023P005N053P058: std_logic_vector(   0 downto 0);
        signal cVar1S7S17N023P005N053P058: std_logic_vector(   0 downto 0);
        signal cVar1S8S17N023P005N053P058: std_logic_vector(   0 downto 0);
        signal cVar1S9S17N023P005N053N058: std_logic_vector(   0 downto 0);
        signal cVar1S10S17N023P005N053N058: std_logic_vector(   0 downto 0);
        signal cVar1S11S17N023P005N053N058: std_logic_vector(   0 downto 0);
        signal cVar1S12S17N023P005N053N058: std_logic_vector(   0 downto 0);
        signal cVar1S13S17N023P005P006P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S17N023P005P006N041: std_logic_vector(   0 downto 0);
        signal cVar1S15S17N023P005P006N041: std_logic_vector(   0 downto 0);
        signal cVar1S0S18P011P058P039P024: std_logic_vector(   0 downto 0);
        signal cVar1S1S18P011P058P039P024: std_logic_vector(   0 downto 0);
        signal cVar1S2S18P011P058P039P024: std_logic_vector(   0 downto 0);
        signal cVar1S3S18P011P058P039P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S18P011N058P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S18P011N058P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S6S18P011N058P046N025: std_logic_vector(   0 downto 0);
        signal cVar1S7S18P011N058N046P021: std_logic_vector(   0 downto 0);
        signal cVar1S8S18P011N058N046P021: std_logic_vector(   0 downto 0);
        signal cVar1S9S18P011N058N046N021: std_logic_vector(   0 downto 0);
        signal cVar1S10S18P011N058N046N021: std_logic_vector(   0 downto 0);
        signal cVar1S11S18P011N058N046N021: std_logic_vector(   0 downto 0);
        signal cVar1S12S18P011P029P066P054nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S18P011P029P066N054: std_logic_vector(   0 downto 0);
        signal cVar1S14S18P011P029P066N054: std_logic_vector(   0 downto 0);
        signal cVar1S15S18P011P029P066N054: std_logic_vector(   0 downto 0);
        signal cVar1S16S18P011N029P013P032: std_logic_vector(   0 downto 0);
        signal cVar1S17S18P011N029P013P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S18P011N029P013P032: std_logic_vector(   0 downto 0);
        signal cVar1S19S18P011N029P013P032: std_logic_vector(   0 downto 0);
        signal cVar1S0S19P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S19P021N040P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S19P021N040N041P056: std_logic_vector(   0 downto 0);
        signal cVar1S3S19P021N040N041P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S19N021P001P058P039: std_logic_vector(   0 downto 0);
        signal cVar1S5S19N021P001P058P039: std_logic_vector(   0 downto 0);
        signal cVar1S6S19N021P001N058P020: std_logic_vector(   0 downto 0);
        signal cVar1S7S19N021P001N058P020: std_logic_vector(   0 downto 0);
        signal cVar1S8S19N021P001N058P020: std_logic_vector(   0 downto 0);
        signal cVar1S9S19N021P001N058N020: std_logic_vector(   0 downto 0);
        signal cVar1S10S19N021P001P051P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S20P032P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S20P032P023N042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S20P032P023N042N005: std_logic_vector(   0 downto 0);
        signal cVar1S3S20P032N023P005P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S20P032N023P005N056: std_logic_vector(   0 downto 0);
        signal cVar1S5S20P032N023P005N056: std_logic_vector(   0 downto 0);
        signal cVar1S6S20P032N023P005N056: std_logic_vector(   0 downto 0);
        signal cVar1S7S20P032N023P005P031: std_logic_vector(   0 downto 0);
        signal cVar1S8S20P032N023P005P031: std_logic_vector(   0 downto 0);
        signal cVar1S9S20P032P008P014P051: std_logic_vector(   0 downto 0);
        signal cVar1S10S20P032P008P014P051: std_logic_vector(   0 downto 0);
        signal cVar1S11S20P032P008N014P012: std_logic_vector(   0 downto 0);
        signal cVar1S12S20P032P008N014P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S20P032P008N014N012: std_logic_vector(   0 downto 0);
        signal cVar1S14S20P032P008N014N012: std_logic_vector(   0 downto 0);
        signal cVar1S15S20P032P008P006P068: std_logic_vector(   0 downto 0);
        signal cVar1S0S21P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S21P023N042P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S21P023N042P024N005: std_logic_vector(   0 downto 0);
        signal cVar1S3S21N023P001P047P024: std_logic_vector(   0 downto 0);
        signal cVar1S4S21N023P001P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S5S21N023P001P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S6S21N023P001P047N024: std_logic_vector(   0 downto 0);
        signal cVar1S7S21N023P001N047P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S21N023P001N047P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S21N023P001N047P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S21N023P001P006P028: std_logic_vector(   0 downto 0);
        signal cVar1S0S22P001P010P028P027: std_logic_vector(   0 downto 0);
        signal cVar1S1S22P001P010P028P027: std_logic_vector(   0 downto 0);
        signal cVar1S2S22P001P010P028N027: std_logic_vector(   0 downto 0);
        signal cVar1S3S22P001P010P028N027: std_logic_vector(   0 downto 0);
        signal cVar1S4S22P001P010P028N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S22P001P010P028P000: std_logic_vector(   0 downto 0);
        signal cVar1S6S22P001P010P028P000: std_logic_vector(   0 downto 0);
        signal cVar1S7S22P001P010P028P034nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S22P001P010N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S22P001P010N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S22P001P010N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S11S22P001P004P051P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S22P001P004P051P024: std_logic_vector(   0 downto 0);
        signal cVar1S0S23P027P000P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S23P027P000N048P035: std_logic_vector(   0 downto 0);
        signal cVar1S2S23P027P000N048P035: std_logic_vector(   0 downto 0);
        signal cVar1S3S23N027P009P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S23N027P009P023N042: std_logic_vector(   0 downto 0);
        signal cVar1S5S23N027P009P023N042: std_logic_vector(   0 downto 0);
        signal cVar1S6S23N027P009N023P035: std_logic_vector(   0 downto 0);
        signal cVar1S7S23N027P009N023P035: std_logic_vector(   0 downto 0);
        signal cVar1S8S23N027P009N023N035: std_logic_vector(   0 downto 0);
        signal cVar1S9S23N027P009N023N035: std_logic_vector(   0 downto 0);
        signal cVar1S10S23N027P009N023N035: std_logic_vector(   0 downto 0);
        signal cVar1S11S23N027P009P068P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S23N027P009P068P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S23N027P009P068P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S23N027P009P068P002: std_logic_vector(   0 downto 0);
        signal cVar1S0S24P008P026P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S1S24P008P026P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S2S24P008P026P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S3S24P008P026P055N057: std_logic_vector(   0 downto 0);
        signal cVar1S4S24P008P026P055N057: std_logic_vector(   0 downto 0);
        signal cVar1S5S24P008P026N055P041: std_logic_vector(   0 downto 0);
        signal cVar1S6S24P008P026N055P041: std_logic_vector(   0 downto 0);
        signal cVar1S7S24P008P026N055P041: std_logic_vector(   0 downto 0);
        signal cVar1S8S24P008P026N055N041: std_logic_vector(   0 downto 0);
        signal cVar1S9S24P008P026P045P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S24P008P026P045N047: std_logic_vector(   0 downto 0);
        signal cVar1S11S24P008P026P004P051nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S24P008P026P004N051: std_logic_vector(   0 downto 0);
        signal cVar1S13S24P008P026P004N051: std_logic_vector(   0 downto 0);
        signal cVar1S14S24P008N026P032P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S24P008N026P032P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S24P008N026P032P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S24P008N026P032P039: std_logic_vector(   0 downto 0);
        signal cVar1S0S25P055P026P030P057: std_logic_vector(   0 downto 0);
        signal cVar1S1S25P055P026P030P057: std_logic_vector(   0 downto 0);
        signal cVar1S2S25P055P026N030P031: std_logic_vector(   0 downto 0);
        signal cVar1S3S25P055P026N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S4S25P055P026N030N031: std_logic_vector(   0 downto 0);
        signal cVar1S5S25N055P057P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S25N055P057P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S7S25N055P057P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S8S25N055P057N041P053: std_logic_vector(   0 downto 0);
        signal cVar1S9S25N055P057N041P053: std_logic_vector(   0 downto 0);
        signal cVar1S10S25N055P057N041P053: std_logic_vector(   0 downto 0);
        signal cVar1S11S25N055P057N041N053: std_logic_vector(   0 downto 0);
        signal cVar1S12S25N055P057N041N053: std_logic_vector(   0 downto 0);
        signal cVar1S13S25N055P057P053P037: std_logic_vector(   0 downto 0);
        signal cVar1S0S26P017P019P037P002: std_logic_vector(   0 downto 0);
        signal cVar1S1S26P017P019P037P002: std_logic_vector(   0 downto 0);
        signal cVar1S2S26P017P019P037P002: std_logic_vector(   0 downto 0);
        signal cVar1S3S26P017P019P037P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S26P017P019P037P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S26P017P019N037P018: std_logic_vector(   0 downto 0);
        signal cVar1S6S26P017P019N037P018: std_logic_vector(   0 downto 0);
        signal cVar1S7S26P017P019N037P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S26P017P019N037P018: std_logic_vector(   0 downto 0);
        signal cVar1S9S26P017P019N037P018: std_logic_vector(   0 downto 0);
        signal cVar1S10S26P017N019P037P064nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S26P017N019P037P064: std_logic_vector(   0 downto 0);
        signal cVar1S12S26P017N019P037P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S26P017N019P037P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S26P017N019P037P003: std_logic_vector(   0 downto 0);
        signal cVar1S15S26P017N019P037P003: std_logic_vector(   0 downto 0);
        signal cVar1S16S26P017N019P037P003: std_logic_vector(   0 downto 0);
        signal cVar1S17S26P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S18S26P017P037P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S19S26P017P037P019N064: std_logic_vector(   0 downto 0);
        signal cVar1S20S26P017P037P019P013: std_logic_vector(   0 downto 0);
        signal cVar1S21S26P017P037P019P013: std_logic_vector(   0 downto 0);
        signal cVar1S22S26P017P037P019P013: std_logic_vector(   0 downto 0);
        signal cVar1S23S26P017P037P019P013: std_logic_vector(   0 downto 0);
        signal cVar1S24S26P017P037P019P013: std_logic_vector(   0 downto 0);
        signal cVar1S25S26P017N037P035P019: std_logic_vector(   0 downto 0);
        signal cVar1S26S26P017N037P035P019: std_logic_vector(   0 downto 0);
        signal cVar1S27S26P017N037P035P019: std_logic_vector(   0 downto 0);
        signal cVar1S28S26P017N037P035P019: std_logic_vector(   0 downto 0);
        signal cVar1S29S26P017N037N035P064: std_logic_vector(   0 downto 0);
        signal cVar1S30S26P017N037N035P064: std_logic_vector(   0 downto 0);
        signal cVar1S31S26P017N037N035P064: std_logic_vector(   0 downto 0);
        signal cVar1S0S27P017P051P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S1S27P017P051P048P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S27P017P051P058P041: std_logic_vector(   0 downto 0);
        signal cVar1S3S27P017P051P058P041: std_logic_vector(   0 downto 0);
        signal cVar1S4S27P017P051P058P041: std_logic_vector(   0 downto 0);
        signal cVar1S5S27N017P019P067P024: std_logic_vector(   0 downto 0);
        signal cVar1S6S27N017P019P067P024: std_logic_vector(   0 downto 0);
        signal cVar1S7S27N017P019N067P037: std_logic_vector(   0 downto 0);
        signal cVar1S8S27N017P019N067P037: std_logic_vector(   0 downto 0);
        signal cVar1S9S27N017P019N067P037: std_logic_vector(   0 downto 0);
        signal cVar1S10S27N017P019N067P037: std_logic_vector(   0 downto 0);
        signal cVar1S11S27N017P019N067N037: std_logic_vector(   0 downto 0);
        signal cVar1S12S27N017N019P068P027: std_logic_vector(   0 downto 0);
        signal cVar1S13S27N017N019P068P027: std_logic_vector(   0 downto 0);
        signal cVar1S14S27N017N019P068P027: std_logic_vector(   0 downto 0);
        signal cVar1S15S27N017N019P068N027: std_logic_vector(   0 downto 0);
        signal cVar1S16S27N017N019P068N027: std_logic_vector(   0 downto 0);
        signal cVar1S17S27N017N019P068N027: std_logic_vector(   0 downto 0);
        signal cVar1S18S27N017N019P068N027: std_logic_vector(   0 downto 0);
        signal cVar1S19S27N017N019P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S20S27N017N019P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S0S28P017P068P064P044: std_logic_vector(   0 downto 0);
        signal cVar1S1S28P017P068P064P044: std_logic_vector(   0 downto 0);
        signal cVar1S2S28P017P068P064P044: std_logic_vector(   0 downto 0);
        signal cVar1S3S28P017P068P064N044: std_logic_vector(   0 downto 0);
        signal cVar1S4S28P017P068P064N044: std_logic_vector(   0 downto 0);
        signal cVar1S5S28P017P068P064P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S28P017P068P064N055: std_logic_vector(   0 downto 0);
        signal cVar1S7S28P017P068P064N055: std_logic_vector(   0 downto 0);
        signal cVar1S8S28P017P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S9S28P017P068P019P064: std_logic_vector(   0 downto 0);
        signal cVar1S10S28P017P068P019N064: std_logic_vector(   0 downto 0);
        signal cVar1S11S28P017P068N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S12S28P017P068N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S13S28P017P068N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S28P017P019P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S28P017P019P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S28P017P019P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S28P017P019P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S18S28P017P019N016P010: std_logic_vector(   0 downto 0);
        signal cVar1S19S28P017P019N016N010: std_logic_vector(   0 downto 0);
        signal cVar1S20S28P017P019N016N010: std_logic_vector(   0 downto 0);
        signal cVar1S21S28P017P019N016N010: std_logic_vector(   0 downto 0);
        signal cVar1S22S28P017P019P064P057: std_logic_vector(   0 downto 0);
        signal cVar1S23S28P017P019P064P057: std_logic_vector(   0 downto 0);
        signal cVar1S24S28P017P019P064P068: std_logic_vector(   0 downto 0);
        signal cVar1S25S28P017P019P064P068: std_logic_vector(   0 downto 0);
        signal cVar1S26S28P017P019P064N068: std_logic_vector(   0 downto 0);
        signal cVar1S27S28P017P019P064N068: std_logic_vector(   0 downto 0);
        signal cVar1S0S29P017P013P011P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S29P017P013P011P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S29P017P013N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S3S29P017P013N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S4S29P017P013N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S5S29P017P013N011P029: std_logic_vector(   0 downto 0);
        signal cVar1S6S29P017P013P067P027: std_logic_vector(   0 downto 0);
        signal cVar1S7S29P017P013P067P051: std_logic_vector(   0 downto 0);
        signal cVar1S8S29N017P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S29N017P044N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S29N017P044N023N025: std_logic_vector(   0 downto 0);
        signal cVar1S11S29N017N044P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S12S29N017N044P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S13S29N017N044P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S14S29N017N044P055P057: std_logic_vector(   0 downto 0);
        signal cVar1S15S29N017N044P055N057: std_logic_vector(   0 downto 0);
        signal cVar1S16S29N017N044N055P041: std_logic_vector(   0 downto 0);
        signal cVar1S17S29N017N044N055P041: std_logic_vector(   0 downto 0);
        signal cVar1S18S29N017N044N055N041: std_logic_vector(   0 downto 0);
        signal cVar1S19S29N017N044N055N041: std_logic_vector(   0 downto 0);
        signal cVar1S0S30P017P036P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S30P017P036P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S30P017P036P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S30P017P036N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S4S30P017P036N044P041: std_logic_vector(   0 downto 0);
        signal cVar1S5S30P017P036N044N041: std_logic_vector(   0 downto 0);
        signal cVar1S6S30P017P036N044N041: std_logic_vector(   0 downto 0);
        signal cVar1S7S30P017P036N044N041: std_logic_vector(   0 downto 0);
        signal cVar1S8S30P017P036P004P013: std_logic_vector(   0 downto 0);
        signal cVar1S9S30P017P036P004P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S30P017P036P004N013: std_logic_vector(   0 downto 0);
        signal cVar1S11S30P017P036P004N013: std_logic_vector(   0 downto 0);
        signal cVar1S12S30P017P036P004P006: std_logic_vector(   0 downto 0);
        signal cVar1S13S30P017P044P063P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S30P017P044P063P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S30P017P044N063P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S30P017P044N063P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S30P017P044N063P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S30P017P044N063P065: std_logic_vector(   0 downto 0);
        signal cVar1S19S30P017P044P034P014: std_logic_vector(   0 downto 0);
        signal cVar1S0S31P033P054P061P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S31P033P054N061P063: std_logic_vector(   0 downto 0);
        signal cVar1S2S31P033P054N061P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S31N033P061P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S31N033P061P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S5S31N033P061P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S6S31N033P061P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S7S31N033P061N029P040: std_logic_vector(   0 downto 0);
        signal cVar1S8S31N033P061N029P040: std_logic_vector(   0 downto 0);
        signal cVar1S9S31N033P061N029P040: std_logic_vector(   0 downto 0);
        signal cVar1S10S31N033P061N029N040: std_logic_vector(   0 downto 0);
        signal cVar1S11S31N033P061N029N040: std_logic_vector(   0 downto 0);
        signal cVar1S12S31N033P061P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S13S31N033P061P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S31N033P061P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S31N033P061P059P032: std_logic_vector(   0 downto 0);
        signal cVar1S16S31N033P061N059P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S31N033P061N059N018: std_logic_vector(   0 downto 0);
        signal cVar1S0S32P061P033P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S1S32P061P033P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S2S32P061P033P060P064: std_logic_vector(   0 downto 0);
        signal cVar1S3S32P061P033P060N064: std_logic_vector(   0 downto 0);
        signal cVar1S4S32P061P033P060N064: std_logic_vector(   0 downto 0);
        signal cVar1S5S32P061P033P060P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S32P061P033P060N032: std_logic_vector(   0 downto 0);
        signal cVar1S7S32P061P033P060N032: std_logic_vector(   0 downto 0);
        signal cVar1S8S32P061P033P065P060: std_logic_vector(   0 downto 0);
        signal cVar1S9S32P061P033P065P060: std_logic_vector(   0 downto 0);
        signal cVar1S10S32P061P033P065N060: std_logic_vector(   0 downto 0);
        signal cVar1S11S32P061P033P065P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S32P061P059P032P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S32P061P059P032P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S32P061P059P032P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S32P061P059P032P064: std_logic_vector(   0 downto 0);
        signal cVar1S16S32P061P059P032P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S32P061P059P032N067: std_logic_vector(   0 downto 0);
        signal cVar1S18S32P061P059P032N067: std_logic_vector(   0 downto 0);
        signal cVar1S19S32P061N059P018P034: std_logic_vector(   0 downto 0);
        signal cVar1S20S32P061N059P018P034: std_logic_vector(   0 downto 0);
        signal cVar1S21S32P061N059N018P063: std_logic_vector(   0 downto 0);
        signal cVar1S0S33P062P013P054P037: std_logic_vector(   0 downto 0);
        signal cVar1S1S33P062P013P054N037: std_logic_vector(   0 downto 0);
        signal cVar1S2S33P062P013P054N037: std_logic_vector(   0 downto 0);
        signal cVar1S3S33P062P013P054P068: std_logic_vector(   0 downto 0);
        signal cVar1S4S33P062P013P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S5S33P062P013P067P059: std_logic_vector(   0 downto 0);
        signal cVar1S6S33P062P013P067P011: std_logic_vector(   0 downto 0);
        signal cVar1S7S33N062P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S33N062P041N020P035: std_logic_vector(   0 downto 0);
        signal cVar1S9S33N062P041N020P035: std_logic_vector(   0 downto 0);
        signal cVar1S10S33N062N041P033P061: std_logic_vector(   0 downto 0);
        signal cVar1S11S33N062N041P033P061: std_logic_vector(   0 downto 0);
        signal cVar1S12S33N062N041P033N061: std_logic_vector(   0 downto 0);
        signal cVar1S13S33N062N041P033N061: std_logic_vector(   0 downto 0);
        signal cVar1S14S33N062N041P033N061: std_logic_vector(   0 downto 0);
        signal cVar1S15S33N062N041N033P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S33N062N041N033P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S33N062N041N033P039: std_logic_vector(   0 downto 0);
        signal cVar1S18S33N062N041N033P039: std_logic_vector(   0 downto 0);
        signal cVar1S0S34P011P029P062P003: std_logic_vector(   0 downto 0);
        signal cVar1S1S34P011P029P062P003: std_logic_vector(   0 downto 0);
        signal cVar1S2S34P011P029P062P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S34P011P029N062P059: std_logic_vector(   0 downto 0);
        signal cVar1S4S34P011P029N062P059: std_logic_vector(   0 downto 0);
        signal cVar1S5S34P011P029N062P059: std_logic_vector(   0 downto 0);
        signal cVar1S6S34P011P029N062N059: std_logic_vector(   0 downto 0);
        signal cVar1S7S34P011P029N062N059: std_logic_vector(   0 downto 0);
        signal cVar1S8S34P011P029N062N059: std_logic_vector(   0 downto 0);
        signal cVar1S9S34P011P029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S34P011P029N052P004: std_logic_vector(   0 downto 0);
        signal cVar1S11S34P011P029N052P004: std_logic_vector(   0 downto 0);
        signal cVar1S12S34P011P013P032P029: std_logic_vector(   0 downto 0);
        signal cVar1S13S34P011P013P032N029: std_logic_vector(   0 downto 0);
        signal cVar1S14S34P011P013P032N029: std_logic_vector(   0 downto 0);
        signal cVar1S15S34P011P013P032N029: std_logic_vector(   0 downto 0);
        signal cVar1S16S34P011P013P004P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S34P011P013P004P008: std_logic_vector(   0 downto 0);
        signal cVar1S0S35P015P022P034P054: std_logic_vector(   0 downto 0);
        signal cVar1S1S35P015P022P034P054: std_logic_vector(   0 downto 0);
        signal cVar1S2S35P015P022P034P054: std_logic_vector(   0 downto 0);
        signal cVar1S3S35P015P022P034P054: std_logic_vector(   0 downto 0);
        signal cVar1S4S35P015P022P034P044: std_logic_vector(   0 downto 0);
        signal cVar1S5S35P015P022P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S35N015P064P043P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S35N015P064P043P033: std_logic_vector(   0 downto 0);
        signal cVar1S8S35N015P064P043P033: std_logic_vector(   0 downto 0);
        signal cVar1S9S35N015P064P043P033: std_logic_vector(   0 downto 0);
        signal cVar1S10S35N015N064P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S35N015N064P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S35N015N064P068P034: std_logic_vector(   0 downto 0);
        signal cVar1S13S35N015N064P068N034: std_logic_vector(   0 downto 0);
        signal cVar1S14S35N015N064P068N034: std_logic_vector(   0 downto 0);
        signal cVar1S15S35N015N064P068N034: std_logic_vector(   0 downto 0);
        signal cVar1S16S35N015N064P068N034: std_logic_vector(   0 downto 0);
        signal cVar1S17S35N015N064P068P011: std_logic_vector(   0 downto 0);
        signal cVar1S18S35N015N064P068P011: std_logic_vector(   0 downto 0);
        signal cVar1S19S35N015N064P068P011: std_logic_vector(   0 downto 0);
        signal cVar1S20S35N015N064P068P011: std_logic_vector(   0 downto 0);
        signal cVar1S0S36P011P015P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S1S36P011P015P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S2S36P011P015P065P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S36P011P015P065N063: std_logic_vector(   0 downto 0);
        signal cVar1S4S36P011P015P065N063: std_logic_vector(   0 downto 0);
        signal cVar1S5S36P011P015P065N063: std_logic_vector(   0 downto 0);
        signal cVar1S6S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S7S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S36P011P015N065P063: std_logic_vector(   0 downto 0);
        signal cVar1S12S36P011P015P022P059: std_logic_vector(   0 downto 0);
        signal cVar1S13S36P011P015P022N059: std_logic_vector(   0 downto 0);
        signal cVar1S14S36P011P015P022N059: std_logic_vector(   0 downto 0);
        signal cVar1S15S36P011P015P022N059: std_logic_vector(   0 downto 0);
        signal cVar1S16S36P011P004P029P054nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S36P011P004P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S18S36P011P004P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S19S36P011P004N029P002: std_logic_vector(   0 downto 0);
        signal cVar1S20S36P011P004N029P002: std_logic_vector(   0 downto 0);
        signal cVar1S21S36P011P004P000P056: std_logic_vector(   0 downto 0);
        signal cVar1S0S37P015P031P022P006: std_logic_vector(   0 downto 0);
        signal cVar1S1S37P015P031P022P006: std_logic_vector(   0 downto 0);
        signal cVar1S2S37P015P031P022P006: std_logic_vector(   0 downto 0);
        signal cVar1S3S37P015P031P022P006: std_logic_vector(   0 downto 0);
        signal cVar1S4S37P015P031P022P012nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S37P015P031P004P030: std_logic_vector(   0 downto 0);
        signal cVar1S6S37P015P031P004P030: std_logic_vector(   0 downto 0);
        signal cVar1S7S37N015P065P007P052nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S37N015P065P007N052: std_logic_vector(   0 downto 0);
        signal cVar1S9S37N015P065P007N052: std_logic_vector(   0 downto 0);
        signal cVar1S10S37N015P065P007P009: std_logic_vector(   0 downto 0);
        signal cVar1S11S37N015N065P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S37N015N065P022N043: std_logic_vector(   0 downto 0);
        signal cVar1S13S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S16S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S17S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S18S37N015N065N022P043: std_logic_vector(   0 downto 0);
        signal cVar1S0S38P006P024P015P014: std_logic_vector(   0 downto 0);
        signal cVar1S1S38P006P024P015P014: std_logic_vector(   0 downto 0);
        signal cVar1S2S38P006P024P015P014: std_logic_vector(   0 downto 0);
        signal cVar1S3S38P006P024P015N014: std_logic_vector(   0 downto 0);
        signal cVar1S4S38P006P024P015N014: std_logic_vector(   0 downto 0);
        signal cVar1S5S38P006P024P015N014: std_logic_vector(   0 downto 0);
        signal cVar1S6S38P006P024P015N014: std_logic_vector(   0 downto 0);
        signal cVar1S7S38P006P024P015P053: std_logic_vector(   0 downto 0);
        signal cVar1S8S38P006P024P015N053: std_logic_vector(   0 downto 0);
        signal cVar1S9S38P006P024P015N053: std_logic_vector(   0 downto 0);
        signal cVar1S10S38P006P024P014P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S38P006P024P014N047: std_logic_vector(   0 downto 0);
        signal cVar1S12S38P006P024P014N047: std_logic_vector(   0 downto 0);
        signal cVar1S13S38P006P024P014P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S38P006P034P024P051: std_logic_vector(   0 downto 0);
        signal cVar1S15S38P006P034N024P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S38P006P034N024P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S38P006P034N024P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S38P006P034P036P011: std_logic_vector(   0 downto 0);
        signal cVar1S0S39P006P067P024P043: std_logic_vector(   0 downto 0);
        signal cVar1S1S39P006P067P024P043: std_logic_vector(   0 downto 0);
        signal cVar1S2S39P006P067P024P043: std_logic_vector(   0 downto 0);
        signal cVar1S3S39P006P067P024P043: std_logic_vector(   0 downto 0);
        signal cVar1S4S39P006P067P024P043: std_logic_vector(   0 downto 0);
        signal cVar1S5S39P006P067P024P014: std_logic_vector(   0 downto 0);
        signal cVar1S6S39P006N067P015P045: std_logic_vector(   0 downto 0);
        signal cVar1S7S39P006N067P015P045: std_logic_vector(   0 downto 0);
        signal cVar1S8S39P006N067P015P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S39P006N067P015P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S39P006N067N015P014: std_logic_vector(   0 downto 0);
        signal cVar1S11S39P006N067N015P014: std_logic_vector(   0 downto 0);
        signal cVar1S12S39P006N067N015N014: std_logic_vector(   0 downto 0);
        signal cVar1S13S39P006N067N015N014: std_logic_vector(   0 downto 0);
        signal cVar1S14S39P006P051P024P011: std_logic_vector(   0 downto 0);
        signal cVar1S15S39P006P051P024P011: std_logic_vector(   0 downto 0);
        signal cVar1S16S39P006P051N024P065: std_logic_vector(   0 downto 0);
        signal cVar1S17S39P006P051N024P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S39P006P051P067P014: std_logic_vector(   0 downto 0);
        signal cVar1S0S40P014P032P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S1S40P014P032P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S40P014P032P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S3S40P014P032P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S4S40P014P032P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S5S40P014P032P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S6S40P014P032N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S7S40P014P032N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S8S40P014P032N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S9S40P014P032N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S10S40P014P032N030P057: std_logic_vector(   0 downto 0);
        signal cVar1S11S40P014P032P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S12S40P014P032P010P012: std_logic_vector(   0 downto 0);
        signal cVar1S13S40P014P032P010N012: std_logic_vector(   0 downto 0);
        signal cVar1S14S40P014P032P010N012: std_logic_vector(   0 downto 0);
        signal cVar1S15S40P014P032P010P017: std_logic_vector(   0 downto 0);
        signal cVar1S16S40P014P024P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S17S40P014P024P044P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S40P014P024P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S40P014P024P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S20S40P014P024P044N032: std_logic_vector(   0 downto 0);
        signal cVar1S21S40P014P024P044P062: std_logic_vector(   0 downto 0);
        signal cVar1S22S40P014P024P054P036: std_logic_vector(   0 downto 0);
        signal cVar1S0S41P035P015P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S41P035P015P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S2S41P035P015N027P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S41P035P015N027P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S41P035P015N027N022: std_logic_vector(   0 downto 0);
        signal cVar1S5S41P035P015N027N022: std_logic_vector(   0 downto 0);
        signal cVar1S6S41P035P015N027N022: std_logic_vector(   0 downto 0);
        signal cVar1S7S41P035P015N027N022: std_logic_vector(   0 downto 0);
        signal cVar1S8S41P035P015P026P061: std_logic_vector(   0 downto 0);
        signal cVar1S9S41P035P015P026P061: std_logic_vector(   0 downto 0);
        signal cVar1S10S41P035P015N026P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S41P035P015N026P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S41P035P015N026P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S41P035P015N026P062: std_logic_vector(   0 downto 0);
        signal cVar1S14S41P035P015N026P062: std_logic_vector(   0 downto 0);
        signal cVar1S15S41P035P045P006P063: std_logic_vector(   0 downto 0);
        signal cVar1S16S41P035P045P006P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S41P035P045P006N063: std_logic_vector(   0 downto 0);
        signal cVar1S18S41P035P045P006N063: std_logic_vector(   0 downto 0);
        signal cVar1S19S41P035P045P006P034: std_logic_vector(   0 downto 0);
        signal cVar1S0S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S1S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S2S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S3S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S42P015P035P001P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S42P015P035P001P013: std_logic_vector(   0 downto 0);
        signal cVar1S7S42P015P035P020P045: std_logic_vector(   0 downto 0);
        signal cVar1S8S42P015P035P020P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S42P015P035P020P045: std_logic_vector(   0 downto 0);
        signal cVar1S10S42P015P009P034P055: std_logic_vector(   0 downto 0);
        signal cVar1S11S42P015P009P034P055: std_logic_vector(   0 downto 0);
        signal cVar1S12S42P015P009P034P055: std_logic_vector(   0 downto 0);
        signal cVar1S13S42P015P009P034N055: std_logic_vector(   0 downto 0);
        signal cVar1S14S42P015P009P034N055: std_logic_vector(   0 downto 0);
        signal cVar1S15S42P015P009P034N055: std_logic_vector(   0 downto 0);
        signal cVar1S16S42P015P009P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S17S42P015P009P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S18S42P015P009P034P063: std_logic_vector(   0 downto 0);
        signal cVar1S19S42P015P009P034N063: std_logic_vector(   0 downto 0);
        signal cVar1S20S42P015P009P041P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S43P015P034P022P016: std_logic_vector(   0 downto 0);
        signal cVar1S1S43P015P034P022P016: std_logic_vector(   0 downto 0);
        signal cVar1S2S43P015P034P022P016: std_logic_vector(   0 downto 0);
        signal cVar1S3S43P015P034P022P016: std_logic_vector(   0 downto 0);
        signal cVar1S4S43P015P034P022P016: std_logic_vector(   0 downto 0);
        signal cVar1S5S43P015P034P022P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S43P015P034P043P044: std_logic_vector(   0 downto 0);
        signal cVar1S7S43N015P027P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S43N015P027N048P005: std_logic_vector(   0 downto 0);
        signal cVar1S9S43N015P027N048P005: std_logic_vector(   0 downto 0);
        signal cVar1S10S43N015N027P030P012: std_logic_vector(   0 downto 0);
        signal cVar1S11S43N015N027P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S12S43N015N027P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S13S43N015N027P030N012: std_logic_vector(   0 downto 0);
        signal cVar1S14S43N015N027N030P040: std_logic_vector(   0 downto 0);
        signal cVar1S15S43N015N027N030P040: std_logic_vector(   0 downto 0);
        signal cVar1S16S43N015N027N030P040: std_logic_vector(   0 downto 0);
        signal cVar1S17S43N015N027N030N040: std_logic_vector(   0 downto 0);
        signal cVar1S0S44P015P027P000P048nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S44P015P027P000N048: std_logic_vector(   0 downto 0);
        signal cVar1S2S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S3S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S4S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S5S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S6S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S7S44P015N027P018P068: std_logic_vector(   0 downto 0);
        signal cVar1S8S44P015N027P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S9S44P015N027P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S10S44P015N027P018P013: std_logic_vector(   0 downto 0);
        signal cVar1S11S44P015N027P018N013: std_logic_vector(   0 downto 0);
        signal cVar1S12S44P015N027P018N013: std_logic_vector(   0 downto 0);
        signal cVar1S13S44P015N027P018N013: std_logic_vector(   0 downto 0);
        signal cVar1S14S44P015P051P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S15S44P015P051P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S16S44P015P051P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S17S44P015P051P068P036: std_logic_vector(   0 downto 0);
        signal cVar1S18S44P015P051P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S19S44P015P051P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S20S44P015P051P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S44P015P051P053P000: std_logic_vector(   0 downto 0);
        signal cVar1S22S44P015P051N053P049: std_logic_vector(   0 downto 0);
        signal cVar1S0S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S1S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S2S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S3S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S5S45P015P018P030P056: std_logic_vector(   0 downto 0);
        signal cVar1S6S45P015P018P030P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S45P015P018P030N069: std_logic_vector(   0 downto 0);
        signal cVar1S8S45P015N018P019P017: std_logic_vector(   0 downto 0);
        signal cVar1S9S45P015N018P019P017: std_logic_vector(   0 downto 0);
        signal cVar1S10S45P015N018P019P017: std_logic_vector(   0 downto 0);
        signal cVar1S11S45P015N018P019P017: std_logic_vector(   0 downto 0);
        signal cVar1S12S45P015N018P019P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S45P015N018N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S14S45P015N018N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S15S45P015N018N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S45P015N018N019P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S45P015P051P068P022: std_logic_vector(   0 downto 0);
        signal cVar1S18S45P015P051P068P022: std_logic_vector(   0 downto 0);
        signal cVar1S19S45P015P051P068P018: std_logic_vector(   0 downto 0);
        signal cVar1S20S45P015P051P068N018: std_logic_vector(   0 downto 0);
        signal cVar1S21S45P015P051P053P000: std_logic_vector(   0 downto 0);
        signal cVar1S22S45P015P051N053P049: std_logic_vector(   0 downto 0);
        signal cVar1S0S46P068P019P057P030: std_logic_vector(   0 downto 0);
        signal cVar1S1S46P068P019P057N030: std_logic_vector(   0 downto 0);
        signal cVar1S2S46P068P019P057N030: std_logic_vector(   0 downto 0);
        signal cVar1S3S46P068P019N057P005: std_logic_vector(   0 downto 0);
        signal cVar1S4S46P068P019N057P005: std_logic_vector(   0 downto 0);
        signal cVar1S5S46P068P019N057N005: std_logic_vector(   0 downto 0);
        signal cVar1S6S46P068P019N057N005: std_logic_vector(   0 downto 0);
        signal cVar1S7S46P068P019N057N005: std_logic_vector(   0 downto 0);
        signal cVar1S8S46P068P019N057N005: std_logic_vector(   0 downto 0);
        signal cVar1S9S46P068P019P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S10S46P068P019P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S11S46P068P019P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S12S46P068P019P006P060: std_logic_vector(   0 downto 0);
        signal cVar1S13S46P068P009P064P053: std_logic_vector(   0 downto 0);
        signal cVar1S14S46P068P009P064P053: std_logic_vector(   0 downto 0);
        signal cVar1S15S46P068P009P064P053: std_logic_vector(   0 downto 0);
        signal cVar1S16S46P068P009N064P056: std_logic_vector(   0 downto 0);
        signal cVar1S17S46P068P009N064P056: std_logic_vector(   0 downto 0);
        signal cVar1S18S46P068P009N064N056: std_logic_vector(   0 downto 0);
        signal cVar1S19S46P068P009N064N056: std_logic_vector(   0 downto 0);
        signal cVar1S20S46P068P009P002P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S46P068P009P002P066: std_logic_vector(   0 downto 0);
        signal cVar1S0S47P019P033P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S1S47P019P033P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S2S47P019P033P006P043: std_logic_vector(   0 downto 0);
        signal cVar1S3S47P019P033P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S4S47P019P033P006P010: std_logic_vector(   0 downto 0);
        signal cVar1S5S47P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S6S47P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S47P019P033P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S8S47P019P033P016N067: std_logic_vector(   0 downto 0);
        signal cVar1S9S47N019P057P041P000: std_logic_vector(   0 downto 0);
        signal cVar1S10S47N019P057P041P000: std_logic_vector(   0 downto 0);
        signal cVar1S11S47N019P057P041P000: std_logic_vector(   0 downto 0);
        signal cVar1S12S47N019P057P041P000: std_logic_vector(   0 downto 0);
        signal cVar1S13S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S14S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S15S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S16S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S17S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S18S47N019N057P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S19S47N019N057P069P029: std_logic_vector(   0 downto 0);
        signal cVar1S20S47N019N057P069N029: std_logic_vector(   0 downto 0);
        signal cVar1S21S47N019N057P069N029: std_logic_vector(   0 downto 0);
        signal cVar1S0S48P019P069P061P007: std_logic_vector(   0 downto 0);
        signal cVar1S1S48P019P069P061P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S48P019P069P061P007: std_logic_vector(   0 downto 0);
        signal cVar1S3S48P019P069P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S4S48P019P069P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S5S48P019P069P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S6S48P019P069P061P033: std_logic_vector(   0 downto 0);
        signal cVar1S7S48P019P069P061N033: std_logic_vector(   0 downto 0);
        signal cVar1S8S48P019P069P061N033: std_logic_vector(   0 downto 0);
        signal cVar1S9S48P019P069P045P043: std_logic_vector(   0 downto 0);
        signal cVar1S10S48P019P069P045P043: std_logic_vector(   0 downto 0);
        signal cVar1S11S48P019P059P041P003: std_logic_vector(   0 downto 0);
        signal cVar1S12S48P019N059P061P033: std_logic_vector(   0 downto 0);
        signal cVar1S13S48P019N059P061P033: std_logic_vector(   0 downto 0);
        signal cVar1S14S48P019N059P061P033: std_logic_vector(   0 downto 0);
        signal cVar1S15S48P019N059P061P033: std_logic_vector(   0 downto 0);
        signal cVar1S16S48P019N059P061P018: std_logic_vector(   0 downto 0);
        signal cVar1S17S48P019N059P061P018: std_logic_vector(   0 downto 0);
        signal cVar1S0S49P019P033P057P013: std_logic_vector(   0 downto 0);
        signal cVar1S1S49P019P033P057P013: std_logic_vector(   0 downto 0);
        signal cVar1S2S49P019P033P057P013: std_logic_vector(   0 downto 0);
        signal cVar1S3S49P019P033P057P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S49P019P033P057P030: std_logic_vector(   0 downto 0);
        signal cVar1S5S49P019P033P057N030: std_logic_vector(   0 downto 0);
        signal cVar1S6S49P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S49P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S8S49P019P033P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S49P019P033P016N067: std_logic_vector(   0 downto 0);
        signal cVar1S10S49N019P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S49N019P007N025P059: std_logic_vector(   0 downto 0);
        signal cVar1S12S49N019P007N025P059: std_logic_vector(   0 downto 0);
        signal cVar1S13S49N019N007P060P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S49N019N007P060P004: std_logic_vector(   0 downto 0);
        signal cVar1S15S49N019N007N060P057: std_logic_vector(   0 downto 0);
        signal cVar1S16S49N019N007N060P057: std_logic_vector(   0 downto 0);
        signal cVar1S17S49N019N007N060P057: std_logic_vector(   0 downto 0);
        signal cVar1S18S49N019N007N060P057: std_logic_vector(   0 downto 0);
        signal cVar1S19S49N019N007N060N057: std_logic_vector(   0 downto 0);
        signal cVar1S20S49N019N007N060N057: std_logic_vector(   0 downto 0);
        signal cVar1S0S50P019P014P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S50P019P014P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S2S50P019P014N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S3S50P019P014N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S4S50P019P014N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S5S50P019P014N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S6S50P019P014P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S7S50P019P014P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S8S50P019P014P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S9S50P019P014P030P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S50P019P014P030P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S50P019P002P020P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S50P019P002P020P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S50P019P002P020N013: std_logic_vector(   0 downto 0);
        signal cVar1S14S50P019P002P020N013: std_logic_vector(   0 downto 0);
        signal cVar1S15S50P019P002P020P013: std_logic_vector(   0 downto 0);
        signal cVar1S16S50P019P002P054P009: std_logic_vector(   0 downto 0);
        signal cVar1S17S50P019P002P054P009: std_logic_vector(   0 downto 0);
        signal cVar1S0S51P019P002P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S1S51P019P002P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S2S51P019P002P020P039: std_logic_vector(   0 downto 0);
        signal cVar1S3S51P019P002P020P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S51P019P002P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S5S51P019P002P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S6S51P019P002P054P000: std_logic_vector(   0 downto 0);
        signal cVar1S7S51N019P017P042P015: std_logic_vector(   0 downto 0);
        signal cVar1S8S51N019P017P042P015: std_logic_vector(   0 downto 0);
        signal cVar1S9S51N019P017P042P015: std_logic_vector(   0 downto 0);
        signal cVar1S10S51N019P017P042P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S51N019N017P005P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S51N019N017P005N023: std_logic_vector(   0 downto 0);
        signal cVar1S13S51N019N017P005N023: std_logic_vector(   0 downto 0);
        signal cVar1S14S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S15S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S16S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S17S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S18S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S19S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S20S51N019N017N005P012: std_logic_vector(   0 downto 0);
        signal cVar1S0S52P019P012P030P050: std_logic_vector(   0 downto 0);
        signal cVar1S1S52P019P012P030P050: std_logic_vector(   0 downto 0);
        signal cVar1S2S52P019P012P030N050: std_logic_vector(   0 downto 0);
        signal cVar1S3S52P019P012P030N050: std_logic_vector(   0 downto 0);
        signal cVar1S4S52P019P012P030N050: std_logic_vector(   0 downto 0);
        signal cVar1S5S52P019P012P030N050: std_logic_vector(   0 downto 0);
        signal cVar1S6S52P019P012P030P010: std_logic_vector(   0 downto 0);
        signal cVar1S7S52P019P012P030N010: std_logic_vector(   0 downto 0);
        signal cVar1S8S52P019P012P030N010: std_logic_vector(   0 downto 0);
        signal cVar1S9S52P019P012P008P031: std_logic_vector(   0 downto 0);
        signal cVar1S10S52P019P012P008P031: std_logic_vector(   0 downto 0);
        signal cVar1S11S52P019P012P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S12S52P019P012P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S13S52P019P012P008N031: std_logic_vector(   0 downto 0);
        signal cVar1S14S52P019P012P008P011: std_logic_vector(   0 downto 0);
        signal cVar1S15S52P019P033P049P028: std_logic_vector(   0 downto 0);
        signal cVar1S16S52P019P033P049P028: std_logic_vector(   0 downto 0);
        signal cVar1S17S52P019P033P049P068: std_logic_vector(   0 downto 0);
        signal cVar1S18S52P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S19S52P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S20S52P019P033P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S0S53P019P033P049P048: std_logic_vector(   0 downto 0);
        signal cVar1S1S53P019P033P049P048: std_logic_vector(   0 downto 0);
        signal cVar1S2S53P019P033P049P048: std_logic_vector(   0 downto 0);
        signal cVar1S3S53P019P033P049P048: std_logic_vector(   0 downto 0);
        signal cVar1S4S53P019P033P049P068: std_logic_vector(   0 downto 0);
        signal cVar1S5S53P019P033P049P068: std_logic_vector(   0 downto 0);
        signal cVar1S6S53P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S7S53P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S8S53P019P033P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S9S53N019P050P021P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S53N019P050P021N027: std_logic_vector(   0 downto 0);
        signal cVar1S11S53N019N050P032P008: std_logic_vector(   0 downto 0);
        signal cVar1S12S53N019N050P032P008: std_logic_vector(   0 downto 0);
        signal cVar1S13S53N019N050P032P008: std_logic_vector(   0 downto 0);
        signal cVar1S14S53N019N050N032P023: std_logic_vector(   0 downto 0);
        signal cVar1S15S53N019N050N032P023: std_logic_vector(   0 downto 0);
        signal cVar1S16S53N019N050N032N023: std_logic_vector(   0 downto 0);
        signal cVar1S17S53N019N050N032N023: std_logic_vector(   0 downto 0);
        signal cVar1S0S54P019P015P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S1S54P019P015P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S2S54P019P015P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S3S54P019P015N017P063: std_logic_vector(   0 downto 0);
        signal cVar1S4S54P019P015N017P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S54P019P015N017P063: std_logic_vector(   0 downto 0);
        signal cVar1S6S54P019P015P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S54P019P015P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S8S54P019P015P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S9S54P019P015P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S10S54P019P015P017N061: std_logic_vector(   0 downto 0);
        signal cVar1S11S54P019P015P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S12S54P019P015P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S13S54P019P033P060P017: std_logic_vector(   0 downto 0);
        signal cVar1S14S54P019P033P060P017: std_logic_vector(   0 downto 0);
        signal cVar1S15S54P019P033P060P017: std_logic_vector(   0 downto 0);
        signal cVar1S16S54P019P033P060N017: std_logic_vector(   0 downto 0);
        signal cVar1S17S54P019P033P060N017: std_logic_vector(   0 downto 0);
        signal cVar1S18S54P019P033P060N017: std_logic_vector(   0 downto 0);
        signal cVar1S19S54P019P033P060P009: std_logic_vector(   0 downto 0);
        signal cVar1S20S54P019P033P060P009: std_logic_vector(   0 downto 0);
        signal cVar1S21S54P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S22S54P019P033P016P065: std_logic_vector(   0 downto 0);
        signal cVar1S23S54P019P033P016P067: std_logic_vector(   0 downto 0);
        signal cVar1S24S54P019P033P016N067: std_logic_vector(   0 downto 0);
        signal cVar1S0S55P015P068P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S1S55P015P068P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S2S55P015P068P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S3S55P015P068P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S4S55P015P068P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S5S55P015P068P051P053: std_logic_vector(   0 downto 0);
        signal cVar1S6S55P015P068P051P053: std_logic_vector(   0 downto 0);
        signal cVar1S7S55P015P068P051N053: std_logic_vector(   0 downto 0);
        signal cVar1S8S55P015P068P009P010: std_logic_vector(   0 downto 0);
        signal cVar1S9S55P015P068P009N010: std_logic_vector(   0 downto 0);
        signal cVar1S10S55P015P068P009P066: std_logic_vector(   0 downto 0);
        signal cVar1S11S55N015P068P003P033: std_logic_vector(   0 downto 0);
        signal cVar1S12S55N015P068P003P033: std_logic_vector(   0 downto 0);
        signal cVar1S13S55N015P068P003P033: std_logic_vector(   0 downto 0);
        signal cVar1S14S55N015P068P003P033: std_logic_vector(   0 downto 0);
        signal cVar1S15S55N015P068P003P065: std_logic_vector(   0 downto 0);
        signal cVar1S16S55N015N068P069P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S55N015N068P069P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S55N015N068P069P008: std_logic_vector(   0 downto 0);
        signal cVar1S19S55N015N068P069P008: std_logic_vector(   0 downto 0);
        signal cVar1S20S55N015N068N069P004: std_logic_vector(   0 downto 0);
        signal cVar1S21S55N015N068N069P004: std_logic_vector(   0 downto 0);
        signal cVar1S22S55N015N068N069N004: std_logic_vector(   0 downto 0);
        signal cVar1S23S55N015N068N069N004: std_logic_vector(   0 downto 0);
        signal cVar1S24S55N015N068N069N004: std_logic_vector(   0 downto 0);
        signal cVar1S0S56P068P015P066P034: std_logic_vector(   0 downto 0);
        signal cVar1S1S56P068P015P066P034: std_logic_vector(   0 downto 0);
        signal cVar1S2S56P068P015P066P034: std_logic_vector(   0 downto 0);
        signal cVar1S3S56P068P015P066N034: std_logic_vector(   0 downto 0);
        signal cVar1S4S56P068P015P066N034: std_logic_vector(   0 downto 0);
        signal cVar1S5S56P068P015P066N034: std_logic_vector(   0 downto 0);
        signal cVar1S6S56P068P015P066N034: std_logic_vector(   0 downto 0);
        signal cVar1S7S56P068P015P066P008: std_logic_vector(   0 downto 0);
        signal cVar1S8S56P068P015P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S9S56P068P015P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S10S56P068P015P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S56P068P015P051P022: std_logic_vector(   0 downto 0);
        signal cVar1S12S56P068P015P051P053: std_logic_vector(   0 downto 0);
        signal cVar1S13S56P068P015P051N053: std_logic_vector(   0 downto 0);
        signal cVar1S14S56P068P009P024P052: std_logic_vector(   0 downto 0);
        signal cVar1S15S56P068P009P024P052: std_logic_vector(   0 downto 0);
        signal cVar1S16S56P068P009P024N052: std_logic_vector(   0 downto 0);
        signal cVar1S17S56P068P009P024N052: std_logic_vector(   0 downto 0);
        signal cVar1S18S56P068P009P024P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S56P068P009P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S20S56P068P009P002P066: std_logic_vector(   0 downto 0);
        signal cVar1S21S56P068P009P002P066: std_logic_vector(   0 downto 0);
        signal cVar1S0S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S1S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S2S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S3S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S4S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S5S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S6S57P015P051P009P037: std_logic_vector(   0 downto 0);
        signal cVar1S7S57P015P051P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S8S57P015P051P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S9S57P015P051P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S10S57P015P051P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S11S57P015P051P053P000: std_logic_vector(   0 downto 0);
        signal cVar1S12S57P015P051N053P014: std_logic_vector(   0 downto 0);
        signal cVar1S13S57N015P033P034P006: std_logic_vector(   0 downto 0);
        signal cVar1S14S57N015P033P034P006: std_logic_vector(   0 downto 0);
        signal cVar1S15S57N015P033N034P027: std_logic_vector(   0 downto 0);
        signal cVar1S16S57N015P033N034P027: std_logic_vector(   0 downto 0);
        signal cVar1S17S57N015P033N034N027: std_logic_vector(   0 downto 0);
        signal cVar1S18S57N015P033N034N027: std_logic_vector(   0 downto 0);
        signal cVar1S19S57N015P033N034N027: std_logic_vector(   0 downto 0);
        signal cVar1S20S57N015P033P064P056: std_logic_vector(   0 downto 0);
        signal cVar1S0S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S1S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S2S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S3S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S4S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S5S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S6S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S7S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S8S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S9S58P066P015P033P018: std_logic_vector(   0 downto 0);
        signal cVar1S10S58P066P015P033N018: std_logic_vector(   0 downto 0);
        signal cVar1S11S58P066P015P007P068: std_logic_vector(   0 downto 0);
        signal cVar1S12S58P066P015P007P068: std_logic_vector(   0 downto 0);
        signal cVar1S13S58P066P015P007P068: std_logic_vector(   0 downto 0);
        signal cVar1S14S58P066P015P007P068: std_logic_vector(   0 downto 0);
        signal cVar1S15S58P066P015P007P059: std_logic_vector(   0 downto 0);
        signal cVar1S16S58P066P009P024P045: std_logic_vector(   0 downto 0);
        signal cVar1S17S58P066P009P024P045: std_logic_vector(   0 downto 0);
        signal cVar1S18S58P066P009P024P045: std_logic_vector(   0 downto 0);
        signal cVar1S19S58P066P009P024P053: std_logic_vector(   0 downto 0);
        signal cVar1S20S58P066P009P002P037: std_logic_vector(   0 downto 0);
        signal cVar1S21S58P066P009P002P037: std_logic_vector(   0 downto 0);
        signal cVar1S22S58P066P009P002N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S59P018P008P050P067: std_logic_vector(   0 downto 0);
        signal cVar1S1S59P018P008P050P067: std_logic_vector(   0 downto 0);
        signal cVar1S2S59P018P008P050P067: std_logic_vector(   0 downto 0);
        signal cVar1S3S59P018P008P050N067: std_logic_vector(   0 downto 0);
        signal cVar1S4S59P018P008P050N067: std_logic_vector(   0 downto 0);
        signal cVar1S5S59P018P008P050P009: std_logic_vector(   0 downto 0);
        signal cVar1S6S59P018P008P050N009: std_logic_vector(   0 downto 0);
        signal cVar1S7S59P018P008P054P015: std_logic_vector(   0 downto 0);
        signal cVar1S8S59P018P008P054P015: std_logic_vector(   0 downto 0);
        signal cVar1S9S59P018P008P054P015: std_logic_vector(   0 downto 0);
        signal cVar1S10S59P018P008P054P015: std_logic_vector(   0 downto 0);
        signal cVar1S11S59N018P061P008P026: std_logic_vector(   0 downto 0);
        signal cVar1S12S59N018P061P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S13S59N018P061P008N026: std_logic_vector(   0 downto 0);
        signal cVar1S14S59N018P061N008P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S59N018P061N008P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S59N018P061N008N039: std_logic_vector(   0 downto 0);
        signal cVar1S17S59N018P061N008N039: std_logic_vector(   0 downto 0);
        signal cVar1S18S59N018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S19S59N018P061N059P063: std_logic_vector(   0 downto 0);
        signal cVar1S20S59N018P061N059N063: std_logic_vector(   0 downto 0);
        signal cVar1S0S60P018P061P067P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S60P018P061P067P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S60P018P061P067P010: std_logic_vector(   0 downto 0);
        signal cVar1S3S60P018P061P067N010: std_logic_vector(   0 downto 0);
        signal cVar1S4S60P018P061P067N010: std_logic_vector(   0 downto 0);
        signal cVar1S5S60P018P061P067N010: std_logic_vector(   0 downto 0);
        signal cVar1S6S60P018P061P067P013: std_logic_vector(   0 downto 0);
        signal cVar1S7S60P018P061P067P013: std_logic_vector(   0 downto 0);
        signal cVar1S8S60P018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S9S60P018P061N059P063: std_logic_vector(   0 downto 0);
        signal cVar1S10S60P018P061N059P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S60P018P061N059N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S60P018P067P019P056nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S60P018P067P019N056: std_logic_vector(   0 downto 0);
        signal cVar1S14S60P018P067P019N056: std_logic_vector(   0 downto 0);
        signal cVar1S15S60P018P067P019N056: std_logic_vector(   0 downto 0);
        signal cVar1S16S60P018P067P019P024: std_logic_vector(   0 downto 0);
        signal cVar1S17S60P018P067P019P024: std_logic_vector(   0 downto 0);
        signal cVar1S18S60P018P067P019P024: std_logic_vector(   0 downto 0);
        signal cVar1S19S60P018N067P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S20S60P018N067P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S21S60P018N067P069P030: std_logic_vector(   0 downto 0);
        signal cVar1S22S60P018N067P069P014: std_logic_vector(   0 downto 0);
        signal cVar1S0S61P018P008P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S1S61P018P008P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S2S61P018P008P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S3S61P018P008P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S4S61P018P008P024P034: std_logic_vector(   0 downto 0);
        signal cVar1S5S61P018P008P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S61P018P008P024N045: std_logic_vector(   0 downto 0);
        signal cVar1S7S61P018P008P024N045: std_logic_vector(   0 downto 0);
        signal cVar1S8S61P018P008P054P022: std_logic_vector(   0 downto 0);
        signal cVar1S9S61P018P008P054P022: std_logic_vector(   0 downto 0);
        signal cVar1S10S61N018P061P050P033: std_logic_vector(   0 downto 0);
        signal cVar1S11S61N018P061P050P033: std_logic_vector(   0 downto 0);
        signal cVar1S12S61N018P061N050P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S61N018P061N050P004: std_logic_vector(   0 downto 0);
        signal cVar1S14S61N018P061N050P004: std_logic_vector(   0 downto 0);
        signal cVar1S15S61N018P061N050N004: std_logic_vector(   0 downto 0);
        signal cVar1S16S61N018P061N050N004: std_logic_vector(   0 downto 0);
        signal cVar1S17S61N018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S18S61N018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S19S61N018P061N059P063: std_logic_vector(   0 downto 0);
        signal cVar1S20S61N018P061N059N063: std_logic_vector(   0 downto 0);
        signal cVar1S0S62P000P018P061P028: std_logic_vector(   0 downto 0);
        signal cVar1S1S62P000P018P061P028: std_logic_vector(   0 downto 0);
        signal cVar1S2S62P000P018P061N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S62P000P018P061N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S62P000P018P061N028: std_logic_vector(   0 downto 0);
        signal cVar1S5S62P000P018P061P059: std_logic_vector(   0 downto 0);
        signal cVar1S6S62P000P018P061N059: std_logic_vector(   0 downto 0);
        signal cVar1S7S62P000P018P061N059: std_logic_vector(   0 downto 0);
        signal cVar1S8S62P000P018P043P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S62P000P018P043P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S62P000P018P043P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S62P000P018P043P045: std_logic_vector(   0 downto 0);
        signal cVar1S12S62P000P030P027P056: std_logic_vector(   0 downto 0);
        signal cVar1S0S63P000P018P028P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S63P000P018P028N010: std_logic_vector(   0 downto 0);
        signal cVar1S2S63P000P018N028P030: std_logic_vector(   0 downto 0);
        signal cVar1S3S63P000P018N028P030: std_logic_vector(   0 downto 0);
        signal cVar1S4S63P000P018N028P030: std_logic_vector(   0 downto 0);
        signal cVar1S5S63P000P018N028P030: std_logic_vector(   0 downto 0);
        signal cVar1S6S63P000P018N028N030: std_logic_vector(   0 downto 0);
        signal cVar1S7S63P000P018N028N030: std_logic_vector(   0 downto 0);
        signal cVar1S8S63P000P018N028N030: std_logic_vector(   0 downto 0);
        signal cVar1S9S63P000P018P036P004: std_logic_vector(   0 downto 0);
        signal cVar1S10S63P000P018P036P004: std_logic_vector(   0 downto 0);
        signal cVar1S11S63P000P018P036P004: std_logic_vector(   0 downto 0);
        signal cVar1S12S63P000P018P036P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S63P000P018N036P057: std_logic_vector(   0 downto 0);
        signal cVar1S14S63P000P018N036P057: std_logic_vector(   0 downto 0);
        signal cVar1S15S63P000P018N036P057: std_logic_vector(   0 downto 0);
        signal cVar1S16S63P000P018N036P057: std_logic_vector(   0 downto 0);
        signal cVar1S17S63P000P030P027P020: std_logic_vector(   0 downto 0);
        signal cVar1S0S64P018P061P059P028: std_logic_vector(   0 downto 0);
        signal cVar1S1S64P018P061P059P028: std_logic_vector(   0 downto 0);
        signal cVar1S2S64P018P061P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S3S64P018P061P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S4S64P018P061P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S5S64P018P061P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S6S64P018P061P059P012: std_logic_vector(   0 downto 0);
        signal cVar1S7S64P018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S8S64P018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S9S64P018P061P059P000: std_logic_vector(   0 downto 0);
        signal cVar1S10S64P018P061N059P063: std_logic_vector(   0 downto 0);
        signal cVar1S11S64P018P061N059N063: std_logic_vector(   0 downto 0);
        signal cVar1S12S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S13S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S14S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S15S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S16S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S17S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S18S64P018P034P039P050: std_logic_vector(   0 downto 0);
        signal cVar1S19S64P018P034P039P068nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S64P018P034P047P069: std_logic_vector(   0 downto 0);
        signal cVar1S21S64P018P034P047P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S64P018P034P047P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S65P018P034P050P039: std_logic_vector(   0 downto 0);
        signal cVar1S1S65P018P034P050P039: std_logic_vector(   0 downto 0);
        signal cVar1S2S65P018P034P050P039: std_logic_vector(   0 downto 0);
        signal cVar1S3S65P018P034P050P039: std_logic_vector(   0 downto 0);
        signal cVar1S4S65P018P034P050P039: std_logic_vector(   0 downto 0);
        signal cVar1S5S65P018P034P050P048: std_logic_vector(   0 downto 0);
        signal cVar1S6S65P018P034P050N048: std_logic_vector(   0 downto 0);
        signal cVar1S7S65P018P034P050N048: std_logic_vector(   0 downto 0);
        signal cVar1S8S65P018P034P047P069: std_logic_vector(   0 downto 0);
        signal cVar1S9S65P018P034P047P069: std_logic_vector(   0 downto 0);
        signal cVar1S10S65N018P028P030P010: std_logic_vector(   0 downto 0);
        signal cVar1S11S65N018P028P030P010: std_logic_vector(   0 downto 0);
        signal cVar1S12S65N018P028P030P010: std_logic_vector(   0 downto 0);
        signal cVar1S13S65N018P028P030N010: std_logic_vector(   0 downto 0);
        signal cVar1S14S65N018N028P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S65N018N028P041P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S65N018N028P041N039: std_logic_vector(   0 downto 0);
        signal cVar1S17S65N018N028N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S18S65N018N028N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S19S65N018N028N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S20S65N018N028N041P039: std_logic_vector(   0 downto 0);
        signal cVar1S0S66P016P000P002P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S66P016P000P002N040: std_logic_vector(   0 downto 0);
        signal cVar1S2S66P016P000P002N040: std_logic_vector(   0 downto 0);
        signal cVar1S3S66P016P000N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S4S66P016P000N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S5S66P016P000N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S6S66P016P000N002P034: std_logic_vector(   0 downto 0);
        signal cVar1S7S66P016P000P053P031: std_logic_vector(   0 downto 0);
        signal cVar1S8S66P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S9S66P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S10S66P016P039P022P019: std_logic_vector(   0 downto 0);
        signal cVar1S11S66P016P039P007P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S66P016P039P007N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S67P014P024P027P044: std_logic_vector(   0 downto 0);
        signal cVar1S1S67P014P024P027P044: std_logic_vector(   0 downto 0);
        signal cVar1S2S67P014P024P027P044: std_logic_vector(   0 downto 0);
        signal cVar1S3S67P014P024P027P044: std_logic_vector(   0 downto 0);
        signal cVar1S4S67P014P024P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S67P014P024P031P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S67N014P027P009P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S67N014P027P009N050: std_logic_vector(   0 downto 0);
        signal cVar1S8S67N014P027N009P000: std_logic_vector(   0 downto 0);
        signal cVar1S9S67N014N027P050P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S67N014N027P050P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S67N014N027P050N024: std_logic_vector(   0 downto 0);
        signal cVar1S12S67N014N027P050N024: std_logic_vector(   0 downto 0);
        signal cVar1S13S67N014N027P050P032: std_logic_vector(   0 downto 0);
        signal cVar1S14S67N014N027P050P032: std_logic_vector(   0 downto 0);
        signal cVar1S15S67N014N027P050P032: std_logic_vector(   0 downto 0);
        signal cVar1S0S68P006P024P049P026: std_logic_vector(   0 downto 0);
        signal cVar1S1S68P006P024P049P026: std_logic_vector(   0 downto 0);
        signal cVar1S2S68P006P024P049P026: std_logic_vector(   0 downto 0);
        signal cVar1S3S68P006P024P049P026: std_logic_vector(   0 downto 0);
        signal cVar1S4S68P006P024P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S68P006P024P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S6S68P006P024P049N026: std_logic_vector(   0 downto 0);
        signal cVar1S7S68P006P024P010P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S68P006P024P010N047: std_logic_vector(   0 downto 0);
        signal cVar1S9S68P006P024P010N047: std_logic_vector(   0 downto 0);
        signal cVar1S10S68P006P024P010P019: std_logic_vector(   0 downto 0);
        signal cVar1S11S68P006P024P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S68P006P024P002P011: std_logic_vector(   0 downto 0);
        signal cVar1S13S68P006N024P065P034: std_logic_vector(   0 downto 0);
        signal cVar1S14S68P006N024P065P034: std_logic_vector(   0 downto 0);
        signal cVar1S15S68P006N024P065P034: std_logic_vector(   0 downto 0);
        signal cVar1S16S68P006N024P065P013: std_logic_vector(   0 downto 0);
        signal cVar1S0S69P055P026P010P057: std_logic_vector(   0 downto 0);
        signal cVar1S1S69P055P026P010P057: std_logic_vector(   0 downto 0);
        signal cVar1S2S69P055P026P010N057: std_logic_vector(   0 downto 0);
        signal cVar1S3S69P055P026N010P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S69P055P026N010N065: std_logic_vector(   0 downto 0);
        signal cVar1S5S69P055P026N010N065: std_logic_vector(   0 downto 0);
        signal cVar1S6S69N055P030P026P004: std_logic_vector(   0 downto 0);
        signal cVar1S7S69N055P030P026P004: std_logic_vector(   0 downto 0);
        signal cVar1S8S69N055P030N026P057: std_logic_vector(   0 downto 0);
        signal cVar1S9S69N055P030N026P057: std_logic_vector(   0 downto 0);
        signal cVar1S10S69N055P030P063P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S69N055P030P063N002: std_logic_vector(   0 downto 0);
        signal cVar1S12S69N055P030P063N002: std_logic_vector(   0 downto 0);
        signal cVar1S13S69N055P030P063N002: std_logic_vector(   0 downto 0);
        signal cVar1S14S69N055P030P063P014: std_logic_vector(   0 downto 0);
        signal cVar1S0S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S1S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S2S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S3S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S4S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S5S70P050P027P048P025: std_logic_vector(   0 downto 0);
        signal cVar1S6S70P050P027P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S70P050P027P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S8S70P050P027P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S9S70P050P027P048N025: std_logic_vector(   0 downto 0);
        signal cVar1S10S70P050P027P000P035: std_logic_vector(   0 downto 0);
        signal cVar1S11S70P050P027P000P035: std_logic_vector(   0 downto 0);
        signal cVar1S12S70P050P043P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S70P050P043P027N009: std_logic_vector(   0 downto 0);
        signal cVar1S14S70P050P043N027P020: std_logic_vector(   0 downto 0);
        signal cVar1S15S70P050P043N027P020: std_logic_vector(   0 downto 0);
        signal cVar1S0S71P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S71P021N040P048P039nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S71P021N040P048N039: std_logic_vector(   0 downto 0);
        signal cVar1S3S71N021P038P040P057: std_logic_vector(   0 downto 0);
        signal cVar1S4S71N021P038P040P057: std_logic_vector(   0 downto 0);
        signal cVar1S5S71N021P038P040N057: std_logic_vector(   0 downto 0);
        signal cVar1S6S71N021P038P040N057: std_logic_vector(   0 downto 0);
        signal cVar1S7S71N021P038P040N057: std_logic_vector(   0 downto 0);
        signal cVar1S8S71N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S71N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S71N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S11S71N021P038P040P015nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S71N021P038P040N015: std_logic_vector(   0 downto 0);
        signal cVar1S13S71N021P038N040P010nsss: std_logic_vector(   0 downto 0);
        signal cVar1S0S72P016P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S72P016P021N038P011: std_logic_vector(   0 downto 0);
        signal cVar1S2S72P016P021N038P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S72P016N021P040P038: std_logic_vector(   0 downto 0);
        signal cVar1S4S72P016N021P040P038: std_logic_vector(   0 downto 0);
        signal cVar1S5S72P016N021P040P038: std_logic_vector(   0 downto 0);
        signal cVar1S6S72P016N021P040P038: std_logic_vector(   0 downto 0);
        signal cVar1S7S72P016N021P040P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S72P016N021P040N002: std_logic_vector(   0 downto 0);
        signal cVar1S9S72P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S10S72P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S72P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S12S72P016P039P041P069: std_logic_vector(   0 downto 0);
        signal cVar1S13S72P016P039P054P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S72P016P039P054N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S73P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S73P021N040P048P056: std_logic_vector(   0 downto 0);
        signal cVar1S2S73P021N040P048P056: std_logic_vector(   0 downto 0);
        signal cVar1S3S73N021P038P040P057: std_logic_vector(   0 downto 0);
        signal cVar1S4S73N021P038P040P057: std_logic_vector(   0 downto 0);
        signal cVar1S5S73N021P038P040N057: std_logic_vector(   0 downto 0);
        signal cVar1S6S73N021P038P040N057: std_logic_vector(   0 downto 0);
        signal cVar1S7S73N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S8S73N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S73N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S73N021P038P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S73N021P038N020P063: std_logic_vector(   0 downto 0);
        signal cVar1S12S73N021P038N020P063: std_logic_vector(   0 downto 0);
        signal cVar1S0S74P014P027P002P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S74P014P027P002N009: std_logic_vector(   0 downto 0);
        signal cVar1S2S74P014P027P002N009: std_logic_vector(   0 downto 0);
        signal cVar1S3S74P014N027P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S4S74P014N027P010P028: std_logic_vector(   0 downto 0);
        signal cVar1S5S74P014N027P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S6S74P014N027P010N028: std_logic_vector(   0 downto 0);
        signal cVar1S7S74P014N027N010P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S74P014N027N010P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S74P014N027N010N024: std_logic_vector(   0 downto 0);
        signal cVar1S10S74P014N027N010N024: std_logic_vector(   0 downto 0);
        signal cVar1S11S74P014N027N010N024: std_logic_vector(   0 downto 0);
        signal cVar1S12S74P014N027N010N024: std_logic_vector(   0 downto 0);
        signal cVar1S13S74P014P024P044P037: std_logic_vector(   0 downto 0);
        signal cVar1S14S74P014P024P044N037: std_logic_vector(   0 downto 0);
        signal cVar1S15S74P014P024P044N037: std_logic_vector(   0 downto 0);
        signal cVar1S16S74P014P024P044N037: std_logic_vector(   0 downto 0);
        signal cVar1S17S74P014P024P044P065: std_logic_vector(   0 downto 0);
        signal cVar1S18S74P014P024P031P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S74P014P024P031N045: std_logic_vector(   0 downto 0);
        signal cVar1S20S74P014P024P031N045: std_logic_vector(   0 downto 0);
        signal cVar1S0S75P010P024P028P003: std_logic_vector(   0 downto 0);
        signal cVar1S1S75P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S2S75P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S3S75P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S4S75P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S5S75P010P024P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S6S75P010P024P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S7S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S11S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S12S75N010P014P024P056: std_logic_vector(   0 downto 0);
        signal cVar1S13S75N010P014P024P051: std_logic_vector(   0 downto 0);
        signal cVar1S14S75N010N014P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S75N010N014P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S16S75N010N014P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S17S75N010N014P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S18S75N010N014N027P024: std_logic_vector(   0 downto 0);
        signal cVar1S19S75N010N014N027P024: std_logic_vector(   0 downto 0);
        signal cVar1S20S75N010N014N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S21S75N010N014N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S22S75N010N014N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S0S76P014P010P032P021: std_logic_vector(   0 downto 0);
        signal cVar1S1S76P014P010P032P021: std_logic_vector(   0 downto 0);
        signal cVar1S2S76P014P010P032P017: std_logic_vector(   0 downto 0);
        signal cVar1S3S76P014N010P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S76P014N010P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S5S76P014N010P027N050: std_logic_vector(   0 downto 0);
        signal cVar1S6S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S8S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S9S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S10S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S76P014N010N027P050: std_logic_vector(   0 downto 0);
        signal cVar1S12S76P014P024P044P027: std_logic_vector(   0 downto 0);
        signal cVar1S13S76P014P024P044P027: std_logic_vector(   0 downto 0);
        signal cVar1S14S76P014P024P044P027: std_logic_vector(   0 downto 0);
        signal cVar1S15S76P014P024P044P027: std_logic_vector(   0 downto 0);
        signal cVar1S16S76P014P024P044P062: std_logic_vector(   0 downto 0);
        signal cVar1S17S76P014P024P031P045nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S76P014P024P031N045: std_logic_vector(   0 downto 0);
        signal cVar1S19S76P014P024P031N045: std_logic_vector(   0 downto 0);
        signal cVar1S0S77P010P024P028P003: std_logic_vector(   0 downto 0);
        signal cVar1S1S77P010P024P028P003: std_logic_vector(   0 downto 0);
        signal cVar1S2S77P010P024P028P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S77P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S4S77P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S5S77P010P024N028P045: std_logic_vector(   0 downto 0);
        signal cVar1S6S77P010P024P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S7S77P010P024P064P019: std_logic_vector(   0 downto 0);
        signal cVar1S8S77N010P025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S77N010P025N046P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S77N010P025N046N007: std_logic_vector(   0 downto 0);
        signal cVar1S11S77N010P025N046N007: std_logic_vector(   0 downto 0);
        signal cVar1S12S77N010N025P046P002: std_logic_vector(   0 downto 0);
        signal cVar1S13S77N010N025P046P002: std_logic_vector(   0 downto 0);
        signal cVar1S14S77N010N025P046P002: std_logic_vector(   0 downto 0);
        signal cVar1S15S77N010N025P046N002: std_logic_vector(   0 downto 0);
        signal cVar1S16S77N010N025P046P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S77N010N025P046N047: std_logic_vector(   0 downto 0);
        signal cVar1S18S77N010N025P046N047: std_logic_vector(   0 downto 0);
        signal cVar1S19S77N010N025P046N047: std_logic_vector(   0 downto 0);
        signal cVar1S0S78P039P041P020P050: std_logic_vector(   0 downto 0);
        signal cVar1S1S78P039P041P020N050: std_logic_vector(   0 downto 0);
        signal cVar1S2S78P039P041P020N050: std_logic_vector(   0 downto 0);
        signal cVar1S3S78P039P041P020N050: std_logic_vector(   0 downto 0);
        signal cVar1S4S78P039P041P020P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S78P039P041P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S6S78P039P041P020N040: std_logic_vector(   0 downto 0);
        signal cVar1S7S78P039P041P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S78P039P020P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S78P039N020P012P060: std_logic_vector(   0 downto 0);
        signal cVar1S10S78P039N020P012P060: std_logic_vector(   0 downto 0);
        signal cVar1S0S79P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S79P021N040P048P060: std_logic_vector(   0 downto 0);
        signal cVar1S2S79N021P038P040P050: std_logic_vector(   0 downto 0);
        signal cVar1S3S79N021P038P040P050: std_logic_vector(   0 downto 0);
        signal cVar1S4S79N021P038P040N050: std_logic_vector(   0 downto 0);
        signal cVar1S5S79N021P038P040N050: std_logic_vector(   0 downto 0);
        signal cVar1S6S79N021P038P040N050: std_logic_vector(   0 downto 0);
        signal cVar1S7S79N021P038P040N050: std_logic_vector(   0 downto 0);
        signal cVar1S8S79N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S9S79N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S10S79N021P038P040P059: std_logic_vector(   0 downto 0);
        signal cVar1S11S79N021P038P065P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S79N021P038P065N020: std_logic_vector(   0 downto 0);
        signal cVar1S13S79N021P038P065N020: std_logic_vector(   0 downto 0);
        signal cVar1S0S80P037P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S80P037P048N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S80P037P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S3S80P037P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S4S80P037P048N025N027: std_logic_vector(   0 downto 0);
        signal cVar1S5S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S6S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S7S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S8S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S9S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S10S80P037N048P046P064: std_logic_vector(   0 downto 0);
        signal cVar1S11S80P037N048P046P003: std_logic_vector(   0 downto 0);
        signal cVar1S12S80P037N048P046P003: std_logic_vector(   0 downto 0);
        signal cVar1S13S80P037P013P048P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S80P037P013P048P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S80P037P013P048N064: std_logic_vector(   0 downto 0);
        signal cVar1S16S80P037P013P048N064: std_logic_vector(   0 downto 0);
        signal cVar1S17S80P037P013P048P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S80P037P013P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S19S80P037P013P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S20S80P037P013P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S21S80P037P013P018P015: std_logic_vector(   0 downto 0);
        signal cVar1S22S80P037P013N018P031nsss: std_logic_vector(   0 downto 0);
        signal cVar1S23S80P037P013N018N031: std_logic_vector(   0 downto 0);
        signal cVar1S24S80P037P013N018N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S81P019P017P055P053: std_logic_vector(   0 downto 0);
        signal cVar1S1S81P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S2S81P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S3S81P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S4S81P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S5S81P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S6S81P019P017P064P029: std_logic_vector(   0 downto 0);
        signal cVar1S7S81P019P017P064P029: std_logic_vector(   0 downto 0);
        signal cVar1S8S81P019P017P064P029: std_logic_vector(   0 downto 0);
        signal cVar1S9S81P019P017P064P029: std_logic_vector(   0 downto 0);
        signal cVar1S10S81P019P017P064P011: std_logic_vector(   0 downto 0);
        signal cVar1S11S81P019P017P064P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S81P019P017P064N011: std_logic_vector(   0 downto 0);
        signal cVar1S13S81N019P037P003P035: std_logic_vector(   0 downto 0);
        signal cVar1S14S81N019P037P003P035: std_logic_vector(   0 downto 0);
        signal cVar1S15S81N019P037P003P035: std_logic_vector(   0 downto 0);
        signal cVar1S16S81N019P037P003P035: std_logic_vector(   0 downto 0);
        signal cVar1S17S81N019P037P003P035: std_logic_vector(   0 downto 0);
        signal cVar1S18S81N019P037P003P034nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S81N019P037P003N034: std_logic_vector(   0 downto 0);
        signal cVar1S20S81N019N037P048P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S81N019N037P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S22S81N019N037P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S23S81N019N037P048N062: std_logic_vector(   0 downto 0);
        signal cVar1S24S81N019N037N048P057: std_logic_vector(   0 downto 0);
        signal cVar1S25S81N019N037N048P057: std_logic_vector(   0 downto 0);
        signal cVar1S26S81N019N037N048P057: std_logic_vector(   0 downto 0);
        signal cVar1S27S81N019N037N048N057: std_logic_vector(   0 downto 0);
        signal cVar1S28S81N019N037N048N057: std_logic_vector(   0 downto 0);
        signal cVar1S29S81N019N037N048N057: std_logic_vector(   0 downto 0);
        signal cVar1S0S82P019P030P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S82P019P030P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S2S82P019P030P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S3S82P019P030N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S4S82P019P030N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S5S82P019P030N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S6S82P019P030P045P056nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S82P019P030P045N056: std_logic_vector(   0 downto 0);
        signal cVar1S8S82P019P030P045N056: std_logic_vector(   0 downto 0);
        signal cVar1S9S82P019P030P045N056: std_logic_vector(   0 downto 0);
        signal cVar1S10S82P019P017P055P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S82P019P017P055N065: std_logic_vector(   0 downto 0);
        signal cVar1S12S82P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S13S82P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S14S82P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S15S82P019P017N055P057: std_logic_vector(   0 downto 0);
        signal cVar1S16S82P019P017P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S17S82P019P017P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S18S82P019P017P053P037: std_logic_vector(   0 downto 0);
        signal cVar1S19S82P019P017P053N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S83P015P051P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S1S83P015P051P017P012: std_logic_vector(   0 downto 0);
        signal cVar1S2S83P015P051P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S3S83P015P051P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S4S83P015P051P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S5S83P015P051P017N012: std_logic_vector(   0 downto 0);
        signal cVar1S6S83P015P051P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S7S83P015P051P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S8S83P015P051P017P061: std_logic_vector(   0 downto 0);
        signal cVar1S9S83P015P051P053P000: std_logic_vector(   0 downto 0);
        signal cVar1S10S83P015P051P053P000: std_logic_vector(   0 downto 0);
        signal cVar1S11S83P015P051N053P014: std_logic_vector(   0 downto 0);
        signal cVar1S12S83N015P021P038nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S83N015P021N038P069: std_logic_vector(   0 downto 0);
        signal cVar1S14S83N015P021N038P069: std_logic_vector(   0 downto 0);
        signal cVar1S15S83N015N021P038P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S83N015N021P038P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S83N015N021P038P067: std_logic_vector(   0 downto 0);
        signal cVar1S18S83N015N021P038N067: std_logic_vector(   0 downto 0);
        signal cVar1S19S83N015N021P038N067: std_logic_vector(   0 downto 0);
        signal cVar1S20S83N015N021P038N067: std_logic_vector(   0 downto 0);
        signal cVar1S21S83N015N021P038P069: std_logic_vector(   0 downto 0);
        signal cVar1S22S83N015N021P038P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S84P067P037P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S84P067P037P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S2S84P067P037P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S3S84P067P037N021P013: std_logic_vector(   0 downto 0);
        signal cVar1S4S84P067P037N021P013: std_logic_vector(   0 downto 0);
        signal cVar1S5S84P067P037N021P013: std_logic_vector(   0 downto 0);
        signal cVar1S6S84P067P037N021N013: std_logic_vector(   0 downto 0);
        signal cVar1S7S84P067P037N021N013: std_logic_vector(   0 downto 0);
        signal cVar1S8S84P067P037N021N013: std_logic_vector(   0 downto 0);
        signal cVar1S9S84P067P037P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S84P067P037N028P013: std_logic_vector(   0 downto 0);
        signal cVar1S11S84P067P037N028P013: std_logic_vector(   0 downto 0);
        signal cVar1S12S84P067P037N028P013: std_logic_vector(   0 downto 0);
        signal cVar1S13S84P067P037N028P013: std_logic_vector(   0 downto 0);
        signal cVar1S14S84P067P037N028P013: std_logic_vector(   0 downto 0);
        signal cVar1S15S84P067P051P065P010: std_logic_vector(   0 downto 0);
        signal cVar1S16S84P067P051P065P010: std_logic_vector(   0 downto 0);
        signal cVar1S17S84P067P051P065P010: std_logic_vector(   0 downto 0);
        signal cVar1S18S84P067P051N065P064: std_logic_vector(   0 downto 0);
        signal cVar1S19S84P067P051N065N064: std_logic_vector(   0 downto 0);
        signal cVar1S20S84P067P051N065N064: std_logic_vector(   0 downto 0);
        signal cVar1S21S84P067P051N065N064: std_logic_vector(   0 downto 0);
        signal cVar1S22S84P067P051P006P034: std_logic_vector(   0 downto 0);
        signal cVar1S0S85P037P013P048P055: std_logic_vector(   0 downto 0);
        signal cVar1S1S85P037P013P048P055: std_logic_vector(   0 downto 0);
        signal cVar1S2S85P037P013P048N055: std_logic_vector(   0 downto 0);
        signal cVar1S3S85P037P013P048N055: std_logic_vector(   0 downto 0);
        signal cVar1S4S85P037P013P048N055: std_logic_vector(   0 downto 0);
        signal cVar1S5S85P037P013P048P035: std_logic_vector(   0 downto 0);
        signal cVar1S6S85P037P013P018P050: std_logic_vector(   0 downto 0);
        signal cVar1S7S85P037P013P018P050: std_logic_vector(   0 downto 0);
        signal cVar1S8S85P037P013P018P050: std_logic_vector(   0 downto 0);
        signal cVar1S9S85P037P013P018P050: std_logic_vector(   0 downto 0);
        signal cVar1S10S85P037P013N018P041: std_logic_vector(   0 downto 0);
        signal cVar1S11S85P037P013N018P041: std_logic_vector(   0 downto 0);
        signal cVar1S12S85N037P058P011P031nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S85N037P058P011N031: std_logic_vector(   0 downto 0);
        signal cVar1S14S85N037P058P011N031: std_logic_vector(   0 downto 0);
        signal cVar1S15S85N037P058P011N031: std_logic_vector(   0 downto 0);
        signal cVar1S16S85N037P058P011N031: std_logic_vector(   0 downto 0);
        signal cVar1S17S85N037P058P011P009: std_logic_vector(   0 downto 0);
        signal cVar1S18S85N037P058P011P009: std_logic_vector(   0 downto 0);
        signal cVar1S19S85N037N058P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar1S20S85N037N058P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S21S85N037N058P021N040: std_logic_vector(   0 downto 0);
        signal cVar1S22S85N037N058N021P048: std_logic_vector(   0 downto 0);
        signal cVar1S23S85N037N058N021P048: std_logic_vector(   0 downto 0);
        signal cVar1S24S85N037N058N021P048: std_logic_vector(   0 downto 0);
        signal cVar1S25S85N037N058N021N048: std_logic_vector(   0 downto 0);
        signal cVar1S0S86P037P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S86P037P048N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S2S86P037P048N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S3S86P037P048N025N050: std_logic_vector(   0 downto 0);
        signal cVar1S4S86P037P048N025N050: std_logic_vector(   0 downto 0);
        signal cVar1S5S86P037N048P046P036: std_logic_vector(   0 downto 0);
        signal cVar1S6S86P037N048P046P036: std_logic_vector(   0 downto 0);
        signal cVar1S7S86P037N048P046P036: std_logic_vector(   0 downto 0);
        signal cVar1S8S86P037N048P046N036: std_logic_vector(   0 downto 0);
        signal cVar1S9S86P037N048P046N036: std_logic_vector(   0 downto 0);
        signal cVar1S10S86P037N048P046N036: std_logic_vector(   0 downto 0);
        signal cVar1S11S86P037N048P046P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S86P037N048P046P062: std_logic_vector(   0 downto 0);
        signal cVar1S13S86P037P004P031P035: std_logic_vector(   0 downto 0);
        signal cVar1S14S86P037P004N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S15S86P037P004N031P055: std_logic_vector(   0 downto 0);
        signal cVar1S16S86P037P004N031N055: std_logic_vector(   0 downto 0);
        signal cVar1S17S86P037P004N031N055: std_logic_vector(   0 downto 0);
        signal cVar1S18S86P037P004P051P036: std_logic_vector(   0 downto 0);
        signal cVar1S19S86P037P004P051P036: std_logic_vector(   0 downto 0);
        signal cVar1S0S87P019P017P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S1S87P019P017P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S2S87P019P017P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S3S87P019P017P035P026: std_logic_vector(   0 downto 0);
        signal cVar1S4S87P019P017N035P066: std_logic_vector(   0 downto 0);
        signal cVar1S5S87P019P017N035P066: std_logic_vector(   0 downto 0);
        signal cVar1S6S87P019P017N035P066: std_logic_vector(   0 downto 0);
        signal cVar1S7S87P019P017N035N066: std_logic_vector(   0 downto 0);
        signal cVar1S8S87P019P017N035N066: std_logic_vector(   0 downto 0);
        signal cVar1S9S87P019P017N035N066: std_logic_vector(   0 downto 0);
        signal cVar1S10S87P019P017P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S11S87P019P017P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S12S87P019P017P053P029: std_logic_vector(   0 downto 0);
        signal cVar1S13S87P019P017P053P037: std_logic_vector(   0 downto 0);
        signal cVar1S14S87N019P009P068P039: std_logic_vector(   0 downto 0);
        signal cVar1S15S87N019P009P068P039: std_logic_vector(   0 downto 0);
        signal cVar1S16S87N019P009P068P039: std_logic_vector(   0 downto 0);
        signal cVar1S17S87N019P009P068P053nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S87N019N009P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar1S19S87N019N009P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S20S87N019N009P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S21S87N019N009P040N021: std_logic_vector(   0 downto 0);
        signal cVar1S22S87N019N009N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S23S87N019N009N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S24S87N019N009N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S25S87N019N009N040P038: std_logic_vector(   0 downto 0);
        signal cVar1S0S88P060P009P068P063: std_logic_vector(   0 downto 0);
        signal cVar1S1S88P060P009P068P063: std_logic_vector(   0 downto 0);
        signal cVar1S2S88P060P009P068P063: std_logic_vector(   0 downto 0);
        signal cVar1S3S88P060P009P068P063: std_logic_vector(   0 downto 0);
        signal cVar1S4S88P060P009P068P063: std_logic_vector(   0 downto 0);
        signal cVar1S5S88P060P009P068P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S88P060P009P068P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S88P060N009P053P055: std_logic_vector(   0 downto 0);
        signal cVar1S8S88P060N009P053N055: std_logic_vector(   0 downto 0);
        signal cVar1S9S88P060N009P053N055: std_logic_vector(   0 downto 0);
        signal cVar1S10S88P060N009P053N055: std_logic_vector(   0 downto 0);
        signal cVar1S11S88P060N009P053P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S88P060N009P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S13S88P060N009P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S14S88P060N009P053N028: std_logic_vector(   0 downto 0);
        signal cVar1S15S88P060P039P062P051: std_logic_vector(   0 downto 0);
        signal cVar1S16S88P060P039P062P051: std_logic_vector(   0 downto 0);
        signal cVar1S17S88P060P039N062P031: std_logic_vector(   0 downto 0);
        signal cVar1S18S88P060P039N062P031: std_logic_vector(   0 downto 0);
        signal cVar1S19S88P060P039N062N031: std_logic_vector(   0 downto 0);
        signal cVar1S20S88P060P039N062N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S89P009P068P063P007: std_logic_vector(   0 downto 0);
        signal cVar1S1S89P009P068P063P007: std_logic_vector(   0 downto 0);
        signal cVar1S2S89P009P068P063N007: std_logic_vector(   0 downto 0);
        signal cVar1S3S89P009P068P063P008: std_logic_vector(   0 downto 0);
        signal cVar1S4S89P009P068P002P047nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S89P009P068P002N047: std_logic_vector(   0 downto 0);
        signal cVar1S6S89P009P068P002N047: std_logic_vector(   0 downto 0);
        signal cVar1S7S89N009P049P023P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S89N009P049P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S9S89N009P049P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S10S89N009P049P023N005: std_logic_vector(   0 downto 0);
        signal cVar1S11S89N009P049N023P043: std_logic_vector(   0 downto 0);
        signal cVar1S12S89N009P049N023P043: std_logic_vector(   0 downto 0);
        signal cVar1S13S89N009P049N023P043: std_logic_vector(   0 downto 0);
        signal cVar1S14S89N009P049N023P043: std_logic_vector(   0 downto 0);
        signal cVar1S15S89N009P049N023P043: std_logic_vector(   0 downto 0);
        signal cVar1S16S89N009P049P026P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S89N009P049N026P024: std_logic_vector(   0 downto 0);
        signal cVar1S18S89N009P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S19S89N009P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S20S89N009P049N026N024: std_logic_vector(   0 downto 0);
        signal cVar1S0S90P049P052P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S90P049P052N065P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S90P049P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S3S90P049P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S4S90P049P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S5S90P049P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S6S90P049N052P029P055: std_logic_vector(   0 downto 0);
        signal cVar1S7S90P049N052P029P055: std_logic_vector(   0 downto 0);
        signal cVar1S8S90P049N052P029N055: std_logic_vector(   0 downto 0);
        signal cVar1S9S90P049N052P029N055: std_logic_vector(   0 downto 0);
        signal cVar1S10S90P049N052P029N055: std_logic_vector(   0 downto 0);
        signal cVar1S11S90P049N052P029N055: std_logic_vector(   0 downto 0);
        signal cVar1S12S90P049N052P029P056: std_logic_vector(   0 downto 0);
        signal cVar1S13S90P049N052P029N056: std_logic_vector(   0 downto 0);
        signal cVar1S14S90P049P026P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S90P049N026P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S90P049N026N027P024: std_logic_vector(   0 downto 0);
        signal cVar1S17S90P049N026N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S18S90P049N026N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S19S90P049N026N027N024: std_logic_vector(   0 downto 0);
        signal cVar1S0S91P052P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S91P052N065P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S91P052N065N062P050: std_logic_vector(   0 downto 0);
        signal cVar1S3S91P052N065N062P050: std_logic_vector(   0 downto 0);
        signal cVar1S4S91P052N065N062N050: std_logic_vector(   0 downto 0);
        signal cVar1S5S91P052N065N062N050: std_logic_vector(   0 downto 0);
        signal cVar1S6S91P052N065N062N050: std_logic_vector(   0 downto 0);
        signal cVar1S7S91N052P048P061P007: std_logic_vector(   0 downto 0);
        signal cVar1S8S91N052P048P061P007: std_logic_vector(   0 downto 0);
        signal cVar1S9S91N052P048P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S10S91N052P048P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S11S91N052P048P061N007: std_logic_vector(   0 downto 0);
        signal cVar1S12S91N052P048P061P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S91N052N048P050P055: std_logic_vector(   0 downto 0);
        signal cVar1S14S91N052N048P050N055: std_logic_vector(   0 downto 0);
        signal cVar1S15S91N052N048P050P004: std_logic_vector(   0 downto 0);
        signal cVar1S0S92P019P068P029P054nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S92P019P068P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S2S92P019P068P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S3S92P019P068P029N054: std_logic_vector(   0 downto 0);
        signal cVar1S4S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S5S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S6S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S7S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S8S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S9S92P019P068N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S10S92P019P068P055P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S92P019P068P055N050: std_logic_vector(   0 downto 0);
        signal cVar1S12S92P019P068P055P010nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S92P019P066P009P046nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S92P019P066P009N046: std_logic_vector(   0 downto 0);
        signal cVar1S15S92P019P066P009N046: std_logic_vector(   0 downto 0);
        signal cVar1S16S92P019P066P009N046: std_logic_vector(   0 downto 0);
        signal cVar1S17S92P019P066P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S18S92P019P066P009P068: std_logic_vector(   0 downto 0);
        signal cVar1S19S92P019N066P051P061: std_logic_vector(   0 downto 0);
        signal cVar1S20S92P019N066P051P061: std_logic_vector(   0 downto 0);
        signal cVar1S21S92P019N066P051P061: std_logic_vector(   0 downto 0);
        signal cVar1S22S92P019N066P051P061: std_logic_vector(   0 downto 0);
        signal cVar1S23S92P019N066P051P061: std_logic_vector(   0 downto 0);
        signal cVar1S24S92P019N066P051P016: std_logic_vector(   0 downto 0);
        signal cVar1S25S92P019N066P051P016: std_logic_vector(   0 downto 0);
        signal cVar1S26S92P019N066P051P016: std_logic_vector(   0 downto 0);
        signal cVar1S0S93P019P051P002P000: std_logic_vector(   0 downto 0);
        signal cVar1S1S93P019P051P002P000: std_logic_vector(   0 downto 0);
        signal cVar1S2S93P019P051P002P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S93P019P051P002N000: std_logic_vector(   0 downto 0);
        signal cVar1S4S93P019P051P002N000: std_logic_vector(   0 downto 0);
        signal cVar1S5S93P019P051P002N000: std_logic_vector(   0 downto 0);
        signal cVar1S6S93P019P051P002N000: std_logic_vector(   0 downto 0);
        signal cVar1S7S93P019P051P002P054: std_logic_vector(   0 downto 0);
        signal cVar1S8S93P019P051P024P037: std_logic_vector(   0 downto 0);
        signal cVar1S9S93P019P051P024N037: std_logic_vector(   0 downto 0);
        signal cVar1S10S93P019P051P024N037: std_logic_vector(   0 downto 0);
        signal cVar1S11S93N019P056P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S93N019P056P054N013: std_logic_vector(   0 downto 0);
        signal cVar1S13S93N019P056N054P058: std_logic_vector(   0 downto 0);
        signal cVar1S14S93N019P056N054P058: std_logic_vector(   0 downto 0);
        signal cVar1S15S93N019P056N054N058: std_logic_vector(   0 downto 0);
        signal cVar1S16S93N019N056P054P037: std_logic_vector(   0 downto 0);
        signal cVar1S17S93N019N056P054P037: std_logic_vector(   0 downto 0);
        signal cVar1S18S93N019N056P054N037: std_logic_vector(   0 downto 0);
        signal cVar1S19S93N019N056P054N037: std_logic_vector(   0 downto 0);
        signal cVar1S20S93N019N056P054N037: std_logic_vector(   0 downto 0);
        signal cVar1S21S93N019N056P054P005: std_logic_vector(   0 downto 0);
        signal cVar1S22S93N019N056P054P005: std_logic_vector(   0 downto 0);
        signal cVar1S0S94P019P037P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S1S94P019P037P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S2S94P019P037P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S94P019P037P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S4S94P019P037P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S5S94P019P037P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S6S94P019P037N029P045: std_logic_vector(   0 downto 0);
        signal cVar1S7S94P019P037N029P045: std_logic_vector(   0 downto 0);
        signal cVar1S8S94P019P037N029P045: std_logic_vector(   0 downto 0);
        signal cVar1S9S94P019P037N029N045: std_logic_vector(   0 downto 0);
        signal cVar1S10S94P019P037N029N045: std_logic_vector(   0 downto 0);
        signal cVar1S11S94P019P037P059P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S94P019P037P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S13S94P019P037P059P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S94P019P037P059P064: std_logic_vector(   0 downto 0);
        signal cVar1S15S94P019P069P051P029: std_logic_vector(   0 downto 0);
        signal cVar1S16S94P019P069P051P029: std_logic_vector(   0 downto 0);
        signal cVar1S17S94P019P069P051P013: std_logic_vector(   0 downto 0);
        signal cVar1S18S94P019N069P057P030: std_logic_vector(   0 downto 0);
        signal cVar1S19S94P019N069P057P030: std_logic_vector(   0 downto 0);
        signal cVar1S20S94P019N069P057P030: std_logic_vector(   0 downto 0);
        signal cVar1S21S94P019N069P057P061: std_logic_vector(   0 downto 0);
        signal cVar1S22S94P019N069P057P061: std_logic_vector(   0 downto 0);
        signal cVar1S23S94P019N069P057P061: std_logic_vector(   0 downto 0);
        signal cVar1S0S95P019P057P036P009: std_logic_vector(   0 downto 0);
        signal cVar1S1S95P019P057P036P009: std_logic_vector(   0 downto 0);
        signal cVar1S2S95P019P057P036P009: std_logic_vector(   0 downto 0);
        signal cVar1S3S95P019P057P036N009: std_logic_vector(   0 downto 0);
        signal cVar1S4S95P019P057P036N009: std_logic_vector(   0 downto 0);
        signal cVar1S5S95P019P057N036P056: std_logic_vector(   0 downto 0);
        signal cVar1S6S95P019P057N036P056: std_logic_vector(   0 downto 0);
        signal cVar1S7S95P019P057N036P056: std_logic_vector(   0 downto 0);
        signal cVar1S8S95P019P057N036P056: std_logic_vector(   0 downto 0);
        signal cVar1S9S95P019P057N036P056: std_logic_vector(   0 downto 0);
        signal cVar1S10S95P019P057P030P056nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S95P019P057P030N056: std_logic_vector(   0 downto 0);
        signal cVar1S12S95P019P057N030P004: std_logic_vector(   0 downto 0);
        signal cVar1S13S95N019P045P062P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S95N019P045P062N005: std_logic_vector(   0 downto 0);
        signal cVar1S15S95N019P045P062N005: std_logic_vector(   0 downto 0);
        signal cVar1S16S95N019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S17S95N019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S18S95N019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S19S95N019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S20S95N019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S21S95N019N045N029P031: std_logic_vector(   0 downto 0);
        signal cVar1S22S95N019N045N029P031: std_logic_vector(   0 downto 0);
        signal cVar1S23S95N019N045N029P031: std_logic_vector(   0 downto 0);
        signal cVar1S24S95N019N045N029N031: std_logic_vector(   0 downto 0);
        signal cVar1S25S95N019N045N029N031: std_logic_vector(   0 downto 0);
        signal cVar1S26S95N019N045N029N031: std_logic_vector(   0 downto 0);
        signal cVar1S0S96P019P037P045P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S96P019P037P045N005: std_logic_vector(   0 downto 0);
        signal cVar1S2S96P019P037P045N005: std_logic_vector(   0 downto 0);
        signal cVar1S3S96P019P037N045P029: std_logic_vector(   0 downto 0);
        signal cVar1S4S96P019P037N045P029: std_logic_vector(   0 downto 0);
        signal cVar1S5S96P019P037N045P029: std_logic_vector(   0 downto 0);
        signal cVar1S6S96P019P037N045N029: std_logic_vector(   0 downto 0);
        signal cVar1S7S96P019P037N045N029: std_logic_vector(   0 downto 0);
        signal cVar1S8S96P019P037N045N029: std_logic_vector(   0 downto 0);
        signal cVar1S9S96P019P037P059P028nsss: std_logic_vector(   0 downto 0);
        signal cVar1S10S96P019P037P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S11S96P019P037P059N028: std_logic_vector(   0 downto 0);
        signal cVar1S12S96P019P037P059P064: std_logic_vector(   0 downto 0);
        signal cVar1S13S96P019P037P059P064: std_logic_vector(   0 downto 0);
        signal cVar1S14S96P019P036P006P009: std_logic_vector(   0 downto 0);
        signal cVar1S15S96P019P036P006N009: std_logic_vector(   0 downto 0);
        signal cVar1S16S96P019P036P006N009: std_logic_vector(   0 downto 0);
        signal cVar1S17S96P019P036P006N009: std_logic_vector(   0 downto 0);
        signal cVar1S18S96P019P036P006P004: std_logic_vector(   0 downto 0);
        signal cVar1S19S96P019P036P006P004: std_logic_vector(   0 downto 0);
        signal cVar1S20S96P019N036P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S21S96P019N036P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S22S96P019N036P009P063: std_logic_vector(   0 downto 0);
        signal cVar1S23S96P019N036P009N063: std_logic_vector(   0 downto 0);
        signal cVar1S24S96P019N036P009N063: std_logic_vector(   0 downto 0);
        signal cVar1S25S96P019N036P009N063: std_logic_vector(   0 downto 0);
        signal cVar1S26S96P019N036P009P028: std_logic_vector(   0 downto 0);
        signal cVar1S0S97P045P035P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S97P045P035N025P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S97P045P035N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S3S97P045P035N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S4S97N045P043P019P023: std_logic_vector(   0 downto 0);
        signal cVar1S5S97N045P043P019P023: std_logic_vector(   0 downto 0);
        signal cVar1S6S97N045P043P019P023: std_logic_vector(   0 downto 0);
        signal cVar1S7S97N045P043N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S97N045P043N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S97N045P043N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S97N045P043N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S97N045P043N019P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S97N045P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S97N045P043N022P057nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S97N045P043N022N057: std_logic_vector(   0 downto 0);
        signal cVar1S0S98P019P045P026P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S98P019P045P026P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S98P019N045P024P029: std_logic_vector(   0 downto 0);
        signal cVar1S3S98P019N045P024P029: std_logic_vector(   0 downto 0);
        signal cVar1S4S98P019N045P024N029: std_logic_vector(   0 downto 0);
        signal cVar1S5S98P019N045P024N029: std_logic_vector(   0 downto 0);
        signal cVar1S6S98P019N045P024N029: std_logic_vector(   0 downto 0);
        signal cVar1S7S98P019N045P024P001: std_logic_vector(   0 downto 0);
        signal cVar1S8S98P019P051P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S98P019P051P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S10S98P019P051P025P016: std_logic_vector(   0 downto 0);
        signal cVar1S11S98P019P051N025P029: std_logic_vector(   0 downto 0);
        signal cVar1S12S98P019P051N025P029: std_logic_vector(   0 downto 0);
        signal cVar1S13S98P019P051N025P029: std_logic_vector(   0 downto 0);
        signal cVar1S14S98P019P051N025P029: std_logic_vector(   0 downto 0);
        signal cVar1S15S98P019P051N025P029: std_logic_vector(   0 downto 0);
        signal cVar1S16S98P019P051P037P024: std_logic_vector(   0 downto 0);
        signal cVar1S17S98P019P051N037P008: std_logic_vector(   0 downto 0);
        signal cVar1S18S98P019P051N037N008: std_logic_vector(   0 downto 0);
        signal cVar1S0S99P045P030P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S99P045P030N025P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S99P045P030N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S3S99P045P030N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S4S99N045P019P043P051: std_logic_vector(   0 downto 0);
        signal cVar1S5S99N045P019P043P051: std_logic_vector(   0 downto 0);
        signal cVar1S6S99N045P019P043P051: std_logic_vector(   0 downto 0);
        signal cVar1S7S99N045P019P043P051: std_logic_vector(   0 downto 0);
        signal cVar1S8S99N045P019P043P051: std_logic_vector(   0 downto 0);
        signal cVar1S9S99N045P019P043P014: std_logic_vector(   0 downto 0);
        signal cVar1S10S99N045P019P043P014: std_logic_vector(   0 downto 0);
        signal cVar1S11S99N045N019P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S12S99N045N019P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S13S99N045N019P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S14S99N045N019P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S15S99N045N019P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S16S99N045N019N029P032: std_logic_vector(   0 downto 0);
        signal cVar1S17S99N045N019N029P032: std_logic_vector(   0 downto 0);
        signal cVar1S18S99N045N019N029N032: std_logic_vector(   0 downto 0);
        signal cVar1S19S99N045N019N029N032: std_logic_vector(   0 downto 0);
        signal cVar1S0S100P019P045P026P062: std_logic_vector(   0 downto 0);
        signal cVar1S1S100P019P045P026P062: std_logic_vector(   0 downto 0);
        signal cVar1S2S100P019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S100P019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S4S100P019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S5S100P019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S6S100P019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S7S100P019N045N029P008: std_logic_vector(   0 downto 0);
        signal cVar1S8S100P019N045N029P008: std_logic_vector(   0 downto 0);
        signal cVar1S9S100P019N045N029P008: std_logic_vector(   0 downto 0);
        signal cVar1S10S100P019N045N029P008: std_logic_vector(   0 downto 0);
        signal cVar1S11S100P019N045N029P008: std_logic_vector(   0 downto 0);
        signal cVar1S12S100P019P013P045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S100P019P013P045N043: std_logic_vector(   0 downto 0);
        signal cVar1S14S100P019P013P045N043: std_logic_vector(   0 downto 0);
        signal cVar1S15S100P019P013N045P067: std_logic_vector(   0 downto 0);
        signal cVar1S16S100P019P013N045P067: std_logic_vector(   0 downto 0);
        signal cVar1S17S100P019P013N045N067: std_logic_vector(   0 downto 0);
        signal cVar1S18S100P019P013N045N067: std_logic_vector(   0 downto 0);
        signal cVar1S19S100P019P013P039P041: std_logic_vector(   0 downto 0);
        signal cVar1S0S101P045P030P035P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S101P045P030P035N025: std_logic_vector(   0 downto 0);
        signal cVar1S2S101P045P030P035N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S101P045P030P035N025: std_logic_vector(   0 downto 0);
        signal cVar1S4S101N045P019P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S5S101N045P019P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S6S101N045P019P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S7S101N045P019P043P023: std_logic_vector(   0 downto 0);
        signal cVar1S8S101N045P019P043P014: std_logic_vector(   0 downto 0);
        signal cVar1S9S101N045P019P043P014: std_logic_vector(   0 downto 0);
        signal cVar1S10S101N045N019P029P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S101N045N019P029P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S101N045N019N029P040: std_logic_vector(   0 downto 0);
        signal cVar1S13S101N045N019N029P040: std_logic_vector(   0 downto 0);
        signal cVar1S0S102P019P045P026P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S102P019P045P026N005: std_logic_vector(   0 downto 0);
        signal cVar1S2S102P019N045P029P061: std_logic_vector(   0 downto 0);
        signal cVar1S3S102P019N045P029P061: std_logic_vector(   0 downto 0);
        signal cVar1S4S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S5S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S6S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S7S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S8S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S9S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S10S102P019N045N029P054: std_logic_vector(   0 downto 0);
        signal cVar1S11S102P019P051P018P057: std_logic_vector(   0 downto 0);
        signal cVar1S12S102P019P051P018P057: std_logic_vector(   0 downto 0);
        signal cVar1S13S102P019P051P018P057: std_logic_vector(   0 downto 0);
        signal cVar1S14S102P019P051P018P057: std_logic_vector(   0 downto 0);
        signal cVar1S15S102P019P051N018P053: std_logic_vector(   0 downto 0);
        signal cVar1S16S102P019P051N018P053: std_logic_vector(   0 downto 0);
        signal cVar1S17S102P019P051N018P053: std_logic_vector(   0 downto 0);
        signal cVar1S18S102P019P051N018P053: std_logic_vector(   0 downto 0);
        signal cVar1S19S102P019P051P024P037: std_logic_vector(   0 downto 0);
        signal cVar1S20S102P019P051P024N037: std_logic_vector(   0 downto 0);
        signal cVar1S0S103P045P030P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S103P045P030N025P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S103P045P030N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S3S103P045P030N025N022: std_logic_vector(   0 downto 0);
        signal cVar1S4S103N045P052P065nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S103N045P052N065P062nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S103N045P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S7S103N045P052N065N062: std_logic_vector(   0 downto 0);
        signal cVar1S8S103N045N052P043P018: std_logic_vector(   0 downto 0);
        signal cVar1S9S103N045N052P043P018: std_logic_vector(   0 downto 0);
        signal cVar1S10S103N045N052P043P018: std_logic_vector(   0 downto 0);
        signal cVar1S11S103N045N052P043P018: std_logic_vector(   0 downto 0);
        signal cVar1S12S103N045N052P043P018: std_logic_vector(   0 downto 0);
        signal cVar1S13S103N045N052P043P063: std_logic_vector(   0 downto 0);
        signal cVar1S14S103N045N052P043P063: std_logic_vector(   0 downto 0);
        signal cVar1S0S104P019P045P026P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S104P019P045P026N005: std_logic_vector(   0 downto 0);
        signal cVar1S2S104P019N045P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S3S104P019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S4S104P019N045P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S5S104P019N045N029P069: std_logic_vector(   0 downto 0);
        signal cVar1S6S104P019N045N029P069: std_logic_vector(   0 downto 0);
        signal cVar1S7S104P019N045N029P069: std_logic_vector(   0 downto 0);
        signal cVar1S8S104P019N045N029P069: std_logic_vector(   0 downto 0);
        signal cVar1S9S104P019N045N029P069: std_logic_vector(   0 downto 0);
        signal cVar1S10S104P019P067P047P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S104P019P067P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S12S104P019P067P047N006: std_logic_vector(   0 downto 0);
        signal cVar1S13S104P019P067N047P069: std_logic_vector(   0 downto 0);
        signal cVar1S14S104P019P067N047P069: std_logic_vector(   0 downto 0);
        signal cVar1S15S104P019P067N047P069: std_logic_vector(   0 downto 0);
        signal cVar1S16S104P019P067N047P069: std_logic_vector(   0 downto 0);
        signal cVar1S17S104P019P067P024P042nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S104P019P067P024N042: std_logic_vector(   0 downto 0);
        signal cVar1S19S104P019P067P024P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S105P045P030P035P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S105P045P030P035N025: std_logic_vector(   0 downto 0);
        signal cVar1S2S105P045P030P035N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S105N045P029P059P028: std_logic_vector(   0 downto 0);
        signal cVar1S4S105N045P029P059P028: std_logic_vector(   0 downto 0);
        signal cVar1S5S105N045N029P043P062: std_logic_vector(   0 downto 0);
        signal cVar1S6S105N045N029P043P062: std_logic_vector(   0 downto 0);
        signal cVar1S7S105N045N029P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S8S105N045N029P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S9S105N045N029P043N062: std_logic_vector(   0 downto 0);
        signal cVar1S10S105N045N029P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S105N045N029P043N022: std_logic_vector(   0 downto 0);
        signal cVar1S0S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S1S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S2S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S3S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S106P020P039P041P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S106P020P039P041P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S106P020P039P012P060: std_logic_vector(   0 downto 0);
        signal cVar1S9S106P020P039P012P060: std_logic_vector(   0 downto 0);
        signal cVar1S10S106P020P039P012P060: std_logic_vector(   0 downto 0);
        signal cVar1S11S106P020P039P041nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S106P020N039P000P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S106P020N039P000P017: std_logic_vector(   0 downto 0);
        signal cVar1S14S106P020N039P000N017: std_logic_vector(   0 downto 0);
        signal cVar1S0S107P051P041P024P053: std_logic_vector(   0 downto 0);
        signal cVar1S1S107P051P041P024N053: std_logic_vector(   0 downto 0);
        signal cVar1S2S107P051P041P024N053: std_logic_vector(   0 downto 0);
        signal cVar1S3S107P051P041P024P067: std_logic_vector(   0 downto 0);
        signal cVar1S4S107N051P053P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S5S107N051P053P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S6S107N051P053P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S7S107N051P053P007N025: std_logic_vector(   0 downto 0);
        signal cVar1S8S107N051P053N007P048: std_logic_vector(   0 downto 0);
        signal cVar1S9S107N051P053N007P048: std_logic_vector(   0 downto 0);
        signal cVar1S10S107N051P053N007P048: std_logic_vector(   0 downto 0);
        signal cVar1S11S107N051P053P027P030: std_logic_vector(   0 downto 0);
        signal cVar1S0S108P061P059P051P039: std_logic_vector(   0 downto 0);
        signal cVar1S1S108P061P059P051P039: std_logic_vector(   0 downto 0);
        signal cVar1S2S108P061P059N051P045: std_logic_vector(   0 downto 0);
        signal cVar1S3S108P061P059N051P045: std_logic_vector(   0 downto 0);
        signal cVar1S4S108P061P059N051P045: std_logic_vector(   0 downto 0);
        signal cVar1S5S108P061P059N051N045: std_logic_vector(   0 downto 0);
        signal cVar1S6S108P061P059N051N045: std_logic_vector(   0 downto 0);
        signal cVar1S7S108P061P059N051N045: std_logic_vector(   0 downto 0);
        signal cVar1S8S108P061P059N051N045: std_logic_vector(   0 downto 0);
        signal cVar1S9S108P061P059P052P062: std_logic_vector(   0 downto 0);
        signal cVar1S10S108P061P059P052P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S108P061P059P052P062: std_logic_vector(   0 downto 0);
        signal cVar1S12S108P061P040P033P015: std_logic_vector(   0 downto 0);
        signal cVar1S13S108P061P040P033N015: std_logic_vector(   0 downto 0);
        signal cVar1S14S108P061P040N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S15S108P061P040N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S16S108P061P040N033P041: std_logic_vector(   0 downto 0);
        signal cVar1S0S109P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S109P022N043P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S109P022N043N002P003: std_logic_vector(   0 downto 0);
        signal cVar1S3S109N022P043P000P056: std_logic_vector(   0 downto 0);
        signal cVar1S4S109N022P043P000P056: std_logic_vector(   0 downto 0);
        signal cVar1S5S109N022P043P000N056: std_logic_vector(   0 downto 0);
        signal cVar1S6S109N022P043P000N056: std_logic_vector(   0 downto 0);
        signal cVar1S7S109N022P043P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S8S109N022P043N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S9S109N022P043N025P050: std_logic_vector(   0 downto 0);
        signal cVar1S0S110P000P051P041P053: std_logic_vector(   0 downto 0);
        signal cVar1S1S110P000P051P041P053: std_logic_vector(   0 downto 0);
        signal cVar1S2S110P000P051P041P053: std_logic_vector(   0 downto 0);
        signal cVar1S3S110P000P051P041N053: std_logic_vector(   0 downto 0);
        signal cVar1S4S110P000P051P041N053: std_logic_vector(   0 downto 0);
        signal cVar1S5S110P000N051P053P044: std_logic_vector(   0 downto 0);
        signal cVar1S6S110P000N051P053P044: std_logic_vector(   0 downto 0);
        signal cVar1S7S110P000N051P053N044: std_logic_vector(   0 downto 0);
        signal cVar1S8S110P000N051P053N044: std_logic_vector(   0 downto 0);
        signal cVar1S9S110P000N051P053N044: std_logic_vector(   0 downto 0);
        signal cVar1S10S110P000N051P053P030: std_logic_vector(   0 downto 0);
        signal cVar1S11S110P000P030P027P060: std_logic_vector(   0 downto 0);
        signal cVar1S0S111P053P004P051P000: std_logic_vector(   0 downto 0);
        signal cVar1S1S111P053P004P051P000: std_logic_vector(   0 downto 0);
        signal cVar1S2S111P053P004P051P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S111P053P004N051P030: std_logic_vector(   0 downto 0);
        signal cVar1S4S111P053P004N051P030: std_logic_vector(   0 downto 0);
        signal cVar1S5S111N053P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S6S111N053P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S7S111N053P044N025N023: std_logic_vector(   0 downto 0);
        signal cVar1S8S111N053N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S9S111N053N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S10S111N053N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S11S111N053N044P042P023: std_logic_vector(   0 downto 0);
        signal cVar1S12S111N053N044P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S111N053N044P042N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S112P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S112P044N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S112P044N023N025P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S112P044N023N025P032: std_logic_vector(   0 downto 0);
        signal cVar1S4S112N044P042P023P051: std_logic_vector(   0 downto 0);
        signal cVar1S5S112N044P042P023P051: std_logic_vector(   0 downto 0);
        signal cVar1S6S112N044P042P023N051: std_logic_vector(   0 downto 0);
        signal cVar1S7S112N044P042P023N051: std_logic_vector(   0 downto 0);
        signal cVar1S8S112N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S112N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S112N044P042P024P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S112N044P042P024P062: std_logic_vector(   0 downto 0);
        signal cVar1S0S113P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S113P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S113P044N025N023P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S113N044P042P023P051: std_logic_vector(   0 downto 0);
        signal cVar1S4S113N044P042P023P051: std_logic_vector(   0 downto 0);
        signal cVar1S5S113N044P042P023N051: std_logic_vector(   0 downto 0);
        signal cVar1S6S113N044P042P023N051: std_logic_vector(   0 downto 0);
        signal cVar1S7S113N044P042P023N051: std_logic_vector(   0 downto 0);
        signal cVar1S8S113N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S113N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S113N044P042P024P062: std_logic_vector(   0 downto 0);
        signal cVar1S11S113N044P042P024P062: std_logic_vector(   0 downto 0);
        signal cVar1S0S114P016P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S114P016P044N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S114P016P044N023N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S114P016N044P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S114P016N044P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S5S114P016N044N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S6S114P016N044N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S7S114P016N044N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S8S114P016N044N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S9S114P016N044N041P020: std_logic_vector(   0 downto 0);
        signal cVar1S10S114P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S11S114P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S12S114P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S13S114P016P039P022P041: std_logic_vector(   0 downto 0);
        signal cVar1S14S114P016P039P022P019: std_logic_vector(   0 downto 0);
        signal cVar1S15S114P016P039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S114P016P039N005P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S115P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S115P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S115P044N025N023P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S115N044P042P023P008: std_logic_vector(   0 downto 0);
        signal cVar1S4S115N044P042P023P008: std_logic_vector(   0 downto 0);
        signal cVar1S5S115N044P042P023P008: std_logic_vector(   0 downto 0);
        signal cVar1S6S115N044P042P023N008: std_logic_vector(   0 downto 0);
        signal cVar1S7S115N044P042P023N008: std_logic_vector(   0 downto 0);
        signal cVar1S8S115N044P042P023N008: std_logic_vector(   0 downto 0);
        signal cVar1S9S115N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S115N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S115N044P042P023P024: std_logic_vector(   0 downto 0);
        signal cVar1S12S115N044P042P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S115N044P042P024N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S116P016P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S116P016P044N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S116P016P044N023N025: std_logic_vector(   0 downto 0);
        signal cVar1S3S116P016N044P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar1S4S116P016N044P041N020: std_logic_vector(   0 downto 0);
        signal cVar1S5S116P016N044N041P004: std_logic_vector(   0 downto 0);
        signal cVar1S6S116P016N044N041P004: std_logic_vector(   0 downto 0);
        signal cVar1S7S116P016N044N041P004: std_logic_vector(   0 downto 0);
        signal cVar1S8S116P016N044N041P004: std_logic_vector(   0 downto 0);
        signal cVar1S9S116P016N044N041P004: std_logic_vector(   0 downto 0);
        signal cVar1S10S116P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S11S116P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S12S116P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S13S116P016P039P041P022: std_logic_vector(   0 downto 0);
        signal cVar1S14S116P016P039P041P069: std_logic_vector(   0 downto 0);
        signal cVar1S15S116P016P039P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S16S116P016P039N005P069: std_logic_vector(   0 downto 0);
        signal cVar1S0S117P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S117P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S117P044N025N023P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S117N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S117N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S117N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S117N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S117N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S8S117N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S117N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S117N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S117N044P023P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S117N044P023P024N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S118P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S118P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S118P044N025N023P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S118N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S4S118N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S5S118N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S6S118N044P023P042P002: std_logic_vector(   0 downto 0);
        signal cVar1S7S118N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S118N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S9S118N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S118N044P023P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S11S118N044P023P024N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S119P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S119P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S119P044N025N023P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S119N044P023P042P053: std_logic_vector(   0 downto 0);
        signal cVar1S4S119N044P023P042N053: std_logic_vector(   0 downto 0);
        signal cVar1S5S119N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S6S119N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S7S119N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S119N044P023P024P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S119N044P023P024N008: std_logic_vector(   0 downto 0);
        signal cVar1S10S119N044P023P024N008: std_logic_vector(   0 downto 0);
        signal cVar1S0S120P044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S120P044N025P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S120P044N025N023P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S120N044P023P042P054: std_logic_vector(   0 downto 0);
        signal cVar1S4S120N044P023P042P054: std_logic_vector(   0 downto 0);
        signal cVar1S5S120N044P023P042P054: std_logic_vector(   0 downto 0);
        signal cVar1S6S120N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S7S120N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S8S120N044P023P024P005nsss: std_logic_vector(   0 downto 0);
        signal cVar1S9S120N044P023P024N005: std_logic_vector(   0 downto 0);
        signal cVar1S0S121P042P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S121P042N023P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S121P042N023N002P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S121P042N023N002N055: std_logic_vector(   0 downto 0);
        signal cVar1S4S121P042N023N002N055: std_logic_vector(   0 downto 0);
        signal cVar1S5S121N042P023P052P065: std_logic_vector(   0 downto 0);
        signal cVar1S6S121N042P023P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S7S121N042P023P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S8S121N042P023P052N065: std_logic_vector(   0 downto 0);
        signal cVar1S9S121N042P023N052P050: std_logic_vector(   0 downto 0);
        signal cVar1S10S121N042P023N052P050: std_logic_vector(   0 downto 0);
        signal cVar1S11S121N042P023N052P050: std_logic_vector(   0 downto 0);
        signal cVar1S12S121N042P023P024P008nsss: std_logic_vector(   0 downto 0);
        signal cVar1S13S121N042P023P024N008: std_logic_vector(   0 downto 0);
        signal cVar1S14S121N042P023P024N008: std_logic_vector(   0 downto 0);
        signal cVar1S0S122P044P026P025nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S122P044P026N025P000: std_logic_vector(   0 downto 0);
        signal cVar1S2S122P044P026N025P000: std_logic_vector(   0 downto 0);
        signal cVar1S3S122N044P023P042P020: std_logic_vector(   0 downto 0);
        signal cVar1S4S122N044P023P042P020: std_logic_vector(   0 downto 0);
        signal cVar1S5S122N044P023P042P020: std_logic_vector(   0 downto 0);
        signal cVar1S6S122N044P023P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S7S122N044P023P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S8S122N044P023P042N020: std_logic_vector(   0 downto 0);
        signal cVar1S9S122N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S10S122N044P023P042P024: std_logic_vector(   0 downto 0);
        signal cVar1S11S122N044P023P024P006nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S122N044P023P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S13S122N044P023P024N006: std_logic_vector(   0 downto 0);
        signal cVar1S0S123P042P023nsss: std_logic_vector(   0 downto 0);
        signal cVar1S1S123P042N023P002nsss: std_logic_vector(   0 downto 0);
        signal cVar1S2S123P042N023N002P055nsss: std_logic_vector(   0 downto 0);
        signal cVar1S3S123P042N023N002N055: std_logic_vector(   0 downto 0);
        signal cVar1S4S123P042N023N002N055: std_logic_vector(   0 downto 0);
        signal cVar1S5S123N042P023P019P006: std_logic_vector(   0 downto 0);
        signal cVar1S6S123N042P023P019P006: std_logic_vector(   0 downto 0);
        signal cVar1S7S123N042P023P019P006: std_logic_vector(   0 downto 0);
        signal cVar1S8S123N042P023P019P006: std_logic_vector(   0 downto 0);
        signal cVar1S9S123N042P023N019P069: std_logic_vector(   0 downto 0);
        signal cVar1S10S123N042P023N019P069: std_logic_vector(   0 downto 0);
        signal cVar1S11S123N042P023N019N069: std_logic_vector(   0 downto 0);
        signal cVar1S12S123N042P023N019N069: std_logic_vector(   0 downto 0);
        signal cVar1S13S123N042P023N019N069: std_logic_vector(   0 downto 0);
        signal cVar1S14S123N042P023P024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar1S15S123N042P023P024N007: std_logic_vector(   0 downto 0);
        signal cVar1S0S124P019P018P067P039: std_logic_vector(   0 downto 0);
        signal cVar1S1S124P019P018P067P039: std_logic_vector(   0 downto 0);
        signal cVar1S2S124P019P018P067P039: std_logic_vector(   0 downto 0);
        signal cVar1S3S124P019P018P067N039: std_logic_vector(   0 downto 0);
        signal cVar1S4S124P019P018P067N039: std_logic_vector(   0 downto 0);
        signal cVar1S5S124P019P018P067N039: std_logic_vector(   0 downto 0);
        signal cVar1S6S124P019P018P067P028: std_logic_vector(   0 downto 0);
        signal cVar1S7S124P019P018P067P028: std_logic_vector(   0 downto 0);
        signal cVar1S8S124P019P018P039P033: std_logic_vector(   0 downto 0);
        signal cVar1S9S124P019P018P039P033: std_logic_vector(   0 downto 0);
        signal cVar1S10S124P019P018P039N033: std_logic_vector(   0 downto 0);
        signal cVar1S11S124P019P018P039N033: std_logic_vector(   0 downto 0);
        signal cVar1S12S124P019P018P039P017: std_logic_vector(   0 downto 0);
        signal cVar1S13S124P019P051P042P067nsss: std_logic_vector(   0 downto 0);
        signal cVar1S14S124P019P051P042N067: std_logic_vector(   0 downto 0);
        signal cVar1S15S124P019P051P042N067: std_logic_vector(   0 downto 0);
        signal cVar1S16S124P019P051N042P029: std_logic_vector(   0 downto 0);
        signal cVar1S17S124P019P051N042P029: std_logic_vector(   0 downto 0);
        signal cVar1S18S124P019P051N042P029: std_logic_vector(   0 downto 0);
        signal cVar1S19S124P019P051N042P029: std_logic_vector(   0 downto 0);
        signal cVar1S20S124P019P051P037P024: std_logic_vector(   0 downto 0);
        signal cVar1S21S124P019P051P037P024: std_logic_vector(   0 downto 0);
        signal cVar1S22S124P019P051N037P000: std_logic_vector(   0 downto 0);
        signal cVar1S23S124P019P051N037P000: std_logic_vector(   0 downto 0);
        signal cVar1S0S125P018P050P029P032: std_logic_vector(   0 downto 0);
        signal cVar1S1S125P018P050P029P032: std_logic_vector(   0 downto 0);
        signal cVar1S2S125P018P050P029P032: std_logic_vector(   0 downto 0);
        signal cVar1S3S125P018P050P029P032: std_logic_vector(   0 downto 0);
        signal cVar1S4S125P018P050P029P032: std_logic_vector(   0 downto 0);
        signal cVar1S5S125P018P050P029P011: std_logic_vector(   0 downto 0);
        signal cVar1S6S125P018P050P029N011: std_logic_vector(   0 downto 0);
        signal cVar1S7S125P018P050P004P012: std_logic_vector(   0 downto 0);
        signal cVar1S8S125P018P050P004P012: std_logic_vector(   0 downto 0);
        signal cVar1S9S125P018P050P004P012: std_logic_vector(   0 downto 0);
        signal cVar1S10S125N018P039P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S11S125N018P039P054P034: std_logic_vector(   0 downto 0);
        signal cVar1S12S125N018N039P014P060: std_logic_vector(   0 downto 0);
        signal cVar1S13S125N018N039P014P060: std_logic_vector(   0 downto 0);
        signal cVar1S14S125N018N039P014P060: std_logic_vector(   0 downto 0);
        signal cVar1S15S125N018N039P014N060: std_logic_vector(   0 downto 0);
        signal cVar1S16S125N018N039P014N060: std_logic_vector(   0 downto 0);
        signal cVar1S17S125N018N039N014P044: std_logic_vector(   0 downto 0);
        signal cVar1S18S125N018N039N014N044: std_logic_vector(   0 downto 0);
        signal cVar1S19S125N018N039N014N044: std_logic_vector(   0 downto 0);
        signal cVar1S20S125N018N039N014N044: std_logic_vector(   0 downto 0);
        signal cVar1S0S126P018P014P037P004: std_logic_vector(   0 downto 0);
        signal cVar1S1S126P018P014P037P004: std_logic_vector(   0 downto 0);
        signal cVar1S2S126P018P014P037P004: std_logic_vector(   0 downto 0);
        signal cVar1S3S126P018P014P037N004: std_logic_vector(   0 downto 0);
        signal cVar1S4S126P018P014P037N004: std_logic_vector(   0 downto 0);
        signal cVar1S5S126P018P014P037N004: std_logic_vector(   0 downto 0);
        signal cVar1S6S126P018P014P037N004: std_logic_vector(   0 downto 0);
        signal cVar1S7S126P018P014P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S8S126P018P014P037P016: std_logic_vector(   0 downto 0);
        signal cVar1S9S126P018P014P037N016: std_logic_vector(   0 downto 0);
        signal cVar1S10S126P018P014P037N016: std_logic_vector(   0 downto 0);
        signal cVar1S11S126P018P014P060P032nsss: std_logic_vector(   0 downto 0);
        signal cVar1S12S126P018P014P060N032: std_logic_vector(   0 downto 0);
        signal cVar1S13S126P018P014P060N032: std_logic_vector(   0 downto 0);
        signal cVar1S14S126P018P014P060N032: std_logic_vector(   0 downto 0);
        signal cVar1S15S126P018P014N060P044: std_logic_vector(   0 downto 0);
        signal cVar1S16S126P018P061P033nsss: std_logic_vector(   0 downto 0);
        signal cVar1S17S126P018P061N033P048: std_logic_vector(   0 downto 0);
        signal cVar1S18S126P018P061N033P048: std_logic_vector(   0 downto 0);
        signal cVar1S19S126P018P061N033P048: std_logic_vector(   0 downto 0);
        signal cVar1S20S126P018N061P042P063nsss: std_logic_vector(   0 downto 0);
        signal cVar1S21S126P018N061P042N063: std_logic_vector(   0 downto 0);
        signal cVar1S22S126P018N061P042N063: std_logic_vector(   0 downto 0);
        signal cVar1S23S126P018N061N042P050: std_logic_vector(   0 downto 0);
        signal cVar1S24S126P018N061N042P050: std_logic_vector(   0 downto 0);
        signal cVar1S25S126P018N061N042P050: std_logic_vector(   0 downto 0);
        signal cVar1S0S127P017P015P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S1S127P017P015P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S2S127P017P015P014P010: std_logic_vector(   0 downto 0);
        signal cVar1S3S127P017P015P014N010: std_logic_vector(   0 downto 0);
        signal cVar1S4S127P017P015P014N010: std_logic_vector(   0 downto 0);
        signal cVar1S5S127P017P015P014N010: std_logic_vector(   0 downto 0);
        signal cVar1S6S127P017P015P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S7S127P017P015P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S8S127P017P015P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S9S127P017P015P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S10S127P017P015P014P066: std_logic_vector(   0 downto 0);
        signal cVar1S11S127P017P015P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S12S127P017P015P000P019: std_logic_vector(   0 downto 0);
        signal cVar1S13S127P017P015P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S14S127P017P015P000N019: std_logic_vector(   0 downto 0);
        signal cVar1S15S127P017P015P000P008: std_logic_vector(   0 downto 0);
        signal cVar1S16S127P017P015P000P008: std_logic_vector(   0 downto 0);
        signal cVar1S17S127N017P018P027P014nsss: std_logic_vector(   0 downto 0);
        signal cVar1S18S127N017P018N027P002: std_logic_vector(   0 downto 0);
        signal cVar1S19S127N017P018N027P002: std_logic_vector(   0 downto 0);
        signal cVar1S20S127N017P018N027N002: std_logic_vector(   0 downto 0);
        signal cVar1S21S127N017P018N027N002: std_logic_vector(   0 downto 0);
        signal cVar1S22S127N017P018N027N002: std_logic_vector(   0 downto 0);
        signal cVar1S23S127N017N018P067P045: std_logic_vector(   0 downto 0);
        signal cVar1S24S127N017N018P067P045: std_logic_vector(   0 downto 0);
        signal cVar1S25S127N017N018P067P045: std_logic_vector(   0 downto 0);
        signal cVar1S26S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar1S27S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar1S28S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar1S29S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar1S30S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar1S31S127N017N018N067P009: std_logic_vector(   0 downto 0);
        signal cVar2S0S0P014P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S0P014P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S0P063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S0P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S0N030P057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S0P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S0P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S0P067P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S0N067P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S0N067N061P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S0P037P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S0N037P034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S0P069P056P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S0P060P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S0P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S0N032P033P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S0P065P063P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S0N065P056P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S1P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S1P014P024P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S1P014P017P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S1P014P017P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S1P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S1P008P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S1N008P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S1P002P000P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S1P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S1P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S1N069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S1N069N012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S1P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S1N060P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S1N060N037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S1P036P017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S1P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S1N028P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S1N028N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S1P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S1N029P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S1N029N027P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S1P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S1N042P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S1N042N064P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S2P036P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S2P036N045P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S2P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S2P065P033P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S2P065N033psss: std_logic_vector(   0 downto 0);
        signal cVar2S7S2P065P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S2P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S2N046P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S2N046N040P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S2P034P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S2N034P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S2P019P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S2P019N067P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S2P019P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S2P011P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S2P011N058P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S2P065P062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S2P065N062P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S2P067P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S2N067P060P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S2N067N060P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S2P044P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S2P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S3P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S3P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S3N028P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S3N028N026P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S3P033P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S3N033psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S3P010P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S3P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S3P046N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S3N046P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S3N046N028P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S3P024P067P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S3P024N067P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S3P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S4P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S4P004P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S4P062P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S4P062N052P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S4P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S4P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S4N028P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S4P059P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S4P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S4N043P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S4N043N024P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S4P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S4N027P056P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S4N027N056psss: std_logic_vector(   0 downto 0);
        signal cVar2S14S4P018P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S4P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S4P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S4P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S4N053P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S4N053N035P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S4P010P035P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S4P010N035P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S4P010P036P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S5P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S5N029P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S5N029N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S5P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S5N052P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S5N052N015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S5P004P055P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S5P004N055psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S5P004P066P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S5P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S5N057P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S5P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S5N043P047P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S5P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S5N048P056P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S5N048N056P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S5P062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S5P069P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S6P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S6P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S6N009P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S6P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S6P026P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S6P026N031P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S6P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S6N051P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S6P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S6P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S6P012P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S6P012N015P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S7P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S7P026N008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S7N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S7P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S7P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S7P068P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S7P002P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S7P002N057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S7P018P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S7P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S7N024P019P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S7P058P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S7P058P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S7N058P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S7P023P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S7P023N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S7N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S8P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S8N026P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S8N026N029P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S8P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S8N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S8N027N024P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S8P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S8N015P041P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S8N015N041psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S8P069P015P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S8P069P015P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S8P024P018P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S8P024P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S8P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S8N029P062P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S8N029N062psss: std_logic_vector(   0 downto 0);
        signal cVar2S18S8P017P066P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S8N017P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S8P018P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S9P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S9N026P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S9P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S9N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S9N027N024P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S9P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S9N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S9N020N021P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S9P065P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S9P053P028P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S9P053N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S9N053P015P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S9N053N015P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S9P012P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S10P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S10N029P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S10N029N026P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S10P014P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S10P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S10N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S10N020N021P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S10P069P016P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S10P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S10N046P002P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S10N046P002P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S10P050P008P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S10P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S10N056P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S10N056N057P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S10P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S10P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S10N063P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S10N063N066P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S10P014P015P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S10P014P015P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S10N014P066P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S10P057P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S11P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S11P026N008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S11N026P009P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S11P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S11P008P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S11P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S11N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S11N025N027P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S11P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S11P030N057P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S11N030P052P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S11N030N052P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S11P007P012P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S12P024P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S12P024N068P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S12P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S12P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S12N034P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S12P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S12P065P067P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S12P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S12N020P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S12P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S12N027P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S12N027P034P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S12P034P014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S12P034N014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S12N034P017P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S12P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S12N061P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S12P051P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S12P051P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S12P060P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S12P060N053P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S12P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S12N058P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S12P017P058P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S13P064P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S13P064N062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S13N064P003P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S13P008P060P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S13P018P067P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S13P018N067P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S13N018P019P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S13P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S13N050P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S13P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S13N048P054P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S13P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S13N029P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S13N029N028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S13P055P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S13P055N030P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S13N055P041P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S13N055N041P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S13P018P009P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S13N018P003P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S14P011P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S14P050P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S14P050P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S14P003P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S14N003P009P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S14N003N009P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S14P003P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S14P003N009P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S14P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S14N043P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S14N043N042P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S14P056P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S14P056N029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S14N056P047P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S14N056N047P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S14P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S14N061P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S14P050P035P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S14P050N035P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S14P033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S14P033N061P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S14N033P035P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S14P068P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S14N068P017P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S15P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S15N047P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S15N047P016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S15P035P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S15P000P063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S15P000N063P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S15P035P051P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S15N035P036P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S15N035N036P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S15P022P008P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S15P022P008P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S15P057P068P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S15P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S15N029P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S15P047P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S15N047P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S15N047N041P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S15P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S16P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S16P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S16N043P014P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S16P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S16P042N040P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S16P060P056P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S16P011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S16P011P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S16P011P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S16P000P065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S16P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S16P003P066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S16N003P009P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S16N003N009P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S16P045P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S16P045N035P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S16P024P057P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S16P036P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S17P062P022P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S17P024P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S17P024N028P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S17P062P017P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S17P011P033P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S17P011N033P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S17P011P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S17P022P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S17P022N004P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S17N022P043P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S17N022P043P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S17P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S17N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S18P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S18N032P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S18N032N033P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S18P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S18P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S18N047P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S18P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S18N040P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S18P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S18P020N039P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S18N020P039P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S18P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S18N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S18N051N052P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S18P003P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S18P003N028P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S18P003P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S18P008P015P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S19P067P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S19P067N006P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S19P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S19P011N013P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S19P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S19N039P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S19N039N040P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S19P039P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S19P060P018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S20P067P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S20P000P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S20P054P035P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S20P054N035psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S20P054P052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S20P006P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S20P006N039P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S20P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S20N060P034P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S20P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S20N064P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S20P059P069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S20P059P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S20P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S21P067P015P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S21P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S21P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S21N026P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S21N026N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S21P056P039P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S21N056P052P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S21P032P043P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S21P051P018P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S22P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S22N050P009P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S22P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S22P050P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S22P050N029P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S22P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S22N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S22P024P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S22P024N029P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S22P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S22P016P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S22P016N035P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S23P062P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S23P062N009P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S23P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S23N045P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S23P062P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S23N062P063P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S23P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S23P022N043P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S23N022P043P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S23P066P036P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S23P066N036P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S23P014P064P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S23P066P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S24P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S24N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S24N030N031P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S24P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S24P013N016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S24P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S24N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S24N020N021P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S24P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S24P055P004P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S24P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S24N050P062P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S24P068P065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S24P068N065P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S24N068P036P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S24N068P036P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S25P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S25P014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S25P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S25P004P010P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S25P004N010P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S25P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S25N021P008P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S25P028P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S25N028P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S25N028N029P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S25P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S25P040N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S25P061P069P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S26P062P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S26P062N064P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S26N062P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S26N062N067P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S26P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S26P067P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S26N067P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S26N067N026P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S26P024P020P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S26P024P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S26P035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S26N035P066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S26N035N066P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S26P018P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S26P018N015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S26N018P016P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S26P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S26N018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S26P006P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S26P009P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S26P009N055P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S26P009P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S26P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S26P062N035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S26P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S26P015P066P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S26P015P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S26P051P002P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S26P003P068P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S26P011P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S26N011P069P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S27P045P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S27P019P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S27P019N018P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S27P019P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S27P000P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S27P000P007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S27P062P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S27P062P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S27N062P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S27N062N007P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S27P008P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S27P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S27N048P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S27N048N009P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S27P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S27P029N011P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S27N029P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S27N029N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S27P055P065P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S27P067P020P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S28P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S28N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S28N023N022P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S28P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S28P042P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S28P067P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S28N067P062P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S28P009P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S28P009N034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S28P035P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S28P063P037P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S28P063P037P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S28P063P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S28P044P012P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S28P044N012P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S28P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S28N065P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S28P000P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S28P013P063P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S28P013N063P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S28P013P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S28P014P051P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S28P014P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S28P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S28N065P069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S28P011P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S28P011N036P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S29P034P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S29P034P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S29P063P034P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S29P063N034P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S29N063P065P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S29P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S29P020P016P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S29P018P069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S29P007P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S29P030P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S29P030P068P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S29N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S29N030N031P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S29P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S29P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S29N020P061P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S29P036P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S29P036P016P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S30P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S30N023P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S30N023N022P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S30P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S30N020P059P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S30P064P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S30P064N062P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S30N064P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S30P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S30N031P062P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S30P052P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S30N052P062P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S30P014P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S30P005P011P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S30P005P011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S30P011P002P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S30N011P026P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S30N011N026P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S30P034P008P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S30P046P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S31P014P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S31P034P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S31P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S31P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S31P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S31N052P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S31N052N008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S31P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S31N021P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S31N021N002P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S31P038P044P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S31P038P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S31P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S31P064P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S31P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S31N069P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S31P034P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S31P063P014P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S32P068P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S32N068P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S32N068N055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S32P062P041P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S32P062N041psss: std_logic_vector(   0 downto 0);
        signal cVar2S6S32P035P034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S32N035P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S32P013P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S32N013P067P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S32P034P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S32P016P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S32P033P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S32N033P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S32N033N034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S32P013P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S32P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S32P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S32N064P068P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S32P008P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S32P008N015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S32P011P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S33P005P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S33P035P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S33N035P001P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S33P015P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S33P030P019P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S33P030P019P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S33P006P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S33P051P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S33P051N021P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S33P032P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S33P032N015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S33P063P034P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S33P063P034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S33P063P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S33P011P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S33P011N029P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S33N011P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S33P008P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S34P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S34P005P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S34P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S34P069P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S34N069P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S34N069P032P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S34P061P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S34P061N004P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S34P061P018P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S34P033P010P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S34P033N010P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S34P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S34P003P015P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S34P003N015P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S34P003P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S34P021P007P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S34P069P006P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S35P063P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S35P063N066P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S35P063P035P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S35P002P056P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S35P043P063P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S35P068P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S35N068P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S35N068N055P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S35P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S35P063P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S35P063P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S35N063P065P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S35P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S35P020N039P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S35N020P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S35N020N011P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S35P008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S35N008P062P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S35N008P062P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S35P065P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S36P060P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S36P060P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S36P060P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S36P016P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S36P016N067P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S36P016P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S36P034P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S36P034P029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S36P034P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S36P034N029P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S36P064P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S36N064P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S36P004P024P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S36P013P041P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S36N013P031P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S36N013P031P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S36P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S36N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S36P021P039P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S36P000P065P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S36P003P008P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S37P045P053P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S37P045N053P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S37P045P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S37P036P054P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S37P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S37N010P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S37P050P060P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S37P050P060P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S37P010P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S37P024P069P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S37P062P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S37P062N052P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S37N062P063P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S37P045P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S37P045N005P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S37N045P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S38P069P060P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S38P069N060psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S38P069P067P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S38P067P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S38P067P035P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S38N067P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S38N067P032P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S38P000P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S38P051P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S38P051P014P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S38P049P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S38P049N000P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S38P026P015P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S38P011P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S38P005P000P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S38P005P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S38P017P010P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S38P068P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S39P065P068P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S39P065P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S39N065P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S39N065P063P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S39P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S39P035P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S39P022P068P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S39P022P068P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S39P022P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S39P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S39P069P060P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S39P069N060psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S39P032P037P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S39P032P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S39P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S39N047P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S39P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S39P014P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S39P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S40P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S40N056P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S40N056P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S40P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S40N010P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S40N010N057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S40P055P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S40P055N027psss: std_logic_vector(   0 downto 0);
        signal cVar2S8S40P055P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S40P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S40N031P000P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S40P036P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S40P036N037P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S40P018P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S40P018N013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S40P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S40P008P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S40P008N060P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S40P069P035P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S40P069P037P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S40P069N037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S40P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S40P003P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S41P014P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S41P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S41N043P017P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S41P043P056P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S41P043N056P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S41P043P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S41P043N005P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S41P004P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S41P004P012P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S41P059P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S41P059N056P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S41N059P012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S41N059N012P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S41P009P008P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S41P012P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S41N012P009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S41P034P022P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S41P034P037P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S41P065P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S42P027P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S42P027N050P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S42N027P049P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S42N027P049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S42P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S42N040P010P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S42P033P007P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S42P067P058P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S42P067P066P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S42P067P066P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S42P066P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S42P066N035P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S42P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S42P065P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S42P065P018P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S42P065N018P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S42P013P019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S42P013P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S42P013P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S42P065P018P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S42P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S43P009P032P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S43P009N032psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S43P009P004P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S43P008P002P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S43P008P018P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S43P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S43P057P063P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S43P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S43N049P035P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S43P018P011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S43P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S43N010P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S43N010N057P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S43P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S43N021P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S43N021N020P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S43P038P002P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S44P005P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S44P014P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S44N014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S44N014P032P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S44P067P032P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S44P067N032P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S44P067P012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S44P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S44N031P061P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S44N031N061P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S44P000P036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S44N000P068P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S44N000N068P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S44P031P065P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S44P031P065P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S44P031P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S44P008P004P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S44P057P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S44P063P016P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S44P063N016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S44P006P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S44P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S45P000P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S45P000N016P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S45N000P069P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S45N000P069P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S45P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S45N064P069P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S45N057P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S45P034P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S45P034N064P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S45N034psss: std_logic_vector(   0 downto 0);
        signal cVar2S11S45P064P029P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S45P064P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S45P014P017P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S45P014N017P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S45N014P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S45N014N027P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S45P025P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S45P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S45P057P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S45P053P063P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S45P006P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S45P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S46P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S46P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S46N031P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S46P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S46N023P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S46P060P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S46P060N062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S46N060P007P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S46N060N007P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S46P049P033P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S46P049P051P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S46P014P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S46P039P010P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S46P069P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S46P069N034P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S46P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S46P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S46N031P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S46P057P008P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S46P057P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S46P037P060P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S46N037P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S47P059P000P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S47N059P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S47P045P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S47P060P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S47P068P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S47P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S47N059P069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S47P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S47P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S47P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S47P010N028P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S47N010P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S47N010N036P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S47P059P061P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S47P059P061P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S47P059P033P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S47P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S47N002P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S47N002N054P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S47P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S47P051P061P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S47P051P053P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S48P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S48N025P009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S48N025N009P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S48P049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S48P049P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S48P049N009P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S48P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S48P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S48N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S48P029P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S48N029P003P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S48P053P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S48P003P064P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S48N003P026P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S48P016P065P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S48P016P067P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S48P034P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S48P034N013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S49P034P032P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S49N034P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S49N034N028psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S49P039P062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S49P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S49P034P053P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S49P017P037P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S49N017P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S49P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S49P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S49P054P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S49P054P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S49P001P033P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S49P001N033P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S49P010P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S49P010N028P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S49N010P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S49N010N036P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S49P030P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S49P030P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S50P037P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S50P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S50N036P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S50N036P013P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S50P004P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S50P011P006P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S50N011P054P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S50N011P054P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S50P065P006P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S50P062P039P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S50P062P064P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S50P034P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S50N034P069P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S50P012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S50P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S50N036P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S51P040P038P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S51P040P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S51P012P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S51P012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S51P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S51N036P008P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S51N036N008P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S51P012P050P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S51N012P050P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S51N012N050P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S51P061P033P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S51P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S51N021P006P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S51P030P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S51P030N046P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S51P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S51P030N057P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S51P057P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S51N057P000P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S51N057N000P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S52P004P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S52P004N048P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S52P048P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S52P048P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S52P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S52P048N025P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S52P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S52P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S52N016P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S52P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S52N058P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S52P030P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S52N030P000P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S52N030N000P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S52P050P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S52P010P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S52N010P009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S52P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S52P017P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S52N017P012P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S52P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S53P010P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S53P010P012P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S53P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S53N026P037P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S53P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S53N008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S53P060P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S53N060P064P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S53P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S53P039P007P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S53P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S53N060P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S53N060N069P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S53P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S53N042P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S53P042P044P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S53P042P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S54P050P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S54P042P065P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S54P042N065psss: std_logic_vector(   0 downto 0);
        signal cVar2S3S54P034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S54P034P037P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S54P035P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S54P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S54N033P011P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S54P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S54N055P062P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S54N055N062P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S54P002P016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S54P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S54P064P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S54P064P011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S54P064P011P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S54P064P058P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S54N064P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S54N064N028P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S54P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S54N031P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S54P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S54N060P064P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S54P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S54P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S55P000P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S55P000N037P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S55N000P004P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S55N000P004P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S55P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S55P006P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S55P006N036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S55P049P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S55P000P036P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S55P006P055P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S55P054P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S55P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S55P041P020P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S55P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S55N008P069P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S55P009P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S55P065P010P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S55N065P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S55N065P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S55P066P024P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S55P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S55N022P016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S55P042P044P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S55P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S55P042N005P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S56P063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S56N063P067P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S56N063N067P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S56P027P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S56P027N009P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S56N027P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S56N027P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S56P050P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S56P000P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S56P000N037P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S56N000P016P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S56P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S56P006P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S56P049P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S56P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S56P016psss: std_logic_vector(   0 downto 0);
        signal cVar2S16S56P064P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S56N064P034P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S56P016P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S56P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S56N050P000P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S57P067P013P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S57P067N013psss: std_logic_vector(   0 downto 0);
        signal cVar2S2S57P067P033P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S57P013P018P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S57P013N018P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S57P013P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S57P013P017P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S57P012P013P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S57P012P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S57P012P016P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S57P066P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S57P006P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S57P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S57P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S57P013P014P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S57P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S57N009P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S57P066P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S57N066P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S57N066N035P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S57P024P002P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S58P004P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S58P004N022P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S58N004P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S58N004P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S58P043P003P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S58P043N003P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S58P043P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S58P019P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S58P019N036P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S58P019P017P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S58P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S58P053P024P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S58N053P051P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S58N053P051P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S58P009P014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S58P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S58P061P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S58P061N033P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S58P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S58P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S58P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S58N014P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S58P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S59P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S59P016P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S59P016N000P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S59P052P062P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S59P052P062P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S59P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S59P024P012P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S59P002P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S59P002P014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S59P063P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S59N063P016P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S59P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S59P003P005P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S59P003P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S59P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S59N020P012P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S59P020P057P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S59P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S59P009P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S59P011P014P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S59P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S60P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S60N028P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S60N028N058P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S60P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S60N004P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S60N004N032P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S60P004P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S60P024P034P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S60P009P007P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S60P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S60N060P014P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S60P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S60P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S60P014P012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S60P014N012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S60P051P065P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S60P051N065P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S60P051P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S60P056P000P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S60P056P034P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S60P061P009P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S60P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S61P061P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S61P061N013P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S61N061P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S61N061N031P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S61P056P007P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S61P014P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S61P014P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S61P015P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S61P015P063P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S61P034P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S61P034N008psss: std_logic_vector(   0 downto 0);
        signal cVar2S12S61P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S61N022P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S61N022N040P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S61P022P028P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S61P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S61P007P069P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S61P007N069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S61P011P014P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S61P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S62P010P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S62N010P030P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S62P026P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S62N026P053P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S62N026P053P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S62P069P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S62P063P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S62N063P036P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S62P045P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S62P045N061P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S62P045P066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S62P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S62P057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S63P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S63P030P006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S63P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S63P012P014P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S63N012P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S63N012N058P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S63P057P054P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S63P057P054P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S63P057P062P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S63P062P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S63P062N069P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S63N062P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S63P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S63P030P056P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S63P030P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S63P068P017P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S63P068P017P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S63P059P057P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S64P010P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S64N010P006P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S64P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S64P041N020P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S64N041P020P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S64N041P020P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S64P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S64P009P012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S64P009N012P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S64P009P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S64P011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S64P036P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S64P064P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S64P064P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S64N064P062P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S64N064P062P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S64P048P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S64N048P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S64N048N029P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S64P055P009P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S64P055N009P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S64P065P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S65P065P006P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S65N065P036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S65N065P036P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S65P016P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S65P016N041P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S65P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S65P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S65N029P005P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S65P055P060P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S65P065P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S65P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S65N057P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S65N057N052P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S65P006P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S65P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S65N020P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S65P036P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S65P020P033P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S65P020P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S65P020N040P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S65P010P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S66P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S66N041P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S66P032P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S66P032N014P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S66N032P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S66P014P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S66P027P034P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S66P043P063P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S66P069P010P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S66P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S66P069P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S67P037P039P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S67N037P069P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S67N037P069P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S67P065P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S67P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S67P053P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S67P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S67N047P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S67P047P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S67P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S67P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S67P008N026P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S67N008P010P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S68P055P065P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S68P055N065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S68N055P057P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S68P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S68P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S68N027P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S68P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S68N000P051P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S68P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S68P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S68N047P013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S68P005P000P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S68P005P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S68P036P011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S68P014P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S69P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S69P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S69P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S69P006P069P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S69P006N069P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S69P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S69N008P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S69P024P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S69N024P047P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S69P056P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S69N056P059P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S69N056N059P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S69P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S70P046P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S70P046N021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S70P046P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S70P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S70N045P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S70N045N024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S70P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S70N047P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S70N047N012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S70P032P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S70P032N003P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S70P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S70P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S70N031P052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S71P060P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S71P030P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S71N030P041P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S71P030P016P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S71P030N016P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S71P030P055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S71P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S71N002P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S71N002N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S71P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S72P019P013P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S72N019P010P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S72P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S72P044N023P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S72N044P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S72P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S72P065P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S72P043P037P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S72P043P065P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S72P019P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S72P010P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S72P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S73P011P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S73P011P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S73P041P030P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S73P041N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S73P030P051P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S73P030P055P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S73P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S73N002P018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S73N002N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S73P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S73N012P018P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S74P010P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S74P010N008P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S74P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S74P066P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S74P013P039P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S74N013P032P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S74P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S74N047P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S74P047P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S74P047P048P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S74P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S74P047N026P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S74P030P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S74P048P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S74P048N062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S74N048P027P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S74P018P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S74P012P003P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S74P012P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S75P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S75P031P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S75N031P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S75N031N029P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S75P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S75P036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S75P036N034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S75P060P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S75P060N034P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S75N060P031P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S75N060P031P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S75P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S75N013P012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S75P068P026P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S75P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S75N046P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S75N046N049P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S75P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S75N047P054P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S75P047P044P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S75P047N044P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S75P047P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S76P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S76N028P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S76P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S76P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S76N046P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S76P052P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S76P052N024P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S76P052P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S76P052N062P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S76P004P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S76P004N008P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S76P043P022P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S76P043P036P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S76P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S76N036P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S76P017P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S76P012P003P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S76P012P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S77P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S77N057P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S77N057N053P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S77P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S77N031P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S77P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S77P036P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S77P036N034P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S77P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S77N024P017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S77P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S77N040P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S77N040P011P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S77P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S77P067P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S77N067P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S77N067N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S78P043P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S78P021P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S78P021N040P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S78N021P038P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S78P022P064P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S78P022P064P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S78P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S78N021P008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S79P057P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S79P043P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S79P043N048P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S79P047P024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S79P047N024P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S79N047P049P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S79N047P049P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S79P018P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S79P018N042P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S79N018P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S79P036P018P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S79P036N018P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S80P062P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S80N062P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S80N062N047P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S80P019P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S80N019P057P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S80N019N057P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S80P017P067P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S80P017N067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S80P017P035P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S80P044P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S80N044P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S80P003P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S80P003P058P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S80P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S80N041P039P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S80P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S80P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S80N014P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S80P014P008P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S80P014P019P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S80P012P051P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S80N012P069P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S81P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S81P053P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S81P053N014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S81N053P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S81N053N035P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S81P016P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S81P063P056P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S81P063P056P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S81P063P024P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S81P012P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S81P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S81N036P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S81P062P063P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S81P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S81N031P013P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S81N031P013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S81P005P067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S81P005P067P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S81P036N016P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S81P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S81N027P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S81N027N025P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S81P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S81N013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S81N013N011P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S81P015P004P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S81P015P004P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S81N015P051P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S82P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S82N002P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S82P021P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S82P021N050P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S82P021P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S82P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S82N002P057P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S82N002N057P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S82P059P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S82P053P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S82P053N014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S82N053P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S82P016P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S82P031P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S82N031P024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S82P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S82P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S83P003P034P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S83P003P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S83P061P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S83P061N033P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S83N061P032P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S83N061N032P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S83P033P009P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S83P033P037P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S83P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S83P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S83N036P069P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S83P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S83P013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S83P013N012P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S83P026P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S83P026P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S83P026P068P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S83P051P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S83P051N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S83N051P053P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S83P014P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S83P014N012P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S84P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S84N064P011P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S84P031P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S84N031P029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S84N031N029P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S84P031P032P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S84P031P032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S84P031P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S84P048P000P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S84P048N000P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S84P048P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S84P018P004P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S84N018P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S84P068P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S84P068P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S84P015P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S84P058P009P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S84P052P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S84N052P063P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S84N052P063P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S84P000P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S85P019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S85N019P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S85P057P035P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S85P057P035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S85P057P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S85P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S85P017P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S85P017N066P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S85P017P015P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S85P017P015P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S85P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S85N031P012P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S85P033P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S85P033N062P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S85N033P010P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S85N033N010P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S85P013P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S85P013N017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S85P061P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S85P061N064P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S85P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S85N025P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S85N025N027P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S85P046P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S86P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S86N027P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S86P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S86N047P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S86P032P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S86P032N056P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S86P032P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S86P009P019P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S86P009N019psss: std_logic_vector(   0 downto 0);
        signal cVar2S10S86P009P016P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S86P019P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S86P019N018P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S86P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S86P019P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S86N019P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S86P057P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S86P057N014P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S86P066P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S86P066P062P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S87P016P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S87P016N064P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S87N016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S87N016N011P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S87P036P010P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S87N036P067P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S87N036N067P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S87P033P045P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S87P033N045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S87P033P012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S87P035P031P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S87P035P032P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S87P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S87P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S87P034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S87N034P006P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S87N034N006P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S87P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S87N020P017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S87N020N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S87P021P068P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S87P021N068P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S87P021P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S87P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S88P007P005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S88N007P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S88N007P012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S88P008P016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S88P008N016P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S88P059P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S88N059P066P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S88P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S88P058P028P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S88P058P028P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S88P058P037P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S88P008P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S88N008P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S88N008N029P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S88P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S88N034P009P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S88P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S88N012P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S88P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S88N069P065P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S89P005P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S89P005P013P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S89P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S89P066P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S89P059P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S89N059P066P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S89P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S89N042P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S89N042N007P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S89P022P045P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S89P022P014P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S89P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S89N022P024P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S89N022N024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S89P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S89P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S89N046P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S89N046N005P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S90P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S90P050P018P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S90P050P018P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S90N050P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S90N050N066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S90P026P010P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S90P026N010P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S90P043P022P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S90P043P022P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S90P043P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S90P043N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S90P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S90P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S90P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S90P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S90N046P016P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S90N046N016P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S91P034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S91P034P016P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S91P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S91N067P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S91N067N066P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S91P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S91N025P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S91P037P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S91P037N062P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S91P037P018P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S91P026P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S91P057P040P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S91P065P001P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S92P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S92N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S92N051N052P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S92P037P007P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S92P037P007P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S92N037P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S92N037N045P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S92P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S92N034P026P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S92P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S92P011P029P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S92P050P061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S92P050N061P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S92P050P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S92P004P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S92P004N006P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S92P015P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S92N015P028P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S92N015N028P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S92P058P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S92N058P067P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S92P036P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S92P036N063P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S92P013P065P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S93P012P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S93P012N036P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S93P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S93P069P065P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S93P069N065P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S93N069P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S93N069N047P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S93P036P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S93P067P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S93P008P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S93N008P017P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S93P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S93P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S93N012P060nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S93P037P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S93P029P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S93P029N028P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S93P007P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S93P007N025P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S93N007P053P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S93P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S93N034P063P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S94P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S94N054P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S94N054N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S94P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S94N034P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S94N034N015P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S94P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S94N005P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S94N005N024P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S94P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S94P022P043P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S94P055P008P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S94P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S94N017P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S94P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S94N042P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S94P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S94P008P063P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S94P008N063P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S94N008P018P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S94P018P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S94P018N030P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S94P018P068P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S95P066P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S95P066P012P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S95P066P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S95P032P004P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S95P032P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S95P009P004P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S95P009N004P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S95P009P017P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S95P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S95N007P010P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S95P017P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S95P060P014P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S95P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S95N007P069P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S95P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S95N054P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S95N054N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S95P055P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S95P055N008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S95P013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S95N013P016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S95N013P016P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S95P054P002P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S95P054N002P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S95P054P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S96P069P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S96P069N024P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S96P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S96N011P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S96N011N034P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S96P040P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S96P040N038P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S96N040P038P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S96P049P064P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S96P049N064P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S96P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S96N017P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S96P060P034P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S96P051P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S96P051N056P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S96P051P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S96P034P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S96P034N037P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S96P064P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S96P064N012P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S96N064P061P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S96P065P031P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S96P065P031P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S96P065P034P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S96P020P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S97P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S97N023P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S97P004P030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S97P004N030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S97P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S97P029P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S97P029N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S97N029P037P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S97N029N037P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S97P014P035P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S97P034P008P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S98P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S98N005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S98P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S98N069P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S98P049P043P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S98P049P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S98P049N026P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S98P027P049P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S98P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S98N012P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S98P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S98P000P012P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S98P000P012P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S98N000P030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S98N000N030P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S98P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S98P067P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S98P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S98P017P014P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S99P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S99N023P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S99P029P067P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S99P029N067P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S99P029P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S99P024P037P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S99P024N037P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S99P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S99N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S99P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S99N054P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S99N054N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S99P055P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S99P055N008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S99P036P013P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S99P036N013P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S99P048P017P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S99N048P031P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S100P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S100N005P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S100P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S100N054P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S100N054N051P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S100P055P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S100P055N034P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S100P053P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S100P053N012P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S100P053P056P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S100P053P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S100N053P006P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S100P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S100N012P066P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S100P018P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S100P018N052P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S100P048P058P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S100P048P016P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S100P020P029P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S101P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S101N022P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S101N022N023P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S101P006P044P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S101P006P044P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S101P006P036P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S101P012P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S101P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S101N017P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S101P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S101N069P028P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S101P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S101N002P021nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S102P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S102P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S102N069P028P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S102P056P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S102P056N053P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S102P056P058P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S102P056N058P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S102P031P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S102P031N068P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S102N031P004P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S102P030P033P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S102P030P033P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S102P030P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S102P008P055P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S102P050P065P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S102N050P024P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S102N050N024P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S102P017P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S102P034P036P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S102P064P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S103P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S103N023P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S103P008P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S103N008P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S103P005P061P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S103P005P008P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S103P039P025P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S103P039P025P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S103P039P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S103P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S103N003P013P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S104P062P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S104P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S104P055P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S104P055N009P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S104P051P011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S104P051N011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S104N051P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S104P009P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S104P009P036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S104P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S104P049P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S104P018P005P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S104N018P054P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S104P014P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S104P014N036P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S104P052nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S104P063P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S105P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S105N022P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S105P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S105N051P000P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S105P052P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S105N052P035P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S105P064P000P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S105P064N000P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S105P064P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S105P050P008P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S106P051P011P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S106P051N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S106N051P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S106N051N045P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S106P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S106N042P007P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S106N042N007P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S106P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S106N003P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S106N003N033P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S106P011P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S106P011N036P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S106P035P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S107P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S107P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S107P069P015P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S107P018P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S107P065P009P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S107P065N009P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S107P065P006P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S107P025P059P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S107P025P010P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S107P037P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S107P016P013P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S108P024nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S108P024P012P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S108P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S108N022P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S108N022N025P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S108P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S108P041N020P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S108N041P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S108N041P043P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S108P057P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S108P057N012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S108N057P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S108P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S108P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S108P059P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S108N059P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S108N059N032P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S109P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S109P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S109N030P013P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S109P054P053P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S109P054P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S109P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S109N023P034P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S110P009P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S110N009P011P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S110N009N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S110P069P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S110P069P015P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S110P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S110N023P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S110P042P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S110P042P023P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S110P042P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S110P064P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S110P056P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S111P011P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S111N011P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S111N011N008P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S111P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S111N064P059P054nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S111P026P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S111P056P004P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S111N056P054P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S111P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S111N045P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S111P009P016P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S112P000P013P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S112P000P013P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S112P041P053P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S112P041N053P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S112P053P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S112P053N041P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S112P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S112N045P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S112P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S112N063P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S113P000P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S113P041P053P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S113P041N053P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S113P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S113P041N020P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S113N041P039P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S113P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S113N045P034P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S113P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S113N063P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S114P026P048P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S114P062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S114P004P008P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S114P004N008P047nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S114P004P003P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S114P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S114N040P064P007nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S114P002P015P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S114P002P066P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S114P002N066P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S114P069P010P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S114P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S114P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S115P000P056P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S115P031P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S115P031P032P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S115P031P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S115P016P022nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S115P016P022P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S115N016P022P043nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S115P006nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S115N006P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S115N006N045P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S115P009P062P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S116P026P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S116P062P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S116P010P028P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S116P010N028P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S116N010P027P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S116N010N027P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S116P003P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S116P002P015P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S116P002P066P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S116P002N066P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S116P019P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S116P010P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S116P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S117P000P056P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S117P005P039P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S117P005P039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S117P005P031P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S117P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S117N038P054P030nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S117P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S117N002P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S117N002N069P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S117P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S118P000P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S118P005P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S118P005P039P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S118P005P031P041nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S118P038nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S118P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S118N002P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S118N002N069P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S118P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S119P032P013P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S119P004P051nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S119P051P041P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S119P002nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S119N002P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S119N002N063P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S119P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S119P069N036P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S120P032P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S120P056P030P057nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S120P056P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S120P056P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S120P062P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S120P062N065P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S120P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S121P006P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S121N006P024P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S121P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S121P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S121N062P050P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S121N062N050P053nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S121P046P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S121N046P025P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S121P004P063P048nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S121P069P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S121P069N036P068nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S122P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S122N023P032P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S122P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S122N039P062P008nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S122N039P062P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S122P039P059P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S122P039N059P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S122P039P012P050nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S122P062P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S122P062N063P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S122P045nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S122N045P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S123P006P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S123N006P024P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S123P067P069nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S123P067P069P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S123P067P024P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S123P046nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S123P045P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S123P045N029P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S123P051P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S123P051N011P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S123N051P038P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S123P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S124P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S124N003P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S124N003N020P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S124P063P058nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S124P063N058P001nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S124N063P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S124P006P021P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S124P006P012P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S124P007P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S124P007P015P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S124P006P066nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S124N006P009P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S124P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S124P037nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S124N037P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S124P013P048P005nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S124P013P048P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S124P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S124N010P067P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S124P061nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S124N061P017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S124P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S124N026P017P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S125P061P033nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S125P061N033P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S125N061P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S125P013P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S125P013P014P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S125P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S125P013nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S125P056P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S125P056N034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S125P016P010nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S125P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S125N020P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S125P032nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S125N032P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S125N032N034P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S125P044P054P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S125P044P054P065nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S125P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S125P042P030P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S125P042N030P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S125P042P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S126P042nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S126N042P013P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S126N042N013P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S126P030P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S126P030N059P031nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S126N030P055P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S126N030P055P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S126P006P062P064nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S126P006N062psss: std_logic_vector(   0 downto 0);
        signal cVar2S9S126P036P006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S126P036N006P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S126P034nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S126N034P016P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S126N034P016P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S126P046P027P017nsss: std_logic_vector(   0 downto 0);
        signal cVar2S17S126P011P067nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S126N011P035P062nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S126N011N035P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S126P010P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S126P010P016P015nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S126P001P009nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S126N001P023P003nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S126P000P049nsss: std_logic_vector(   0 downto 0);
        signal cVar2S0S127P036nsss: std_logic_vector(   0 downto 0);
        signal cVar2S1S127N036P028nsss: std_logic_vector(   0 downto 0);
        signal cVar2S2S127N036N028P035nsss: std_logic_vector(   0 downto 0);
        signal cVar2S3S127P032P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S4S127P032P019P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S5S127N032P023nsss: std_logic_vector(   0 downto 0);
        signal cVar2S6S127P010P032P056nsss: std_logic_vector(   0 downto 0);
        signal cVar2S7S127P010P032P059nsss: std_logic_vector(   0 downto 0);
        signal cVar2S8S127P010P006P019nsss: std_logic_vector(   0 downto 0);
        signal cVar2S9S127P068P013P018nsss: std_logic_vector(   0 downto 0);
        signal cVar2S10S127P068N013P012nsss: std_logic_vector(   0 downto 0);
        signal cVar2S11S127P028P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S12S127P028P016P040nsss: std_logic_vector(   0 downto 0);
        signal cVar2S13S127P061P020nsss: std_logic_vector(   0 downto 0);
        signal cVar2S14S127P061P013P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S15S127P063nsss: std_logic_vector(   0 downto 0);
        signal cVar2S16S127N063P010P016nsss: std_logic_vector(   0 downto 0);
        signal cVar2S18S127P004nsss: std_logic_vector(   0 downto 0);
        signal cVar2S19S127N004P016P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S20S127P050P044nsss: std_logic_vector(   0 downto 0);
        signal cVar2S21S127P050N044P025nsss: std_logic_vector(   0 downto 0);
        signal cVar2S22S127P050P029nsss: std_logic_vector(   0 downto 0);
        signal cVar2S23S127P036P035P039nsss: std_logic_vector(   0 downto 0);
        signal cVar2S24S127P036P035P014nsss: std_logic_vector(   0 downto 0);
        signal cVar2S25S127P036P016P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S26S127P011P055nsss: std_logic_vector(   0 downto 0);
        signal cVar2S27S127P011N055P000nsss: std_logic_vector(   0 downto 0);
        signal cVar2S28S127N011P036P026nsss: std_logic_vector(   0 downto 0);
        signal cVar2S29S127P027nsss: std_logic_vector(   0 downto 0);
        signal cVar2S30S127N027P007P011nsss: std_logic_vector(   0 downto 0);
        signal cVar2S31S127N027N007P065nsss: std_logic_vector(   0 downto 0);
        signal oVar1S0: std_logic_vector(   0 downto 0);
        signal oVar1S1: std_logic_vector(   0 downto 0);
        signal oVar1S2: std_logic_vector(   0 downto 0);
        signal oVar1S3: std_logic_vector(   0 downto 0);
        signal oVar1S4: std_logic_vector(   0 downto 0);
        signal oVar1S5: std_logic_vector(   0 downto 0);
        signal oVar1S6: std_logic_vector(   0 downto 0);
        signal oVar1S7: std_logic_vector(   0 downto 0);
        signal oVar1S8: std_logic_vector(   0 downto 0);
        signal oVar1S9: std_logic_vector(   0 downto 0);
        signal oVar1S10: std_logic_vector(   0 downto 0);
        signal oVar1S11: std_logic_vector(   0 downto 0);
        signal oVar1S12: std_logic_vector(   0 downto 0);
        signal oVar1S13: std_logic_vector(   0 downto 0);
        signal oVar1S14: std_logic_vector(   0 downto 0);
        signal oVar1S15: std_logic_vector(   0 downto 0);
        signal oVar1S16: std_logic_vector(   0 downto 0);
        signal oVar1S17: std_logic_vector(   0 downto 0);
        signal oVar1S18: std_logic_vector(   0 downto 0);
        signal oVar1S19: std_logic_vector(   0 downto 0);
        signal oVar1S20: std_logic_vector(   0 downto 0);
        signal oVar1S21: std_logic_vector(   0 downto 0);
        signal oVar1S22: std_logic_vector(   0 downto 0);
        signal oVar1S23: std_logic_vector(   0 downto 0);
        signal oVar1S24: std_logic_vector(   0 downto 0);
        signal oVar1S25: std_logic_vector(   0 downto 0);
        signal oVar1S26: std_logic_vector(   0 downto 0);
        signal oVar1S27: std_logic_vector(   0 downto 0);
        signal oVar1S28: std_logic_vector(   0 downto 0);
        signal oVar1S29: std_logic_vector(   0 downto 0);
        signal oVar1S30: std_logic_vector(   0 downto 0);
        signal oVar1S31: std_logic_vector(   0 downto 0);
        signal oVar1S32: std_logic_vector(   0 downto 0);
        signal oVar1S33: std_logic_vector(   0 downto 0);
        signal oVar1S34: std_logic_vector(   0 downto 0);
        signal oVar1S35: std_logic_vector(   0 downto 0);
        signal oVar1S36: std_logic_vector(   0 downto 0);
        signal oVar1S37: std_logic_vector(   0 downto 0);
        signal oVar1S38: std_logic_vector(   0 downto 0);
        signal oVar1S39: std_logic_vector(   0 downto 0);
        signal oVar1S40: std_logic_vector(   0 downto 0);
        signal oVar1S41: std_logic_vector(   0 downto 0);
        signal oVar1S42: std_logic_vector(   0 downto 0);
        signal oVar1S43: std_logic_vector(   0 downto 0);
        signal oVar1S44: std_logic_vector(   0 downto 0);
        signal oVar1S45: std_logic_vector(   0 downto 0);
        signal oVar1S47: std_logic_vector(   0 downto 0);
        signal oVar1S48: std_logic_vector(   0 downto 0);
        signal oVar1S49: std_logic_vector(   0 downto 0);
        signal oVar1S50: std_logic_vector(   0 downto 0);
        signal oVar1S51: std_logic_vector(   0 downto 0);
        signal oVar1S52: std_logic_vector(   0 downto 0);
        signal oVar1S53: std_logic_vector(   0 downto 0);
        signal oVar1S54: std_logic_vector(   0 downto 0);
        signal oVar1S55: std_logic_vector(   0 downto 0);
        signal oVar1S56: std_logic_vector(   0 downto 0);
        signal oVar1S57: std_logic_vector(   0 downto 0);
        signal oVar1S58: std_logic_vector(   0 downto 0);
        signal oVar1S59: std_logic_vector(   0 downto 0);
        signal oVar1S60: std_logic_vector(   0 downto 0);
        signal oVar1S61: std_logic_vector(   0 downto 0);
        signal oVar1S62: std_logic_vector(   0 downto 0);
        signal oVar1S63: std_logic_vector(   0 downto 0);
        signal oVar1S65: std_logic_vector(   0 downto 0);
        signal oVar1S66: std_logic_vector(   0 downto 0);
        signal oVar1S67: std_logic_vector(   0 downto 0);
        signal oVar1S68: std_logic_vector(   0 downto 0);
        signal oVar1S69: std_logic_vector(   0 downto 0);
        signal oVar1S70: std_logic_vector(   0 downto 0);
        signal oVar1S71: std_logic_vector(   0 downto 0);
        signal oVar1S72: std_logic_vector(   0 downto 0);
        signal oVar1S73: std_logic_vector(   0 downto 0);
        signal oVar1S74: std_logic_vector(   0 downto 0);
        signal oVar1S75: std_logic_vector(   0 downto 0);
        signal oVar1S77: std_logic_vector(   0 downto 0);
        signal oVar1S78: std_logic_vector(   0 downto 0);
        signal oVar1S79: std_logic_vector(   0 downto 0);
        signal oVar1S80: std_logic_vector(   0 downto 0);
        signal oVar1S81: std_logic_vector(   0 downto 0);
        signal oVar1S83: std_logic_vector(   0 downto 0);
        signal oVar1S84: std_logic_vector(   0 downto 0);
        signal oVar1S85: std_logic_vector(   0 downto 0);
        signal oVar1S86: std_logic_vector(   0 downto 0);
        signal oVar1S87: std_logic_vector(   0 downto 0);
        signal oVar1S88: std_logic_vector(   0 downto 0);
        signal oVar1S89: std_logic_vector(   0 downto 0);
        signal oVar1S90: std_logic_vector(   0 downto 0);
        signal oVar1S91: std_logic_vector(   0 downto 0);
        signal oVar1S92: std_logic_vector(   0 downto 0);
        signal oVar1S93: std_logic_vector(   0 downto 0);
        signal oVar1S94: std_logic_vector(   0 downto 0);
        signal oVar1S96: std_logic_vector(   0 downto 0);
        signal oVar1S97: std_logic_vector(   0 downto 0);
        signal oVar1S98: std_logic_vector(   0 downto 0);
        signal oVar1S99: std_logic_vector(   0 downto 0);
        signal oVar1S100: std_logic_vector(   0 downto 0);
        signal oVar1S101: std_logic_vector(   0 downto 0);
        signal oVar1S102: std_logic_vector(   0 downto 0);
        signal oVar1S103: std_logic_vector(   0 downto 0);
        signal oVar1S104: std_logic_vector(   0 downto 0);
        signal oVar1S106: std_logic_vector(   0 downto 0);
        signal oVar1S107: std_logic_vector(   0 downto 0);
        signal oVar1S108: std_logic_vector(   0 downto 0);
        signal oVar1S109: std_logic_vector(   0 downto 0);
        signal oVar1S110: std_logic_vector(   0 downto 0);
        signal oVar1S112: std_logic_vector(   0 downto 0);
        signal oVar1S113: std_logic_vector(   0 downto 0);
        signal oVar1S114: std_logic_vector(   0 downto 0);
        signal oVar1S115: std_logic_vector(   0 downto 0);
        signal oVar1S116: std_logic_vector(   0 downto 0);
        signal oVar1S117: std_logic_vector(   0 downto 0);
        signal oVar1S118: std_logic_vector(   0 downto 0);
        signal oVar1S120: std_logic_vector(   0 downto 0);
        signal oVar1S121: std_logic_vector(   0 downto 0);
        signal oVar1S122: std_logic_vector(   0 downto 0);
        signal oVar1S123: std_logic_vector(   0 downto 0);
        signal oVar1S124: std_logic_vector(   0 downto 0);
        signal oVar1S125: std_logic_vector(   0 downto 0);
        signal oVar1S126: std_logic_vector(   0 downto 0);
        signal oVar1S127: std_logic_vector(   0 downto 0);
        signal oVar1S128: std_logic_vector(   0 downto 0);
        signal oVar1S129: std_logic_vector(   0 downto 0);
        signal oVar1S130: std_logic_vector(   0 downto 0);
        signal oVar1S131: std_logic_vector(   0 downto 0);
        signal oVar1S132: std_logic_vector(   0 downto 0);
        signal oVar1S133: std_logic_vector(   0 downto 0);
        signal oVar1S134: std_logic_vector(   0 downto 0);
        signal oVar1S135: std_logic_vector(   0 downto 0);
        signal oVar1S136: std_logic_vector(   0 downto 0);
        signal oVar1S137: std_logic_vector(   0 downto 0);
        signal oVar1S138: std_logic_vector(   0 downto 0);
        signal oVar1S139: std_logic_vector(   0 downto 0);
        signal oVar1S140: std_logic_vector(   0 downto 0);
        signal oVar1S141: std_logic_vector(   0 downto 0);
        signal oVar1S142: std_logic_vector(   0 downto 0);
        signal oVar1S143: std_logic_vector(   0 downto 0);
        signal oVar1S144: std_logic_vector(   0 downto 0);
        signal oVar1S145: std_logic_vector(   0 downto 0);
        signal oVar1S146: std_logic_vector(   0 downto 0);
        signal oVar1S147: std_logic_vector(   0 downto 0);
        signal oVar1S149: std_logic_vector(   0 downto 0);
        signal oVar1S150: std_logic_vector(   0 downto 0);
        signal oVar1S151: std_logic_vector(   0 downto 0);
        signal oVar1S152: std_logic_vector(   0 downto 0);
        signal oVar1S153: std_logic_vector(   0 downto 0);
        signal oVar1S154: std_logic_vector(   0 downto 0);
        signal oVar1S155: std_logic_vector(   0 downto 0);
        signal oVar1S156: std_logic_vector(   0 downto 0);
        signal oVar1S157: std_logic_vector(   0 downto 0);
        signal oVar1S158: std_logic_vector(   0 downto 0);
        signal oVar1S159: std_logic_vector(   0 downto 0);
        signal oVar1S160: std_logic_vector(   0 downto 0);
        signal oVar1S161: std_logic_vector(   0 downto 0);
        signal oVar1S163: std_logic_vector(   0 downto 0);
        signal oVar1S164: std_logic_vector(   0 downto 0);
        signal oVar1S165: std_logic_vector(   0 downto 0);
        signal oVar1S166: std_logic_vector(   0 downto 0);
        signal oVar1S167: std_logic_vector(   0 downto 0);
        signal oVar1S169: std_logic_vector(   0 downto 0);
        signal oVar1S170: std_logic_vector(   0 downto 0);
        signal oVar1S171: std_logic_vector(   0 downto 0);
        signal oVar1S172: std_logic_vector(   0 downto 0);
        signal oVar1S173: std_logic_vector(   0 downto 0);
        signal oVar1S175: std_logic_vector(   0 downto 0);
        signal oVar1S176: std_logic_vector(   0 downto 0);
        signal oVar1S177: std_logic_vector(   0 downto 0);
        signal oVar1S178: std_logic_vector(   0 downto 0);
        signal oVar1S179: std_logic_vector(   0 downto 0);
        signal oVar1S180: std_logic_vector(   0 downto 0);
        signal oVar1S181: std_logic_vector(   0 downto 0);
        signal oVar1S182: std_logic_vector(   0 downto 0);
        signal oVar1S183: std_logic_vector(   0 downto 0);
        signal oVar1S184: std_logic_vector(   0 downto 0);
        signal oVar1S185: std_logic_vector(   0 downto 0);
        signal oVar1S186: std_logic_vector(   0 downto 0);
        signal oVar1S187: std_logic_vector(   0 downto 0);
        signal oVar1S188: std_logic_vector(   0 downto 0);
        signal oVar1S189: std_logic_vector(   0 downto 0);
        signal oVar1S190: std_logic_vector(   0 downto 0);
        signal oVar1S191: std_logic_vector(   0 downto 0);
        signal oVar1S192: std_logic_vector(   0 downto 0);
        signal oVar1S193: std_logic_vector(   0 downto 0);
        signal oVar1S194: std_logic_vector(   0 downto 0);
        signal oVar1S195: std_logic_vector(   0 downto 0);
        signal oVar1S196: std_logic_vector(   0 downto 0);
        signal oVar1S197: std_logic_vector(   0 downto 0);
        signal oVar1S198: std_logic_vector(   0 downto 0);
        signal oVar1S199: std_logic_vector(   0 downto 0);
        signal oVar1S200: std_logic_vector(   0 downto 0);
        signal oVar1S201: std_logic_vector(   0 downto 0);
        signal oVar1S202: std_logic_vector(   0 downto 0);
        signal oVar1S203: std_logic_vector(   0 downto 0);
        signal oVar1S204: std_logic_vector(   0 downto 0);
        signal oVar1S205: std_logic_vector(   0 downto 0);
        signal oVar1S206: std_logic_vector(   0 downto 0);
        signal oVar1S207: std_logic_vector(   0 downto 0);
        signal oVar1S208: std_logic_vector(   0 downto 0);
        signal oVar1S209: std_logic_vector(   0 downto 0);
        signal oVar1S210: std_logic_vector(   0 downto 0);
        signal oVar1S211: std_logic_vector(   0 downto 0);
        signal oVar1S212: std_logic_vector(   0 downto 0);
        signal oVar1S213: std_logic_vector(   0 downto 0);
        signal oVar1S214: std_logic_vector(   0 downto 0);
        signal oVar1S215: std_logic_vector(   0 downto 0);
        signal oVar1S216: std_logic_vector(   0 downto 0);
        signal oVar1S217: std_logic_vector(   0 downto 0);
        signal oVar1S218: std_logic_vector(   0 downto 0);
        signal oVar1S219: std_logic_vector(   0 downto 0);
        signal oVar1S220: std_logic_vector(   0 downto 0);
        signal oVar1S221: std_logic_vector(   0 downto 0);
        signal oVar1S222: std_logic_vector(   0 downto 0);
        signal oVar1S223: std_logic_vector(   0 downto 0);
        signal oVar1S224: std_logic_vector(   0 downto 0);
        signal oVar1S225: std_logic_vector(   0 downto 0);
        signal oVar1S226: std_logic_vector(   0 downto 0);
        signal oVar1S227: std_logic_vector(   0 downto 0);
        signal oVar1S228: std_logic_vector(   0 downto 0);
        signal oVar1S229: std_logic_vector(   0 downto 0);
        signal oVar1S230: std_logic_vector(   0 downto 0);
        signal oVar1S231: std_logic_vector(   0 downto 0);
        signal oVar1S232: std_logic_vector(   0 downto 0);
        signal oVar1S233: std_logic_vector(   0 downto 0);
        signal oVar1S235: std_logic_vector(   0 downto 0);
        signal oVar1S236: std_logic_vector(   0 downto 0);
        signal oVar1S237: std_logic_vector(   0 downto 0);
        signal oVar1S238: std_logic_vector(   0 downto 0);
        signal oVar1S239: std_logic_vector(   0 downto 0);
        signal oVar1S240: std_logic_vector(   0 downto 0);
        signal oVar1S241: std_logic_vector(   0 downto 0);
        signal oVar1S242: std_logic_vector(   0 downto 0);
        signal oVar1S243: std_logic_vector(   0 downto 0);
        signal oVar1S244: std_logic_vector(   0 downto 0);
        signal oVar1S245: std_logic_vector(   0 downto 0);
        signal oVar1S246: std_logic_vector(   0 downto 0);
        signal oVar1S247: std_logic_vector(   0 downto 0);
        signal oVar1S248: std_logic_vector(   0 downto 0);
        signal oVar1S249: std_logic_vector(   0 downto 0);
        signal oVar1S250: std_logic_vector(   0 downto 0);
        signal oVar1S251: std_logic_vector(   0 downto 0);
        signal oVar1S252: std_logic_vector(   0 downto 0);
        signal oVar1S253: std_logic_vector(   0 downto 0);
        signal oVar1S254: std_logic_vector(   0 downto 0);
        signal oVar1S255: std_logic_vector(   0 downto 0);
        signal oVar1S256: std_logic_vector(   0 downto 0);
        signal oVar1S257: std_logic_vector(   0 downto 0);
        signal oVar1S258: std_logic_vector(   0 downto 0);
        signal oVar1S259: std_logic_vector(   0 downto 0);
        signal oVar1S260: std_logic_vector(   0 downto 0);
        signal oVar1S261: std_logic_vector(   0 downto 0);
        signal oVar1S262: std_logic_vector(   0 downto 0);
        signal oVar1S263: std_logic_vector(   0 downto 0);
        signal oVar1S264: std_logic_vector(   0 downto 0);
        signal oVar1S265: std_logic_vector(   0 downto 0);
        signal oVar1S266: std_logic_vector(   0 downto 0);
        signal oVar1S267: std_logic_vector(   0 downto 0);
        signal oVar1S268: std_logic_vector(   0 downto 0);
        signal oVar1S269: std_logic_vector(   0 downto 0);
        signal oVar1S270: std_logic_vector(   0 downto 0);
        signal oVar1S271: std_logic_vector(   0 downto 0);
        signal oVar1S272: std_logic_vector(   0 downto 0);
        signal oVar1S273: std_logic_vector(   0 downto 0);
        signal oVar1S274: std_logic_vector(   0 downto 0);
        signal oVar1S275: std_logic_vector(   0 downto 0);
        signal oVar1S276: std_logic_vector(   0 downto 0);
        signal oVar1S277: std_logic_vector(   0 downto 0);
        signal oVar1S278: std_logic_vector(   0 downto 0);
        signal oVar1S279: std_logic_vector(   0 downto 0);
        signal oVar1S280: std_logic_vector(   0 downto 0);
        signal oVar1S281: std_logic_vector(   0 downto 0);
        signal oVar1S282: std_logic_vector(   0 downto 0);
        signal oVar1S283: std_logic_vector(   0 downto 0);
        signal oVar1S284: std_logic_vector(   0 downto 0);
        signal oVar1S285: std_logic_vector(   0 downto 0);
        signal oVar1S286: std_logic_vector(   0 downto 0);
        signal oVar1S287: std_logic_vector(   0 downto 0);
        signal oVar1S288: std_logic_vector(   0 downto 0);
        signal oVar1S289: std_logic_vector(   0 downto 0);
        signal oVar1S290: std_logic_vector(   0 downto 0);
        signal oVar1S291: std_logic_vector(   0 downto 0);
        signal oVar1S292: std_logic_vector(   0 downto 0);
        signal oVar1S293: std_logic_vector(   0 downto 0);
        signal oVar1S294: std_logic_vector(   0 downto 0);
        signal oVar1S295: std_logic_vector(   0 downto 0);
        signal oVar1S296: std_logic_vector(   0 downto 0);
        signal oVar1S297: std_logic_vector(   0 downto 0);
        signal oVar1S298: std_logic_vector(   0 downto 0);
        signal oVar1S299: std_logic_vector(   0 downto 0);
        signal oVar1S300: std_logic_vector(   0 downto 0);
        signal oVar1S301: std_logic_vector(   0 downto 0);
        signal oVar1S302: std_logic_vector(   0 downto 0);
        signal oVar1S303: std_logic_vector(   0 downto 0);
        signal oVar1S304: std_logic_vector(   0 downto 0);
        signal oVar1S305: std_logic_vector(   0 downto 0);
        signal oVar1S306: std_logic_vector(   0 downto 0);
        signal oVar1S307: std_logic_vector(   0 downto 0);
        signal oVar1S308: std_logic_vector(   0 downto 0);
        signal oVar1S309: std_logic_vector(   0 downto 0);
        signal oVar1S310: std_logic_vector(   0 downto 0);
        signal oVar1S311: std_logic_vector(   0 downto 0);
        signal oVar1S312: std_logic_vector(   0 downto 0);
        signal oVar1S313: std_logic_vector(   0 downto 0);
        signal oVar1S314: std_logic_vector(   0 downto 0);
        signal oVar1S315: std_logic_vector(   0 downto 0);
        signal oVar1S316: std_logic_vector(   0 downto 0);
        signal oVar1S317: std_logic_vector(   0 downto 0);
        signal oVar1S318: std_logic_vector(   0 downto 0);
        signal oVar1S319: std_logic_vector(   0 downto 0);
        signal oVar1S320: std_logic_vector(   0 downto 0);
        signal oVar1S321: std_logic_vector(   0 downto 0);
        signal oVar1S322: std_logic_vector(   0 downto 0);
        signal oVar1S323: std_logic_vector(   0 downto 0);
        signal oVar1S324: std_logic_vector(   0 downto 0);
        signal oVar1S325: std_logic_vector(   0 downto 0);
        signal oVar1S326: std_logic_vector(   0 downto 0);
        signal oVar1S327: std_logic_vector(   0 downto 0);
        signal oVar1S328: std_logic_vector(   0 downto 0);
        signal oVar1S329: std_logic_vector(   0 downto 0);
        signal oVar1S330: std_logic_vector(   0 downto 0);
        signal oVar1S331: std_logic_vector(   0 downto 0);
        signal oVar1S332: std_logic_vector(   0 downto 0);
        signal oVar1S333: std_logic_vector(   0 downto 0);
        signal oVar1S334: std_logic_vector(   0 downto 0);
        signal oVar1S335: std_logic_vector(   0 downto 0);
        signal oVar1S336: std_logic_vector(   0 downto 0);
        signal oVar1S337: std_logic_vector(   0 downto 0);
        signal oVar1S338: std_logic_vector(   0 downto 0);
        signal oVar1S339: std_logic_vector(   0 downto 0);
        signal oVar1S340: std_logic_vector(   0 downto 0);
        signal oVar1S341: std_logic_vector(   0 downto 0);
        signal oVar1S342: std_logic_vector(   0 downto 0);
        signal oVar1S343: std_logic_vector(   0 downto 0);
        signal oVar1S344: std_logic_vector(   0 downto 0);
        signal oVar1S345: std_logic_vector(   0 downto 0);
        signal oVar1S346: std_logic_vector(   0 downto 0);
        signal oVar1S347: std_logic_vector(   0 downto 0);
        signal oVar1S348: std_logic_vector(   0 downto 0);
        signal oVar1S349: std_logic_vector(   0 downto 0);
        signal oVar1S350: std_logic_vector(   0 downto 0);
        signal oVar1S351: std_logic_vector(   0 downto 0);
        signal oVar1S352: std_logic_vector(   0 downto 0);
        signal oVar1S353: std_logic_vector(   0 downto 0);
        signal oVar1S354: std_logic_vector(   0 downto 0);
        signal oVar1S355: std_logic_vector(   0 downto 0);
        signal oVar1S356: std_logic_vector(   0 downto 0);
        signal oVar1S357: std_logic_vector(   0 downto 0);
        signal oVar1S358: std_logic_vector(   0 downto 0);
        signal oVar1S359: std_logic_vector(   0 downto 0);
        signal oVar1S360: std_logic_vector(   0 downto 0);
        signal oVar1S361: std_logic_vector(   0 downto 0);
        signal oVar1S362: std_logic_vector(   0 downto 0);
        signal oVar1S363: std_logic_vector(   0 downto 0);
        signal oVar1S364: std_logic_vector(   0 downto 0);
        signal oVar1S365: std_logic_vector(   0 downto 0);
        signal oVar1S366: std_logic_vector(   0 downto 0);
        signal oVar1S367: std_logic_vector(   0 downto 0);
        signal oVar1S368: std_logic_vector(   0 downto 0);
        signal oVar1S369: std_logic_vector(   0 downto 0);
        signal oVar1S370: std_logic_vector(   0 downto 0);
        signal oVar1S371: std_logic_vector(   0 downto 0);
        signal oVar1S372: std_logic_vector(   0 downto 0);
        signal oVar1S373: std_logic_vector(   0 downto 0);
        signal oVar1S374: std_logic_vector(   0 downto 0);
        signal oVar1S375: std_logic_vector(   0 downto 0);
        signal oVar1S376: std_logic_vector(   0 downto 0);
        signal oVar1S377: std_logic_vector(   0 downto 0);
        signal oVar1S378: std_logic_vector(   0 downto 0);
        signal oVar1S379: std_logic_vector(   0 downto 0);
        signal oVar1S380: std_logic_vector(   0 downto 0);
        signal oVar1S381: std_logic_vector(   0 downto 0);
        signal oVar1S383: std_logic_vector(   0 downto 0);
        signal oVar1S384: std_logic_vector(   0 downto 0);
        signal oVar1S385: std_logic_vector(   0 downto 0);
        signal oVar1S386: std_logic_vector(   0 downto 0);
        signal oVar1S387: std_logic_vector(   0 downto 0);
        signal oVar1S388: std_logic_vector(   0 downto 0);
        signal oVar1S389: std_logic_vector(   0 downto 0);
        signal oVar1S390: std_logic_vector(   0 downto 0);
        signal oVar1S391: std_logic_vector(   0 downto 0);
        signal oVar1S392: std_logic_vector(   0 downto 0);
        signal oVar1S393: std_logic_vector(   0 downto 0);
        signal oVar1S394: std_logic_vector(   0 downto 0);
        signal oVar1S395: std_logic_vector(   0 downto 0);
        signal oVar1S397: std_logic_vector(   0 downto 0);
        signal oVar1S398: std_logic_vector(   0 downto 0);
        signal oVar1S399: std_logic_vector(   0 downto 0);
        signal oVar1S400: std_logic_vector(   0 downto 0);
        signal oVar1S401: std_logic_vector(   0 downto 0);
        signal oVar1S402: std_logic_vector(   0 downto 0);
        signal oVar1S403: std_logic_vector(   0 downto 0);
        signal oVar1S404: std_logic_vector(   0 downto 0);
        signal oVar1S405: std_logic_vector(   0 downto 0);
        signal oVar1S406: std_logic_vector(   0 downto 0);
        signal oVar1S407: std_logic_vector(   0 downto 0);
        signal oVar1S408: std_logic_vector(   0 downto 0);
        signal oVar1S409: std_logic_vector(   0 downto 0);
        signal oVar1S410: std_logic_vector(   0 downto 0);
        signal oVar1S411: std_logic_vector(   0 downto 0);
        signal oVar1S412: std_logic_vector(   0 downto 0);
        signal oVar1S413: std_logic_vector(   0 downto 0);
        signal oVar1S414: std_logic_vector(   0 downto 0);
        signal oVar1S415: std_logic_vector(   0 downto 0);
        signal oVar1S416: std_logic_vector(   0 downto 0);
        signal oVar1S417: std_logic_vector(   0 downto 0);
        signal oVar1S418: std_logic_vector(   0 downto 0);
        signal oVar1S419: std_logic_vector(   0 downto 0);
        signal oVar1S420: std_logic_vector(   0 downto 0);
        signal oVar1S421: std_logic_vector(   0 downto 0);
        signal oVar1S422: std_logic_vector(   0 downto 0);
        signal oVar1S423: std_logic_vector(   0 downto 0);
        signal oVar1S424: std_logic_vector(   0 downto 0);
        signal oVar1S425: std_logic_vector(   0 downto 0);
        signal oVar1S427: std_logic_vector(   0 downto 0);
        signal oVar1S428: std_logic_vector(   0 downto 0);
        signal oVar1S429: std_logic_vector(   0 downto 0);
        signal oVar1S430: std_logic_vector(   0 downto 0);
        signal oVar1S431: std_logic_vector(   0 downto 0);
        signal oVar1S433: std_logic_vector(   0 downto 0);
        signal oVar1S434: std_logic_vector(   0 downto 0);
        signal oVar1S435: std_logic_vector(   0 downto 0);
        signal oVar1S436: std_logic_vector(   0 downto 0);
        signal oVar1S437: std_logic_vector(   0 downto 0);
        signal oVar1S438: std_logic_vector(   0 downto 0);
        signal oVar1S439: std_logic_vector(   0 downto 0);
        signal oVar1S440: std_logic_vector(   0 downto 0);
        signal oVar1S441: std_logic_vector(   0 downto 0);
        signal oVar1S442: std_logic_vector(   0 downto 0);
        signal oVar1S443: std_logic_vector(   0 downto 0);
        signal oVar1S444: std_logic_vector(   0 downto 0);
        signal oVar1S445: std_logic_vector(   0 downto 0);
        signal oVar1S446: std_logic_vector(   0 downto 0);
        signal oVar1S447: std_logic_vector(   0 downto 0);
        signal oVar1S448: std_logic_vector(   0 downto 0);
        signal oVar1S449: std_logic_vector(   0 downto 0);
        signal oVar1S450: std_logic_vector(   0 downto 0);
        signal oVar1S451: std_logic_vector(   0 downto 0);
        signal oVar1S452: std_logic_vector(   0 downto 0);
        signal oVar1S453: std_logic_vector(   0 downto 0);
        signal oVar1S454: std_logic_vector(   0 downto 0);
        signal oVar1S455: std_logic_vector(   0 downto 0);
        signal oVar1S456: std_logic_vector(   0 downto 0);
        signal oVar1S457: std_logic_vector(   0 downto 0);
        signal oVar1S458: std_logic_vector(   0 downto 0);
        signal oVar1S459: std_logic_vector(   0 downto 0);
        signal oVar1S461: std_logic_vector(   0 downto 0);
        signal oVar1S462: std_logic_vector(   0 downto 0);
        signal oVar1S463: std_logic_vector(   0 downto 0);
        signal oVar1S464: std_logic_vector(   0 downto 0);
        signal oVar1S465: std_logic_vector(   0 downto 0);
        signal oVar1S466: std_logic_vector(   0 downto 0);
        signal oVar1S467: std_logic_vector(   0 downto 0);
        signal oVar1S468: std_logic_vector(   0 downto 0);
        signal oVar1S469: std_logic_vector(   0 downto 0);
        signal oVar1S470: std_logic_vector(   0 downto 0);
        signal oVar1S471: std_logic_vector(   0 downto 0);
        signal oVar1S472: std_logic_vector(   0 downto 0);
        signal oVar1S473: std_logic_vector(   0 downto 0);
        signal oVar1S474: std_logic_vector(   0 downto 0);
        signal oVar1S475: std_logic_vector(   0 downto 0);
        signal oVar1S476: std_logic_vector(   0 downto 0);
        signal oVar1S477: std_logic_vector(   0 downto 0);
        signal oVar1S478: std_logic_vector(   0 downto 0);
        signal oVar1S479: std_logic_vector(   0 downto 0);
        signal oVar1S480: std_logic_vector(   0 downto 0);
        signal oVar1S481: std_logic_vector(   0 downto 0);
        signal oVar1S482: std_logic_vector(   0 downto 0);
        signal oVar1S483: std_logic_vector(   0 downto 0);
        signal oVar1S484: std_logic_vector(   0 downto 0);
        signal oVar1S486: std_logic_vector(   0 downto 0);
        signal oVar1S487: std_logic_vector(   0 downto 0);
        signal oVar1S488: std_logic_vector(   0 downto 0);
        signal oVar1S489: std_logic_vector(   0 downto 0);
        signal oVar1S490: std_logic_vector(   0 downto 0);
        signal oVar1S491: std_logic_vector(   0 downto 0);
        signal oVar1S492: std_logic_vector(   0 downto 0);
        signal oVar1S493: std_logic_vector(   0 downto 0);
        signal oVar1S494: std_logic_vector(   0 downto 0);
        signal oVar1S495: std_logic_vector(   0 downto 0);
        signal oVar1S496: std_logic_vector(   0 downto 0);
        signal oVar1S497: std_logic_vector(   0 downto 0);
        signal oVar1S498: std_logic_vector(   0 downto 0);
        signal oVar1S499: std_logic_vector(   0 downto 0);
        signal oVar1S500: std_logic_vector(   0 downto 0);
        signal oVar1S501: std_logic_vector(   0 downto 0);
        signal oVar1S502: std_logic_vector(   0 downto 0);
        signal oVar1S503: std_logic_vector(   0 downto 0);
        signal oVar1S504: std_logic_vector(   0 downto 0);
        signal oVar1S505: std_logic_vector(   0 downto 0);
        signal oVar1S506: std_logic_vector(   0 downto 0);
        signal oVar1S507: std_logic_vector(   0 downto 0);
        signal oVar1S508: std_logic_vector(   0 downto 0);
        signal oVar1S509: std_logic_vector(   0 downto 0);
        signal oVar1S511: std_logic_vector(   0 downto 0);
        signal oVar1S512: std_logic_vector(   0 downto 0);
        signal oVar1S513: std_logic_vector(   0 downto 0);
        signal oVar1S514: std_logic_vector(   0 downto 0);
        signal oVar1S516: std_logic_vector(   0 downto 0);
        signal oVar1S517: std_logic_vector(   0 downto 0);
        signal oVar1S518: std_logic_vector(   0 downto 0);
        signal oVar1S519: std_logic_vector(   0 downto 0);
        signal oVar1S520: std_logic_vector(   0 downto 0);
        signal oVar1S521: std_logic_vector(   0 downto 0);
        signal oVar1S522: std_logic_vector(   0 downto 0);
        signal oVar1S523: std_logic_vector(   0 downto 0);
        signal oVar1S524: std_logic_vector(   0 downto 0);
        signal oVar1S525: std_logic_vector(   0 downto 0);
        signal oVar1S526: std_logic_vector(   0 downto 0);
        signal oVar1S527: std_logic_vector(   0 downto 0);
        signal oVar1S528: std_logic_vector(   0 downto 0);
        signal oVar1S529: std_logic_vector(   0 downto 0);
        signal oVar1S530: std_logic_vector(   0 downto 0);
        signal oVar1S531: std_logic_vector(   0 downto 0);
        signal oVar1S532: std_logic_vector(   0 downto 0);
        signal oVar1S533: std_logic_vector(   0 downto 0);
        signal oVar1S534: std_logic_vector(   0 downto 0);
        signal oVar1S536: std_logic_vector(   0 downto 0);
        signal oVar1S537: std_logic_vector(   0 downto 0);
        signal oVar1S538: std_logic_vector(   0 downto 0);
        signal oVar1S539: std_logic_vector(   0 downto 0);
        signal oVar1S540: std_logic_vector(   0 downto 0);
        signal oVar1S541: std_logic_vector(   0 downto 0);
        signal oVar1S542: std_logic_vector(   0 downto 0);
        signal oVar1S543: std_logic_vector(   0 downto 0);
        signal oVar1S544: std_logic_vector(   0 downto 0);
        signal oVar1S545: std_logic_vector(   0 downto 0);
        signal oVar1S546: std_logic_vector(   0 downto 0);
        signal oVar1S547: std_logic_vector(   0 downto 0);
        signal oVar1S548: std_logic_vector(   0 downto 0);
        signal oVar1S549: std_logic_vector(   0 downto 0);
        signal oVar1S550: std_logic_vector(   0 downto 0);
        signal oVar1S551: std_logic_vector(   0 downto 0);
        signal oVar1S552: std_logic_vector(   0 downto 0);
        signal oVar1S553: std_logic_vector(   0 downto 0);
        signal oVar1S554: std_logic_vector(   0 downto 0);
        signal oVar1S555: std_logic_vector(   0 downto 0);
        signal oVar1S556: std_logic_vector(   0 downto 0);
        signal oVar1S557: std_logic_vector(   0 downto 0);
        signal oVar1S558: std_logic_vector(   0 downto 0);
        signal oVar1S559: std_logic_vector(   0 downto 0);
        signal oVar1S560: std_logic_vector(   0 downto 0);
        signal oVar1S561: std_logic_vector(   0 downto 0);
        signal oVar1S562: std_logic_vector(   0 downto 0);
        signal oVar1S563: std_logic_vector(   0 downto 0);
        signal oVar1S565: std_logic_vector(   0 downto 0);
        signal oVar1S566: std_logic_vector(   0 downto 0);
        signal oVar1S567: std_logic_vector(   0 downto 0);
        signal oVar1S568: std_logic_vector(   0 downto 0);
        signal oVar1S569: std_logic_vector(   0 downto 0);
        signal oVar1S571: std_logic_vector(   0 downto 0);
        signal oVar1S572: std_logic_vector(   0 downto 0);
        signal oVar1S573: std_logic_vector(   0 downto 0);
        signal oVar1S574: std_logic_vector(   0 downto 0);
        signal oVar1S575: std_logic_vector(   0 downto 0);
        signal oVar1S576: std_logic_vector(   0 downto 0);
        signal oVar1S577: std_logic_vector(   0 downto 0);
        signal oVar1S578: std_logic_vector(   0 downto 0);
        signal oVar1S579: std_logic_vector(   0 downto 0);
        signal oVar1S580: std_logic_vector(   0 downto 0);
        signal oVar1S581: std_logic_vector(   0 downto 0);
        signal oVar1S582: std_logic_vector(   0 downto 0);
        signal oVar1S583: std_logic_vector(   0 downto 0);
        signal oVar1S584: std_logic_vector(   0 downto 0);
        signal oVar1S585: std_logic_vector(   0 downto 0);
        signal oVar1S586: std_logic_vector(   0 downto 0);
        signal oVar1S587: std_logic_vector(   0 downto 0);
        signal oVar1S588: std_logic_vector(   0 downto 0);
        signal oVar1S589: std_logic_vector(   0 downto 0);
        signal oVar1S591: std_logic_vector(   0 downto 0);
        signal oVar1S592: std_logic_vector(   0 downto 0);
        signal oVar1S593: std_logic_vector(   0 downto 0);
        signal oVar1S595: std_logic_vector(   0 downto 0);
        signal oVar1S596: std_logic_vector(   0 downto 0);
        signal oVar1S597: std_logic_vector(   0 downto 0);
        signal oVar1S598: std_logic_vector(   0 downto 0);
        signal oVar1S599: std_logic_vector(   0 downto 0);
        signal oVar1S600: std_logic_vector(   0 downto 0);
        signal oVar1S601: std_logic_vector(   0 downto 0);
        signal oVar1S603: std_logic_vector(   0 downto 0);
        signal oVar1S604: std_logic_vector(   0 downto 0);
        signal oVar1S605: std_logic_vector(   0 downto 0);
        signal oVar1S606: std_logic_vector(   0 downto 0);
        signal oVar1S607: std_logic_vector(   0 downto 0);
        signal oVar1S608: std_logic_vector(   0 downto 0);
        signal oVar1S609: std_logic_vector(   0 downto 0);
        signal oVar1S610: std_logic_vector(   0 downto 0);
        signal oVar1S611: std_logic_vector(   0 downto 0);
        signal oVar1S612: std_logic_vector(   0 downto 0);
        signal oVar1S613: std_logic_vector(   0 downto 0);
        signal oVar1S615: std_logic_vector(   0 downto 0);
        signal oVar1S616: std_logic_vector(   0 downto 0);
        signal oVar1S617: std_logic_vector(   0 downto 0);
        signal oVar1S618: std_logic_vector(   0 downto 0);
        signal oVar1S619: std_logic_vector(   0 downto 0);
        signal oVar1S620: std_logic_vector(   0 downto 0);
        signal oVar1S621: std_logic_vector(   0 downto 0);
        signal oVar1S623: std_logic_vector(   0 downto 0);
        signal oVar1S624: std_logic_vector(   0 downto 0);
        signal oVar1S625: std_logic_vector(   0 downto 0);
        signal oVar1S627: std_logic_vector(   0 downto 0);
        signal oVar1S628: std_logic_vector(   0 downto 0);
        signal oVar1S629: std_logic_vector(   0 downto 0);
        signal oVar1S630: std_logic_vector(   0 downto 0);
        signal oVar1S631: std_logic_vector(   0 downto 0);
        signal oVar1S632: std_logic_vector(   0 downto 0);
        signal oVar1S633: std_logic_vector(   0 downto 0);
        signal oVar1S634: std_logic_vector(   0 downto 0);
        signal oVar1S635: std_logic_vector(   0 downto 0);
        signal oVar1S636: std_logic_vector(   0 downto 0);
        signal oVar1S637: std_logic_vector(   0 downto 0);
        signal oVar1S638: std_logic_vector(   0 downto 0);
        signal oVar1S639: std_logic_vector(   0 downto 0);
        signal oVar1S640: std_logic_vector(   0 downto 0);
        signal oVar1S641: std_logic_vector(   0 downto 0);
        signal oVar1S642: std_logic_vector(   0 downto 0);
        signal oVar1S643: std_logic_vector(   0 downto 0);
        signal oVar1S644: std_logic_vector(   0 downto 0);
        signal oVar1S645: std_logic_vector(   0 downto 0);
        signal oVar1S646: std_logic_vector(   0 downto 0);
        signal oVar1S647: std_logic_vector(   0 downto 0);
        signal oVar1S649: std_logic_vector(   0 downto 0);
        signal oVar1S650: std_logic_vector(   0 downto 0);
        signal oVar1S651: std_logic_vector(   0 downto 0);
        signal oVar1S652: std_logic_vector(   0 downto 0);
        signal oVar1S653: std_logic_vector(   0 downto 0);
        signal oVar1S654: std_logic_vector(   0 downto 0);
        signal oVar1S655: std_logic_vector(   0 downto 0);
        signal oVar1S656: std_logic_vector(   0 downto 0);
        signal oVar1S657: std_logic_vector(   0 downto 0);
        signal oVar1S658: std_logic_vector(   0 downto 0);
        signal oVar1S659: std_logic_vector(   0 downto 0);
        signal oVar1S660: std_logic_vector(   0 downto 0);
        signal oVar1S661: std_logic_vector(   0 downto 0);
        signal oVar1S662: std_logic_vector(   0 downto 0);
        signal oVar1S663: std_logic_vector(   0 downto 0);
        signal oVar1S664: std_logic_vector(   0 downto 0);
        signal oVar1S665: std_logic_vector(   0 downto 0);
        signal oVar1S666: std_logic_vector(   0 downto 0);
        signal oVar1S668: std_logic_vector(   0 downto 0);
        signal oVar1S669: std_logic_vector(   0 downto 0);
        signal oVar1S670: std_logic_vector(   0 downto 0);
        signal oVar1S671: std_logic_vector(   0 downto 0);
        signal oVar1S672: std_logic_vector(   0 downto 0);
        signal oVar1S673: std_logic_vector(   0 downto 0);
        signal oVar1S675: std_logic_vector(   0 downto 0);
        signal oVar1S676: std_logic_vector(   0 downto 0);
        signal oVar1S677: std_logic_vector(   0 downto 0);
        signal oVar1S678: std_logic_vector(   0 downto 0);
        signal oVar1S679: std_logic_vector(   0 downto 0);
        signal oVar1S680: std_logic_vector(   0 downto 0);
        signal oVar1S681: std_logic_vector(   0 downto 0);
        signal oVar1S682: std_logic_vector(   0 downto 0);
        signal oVar1S683: std_logic_vector(   0 downto 0);
        signal oVar1S684: std_logic_vector(   0 downto 0);
        signal oVar1S685: std_logic_vector(   0 downto 0);
        signal oVar1S686: std_logic_vector(   0 downto 0);
        signal oVar1S687: std_logic_vector(   0 downto 0);
        signal oVar1S688: std_logic_vector(   0 downto 0);
        signal oVar1S689: std_logic_vector(   0 downto 0);
        signal oVar1S690: std_logic_vector(   0 downto 0);
        signal oVar1S691: std_logic_vector(   0 downto 0);
        signal oVar1S692: std_logic_vector(   0 downto 0);
        signal oVar1S693: std_logic_vector(   0 downto 0);
        signal oVar1S694: std_logic_vector(   0 downto 0);
        signal oVar1S695: std_logic_vector(   0 downto 0);
        signal oVar2S0: std_logic_vector(   0 downto 0);
        signal oVar2S1: std_logic_vector(   0 downto 0);
        signal oVar2S2: std_logic_vector(   0 downto 0);
        signal oVar2S3: std_logic_vector(   0 downto 0);
        signal oVar2S4: std_logic_vector(   0 downto 0);
        signal oVar2S5: std_logic_vector(   0 downto 0);
        signal oVar2S6: std_logic_vector(   0 downto 0);
        signal oVar2S7: std_logic_vector(   0 downto 0);
        signal oVar2S8: std_logic_vector(   0 downto 0);
        signal oVar2S9: std_logic_vector(   0 downto 0);
        signal oVar2S10: std_logic_vector(   0 downto 0);
        signal oVar2S11: std_logic_vector(   0 downto 0);
        signal oVar2S12: std_logic_vector(   0 downto 0);
        signal oVar2S14: std_logic_vector(   0 downto 0);
        signal oVar2S15: std_logic_vector(   0 downto 0);
        signal oVar2S16: std_logic_vector(   0 downto 0);
        signal oVar2S17: std_logic_vector(   0 downto 0);
        signal oVar2S18: std_logic_vector(   0 downto 0);
        signal oVar2S19: std_logic_vector(   0 downto 0);
        signal oVar2S20: std_logic_vector(   0 downto 0);
        signal oVar2S21: std_logic_vector(   0 downto 0);
        signal oVar2S22: std_logic_vector(   0 downto 0);
        signal oVar2S23: std_logic_vector(   0 downto 0);
        signal oVar2S24: std_logic_vector(   0 downto 0);
        signal oVar2S25: std_logic_vector(   0 downto 0);
        signal oVar2S26: std_logic_vector(   0 downto 0);
        signal oVar2S27: std_logic_vector(   0 downto 0);
        signal oVar2S28: std_logic_vector(   0 downto 0);
        signal oVar2S29: std_logic_vector(   0 downto 0);
        signal oVar2S30: std_logic_vector(   0 downto 0);
        signal oVar2S31: std_logic_vector(   0 downto 0);
        signal oVar2S32: std_logic_vector(   0 downto 0);
        signal oVar2S33: std_logic_vector(   0 downto 0);
        signal oVar2S34: std_logic_vector(   0 downto 0);
        signal oVar2S36: std_logic_vector(   0 downto 0);
        signal oVar2S37: std_logic_vector(   0 downto 0);
        signal oVar2S38: std_logic_vector(   0 downto 0);
        signal oVar2S39: std_logic_vector(   0 downto 0);
        signal oVar2S41: std_logic_vector(   0 downto 0);
        signal oVar2S42: std_logic_vector(   0 downto 0);
        signal oVar2S44: std_logic_vector(   0 downto 0);
        signal oVar2S46: std_logic_vector(   0 downto 0);
        signal oVar2S47: std_logic_vector(   0 downto 0);
        signal oVar2S48: std_logic_vector(   0 downto 0);
        signal oVar2S50: std_logic_vector(   0 downto 0);
        signal oVar2S51: std_logic_vector(   0 downto 0);
        signal oVar2S53: std_logic_vector(   0 downto 0);
        signal oVar2S54: std_logic_vector(   0 downto 0);
        signal oVar2S55: std_logic_vector(   0 downto 0);
        signal oVar2S56: std_logic_vector(   0 downto 0);
        signal oVar2S58: std_logic_vector(   0 downto 0);
        signal oVar2S59: std_logic_vector(   0 downto 0);
        signal oVar2S60: std_logic_vector(   0 downto 0);
        signal oVar2S61: std_logic_vector(   0 downto 0);
        signal oVar2S62: std_logic_vector(   0 downto 0);
        signal oVar2S63: std_logic_vector(   0 downto 0);
        signal oVar2S64: std_logic_vector(   0 downto 0);
        signal oVar2S65: std_logic_vector(   0 downto 0);
        signal oVar2S66: std_logic_vector(   0 downto 0);
        signal oVar2S67: std_logic_vector(   0 downto 0);
        signal oVar2S68: std_logic_vector(   0 downto 0);
        signal oVar2S69: std_logic_vector(   0 downto 0);
        signal oVar2S70: std_logic_vector(   0 downto 0);
        signal oVar2S71: std_logic_vector(   0 downto 0);
        signal oVar2S72: std_logic_vector(   0 downto 0);
        signal oVar2S73: std_logic_vector(   0 downto 0);
        signal oVar2S74: std_logic_vector(   0 downto 0);
        signal oVar2S75: std_logic_vector(   0 downto 0);
        signal oVar2S76: std_logic_vector(   0 downto 0);
        signal oVar2S77: std_logic_vector(   0 downto 0);
        signal oVar2S78: std_logic_vector(   0 downto 0);
        signal oVar2S79: std_logic_vector(   0 downto 0);
        signal oVar2S80: std_logic_vector(   0 downto 0);
        signal oVar2S81: std_logic_vector(   0 downto 0);
        signal oVar2S82: std_logic_vector(   0 downto 0);
        signal oVar2S83: std_logic_vector(   0 downto 0);
        signal oVar2S84: std_logic_vector(   0 downto 0);
        signal oVar2S85: std_logic_vector(   0 downto 0);
        signal oVar2S86: std_logic_vector(   0 downto 0);
        signal oVar2S87: std_logic_vector(   0 downto 0);
        signal oVar2S88: std_logic_vector(   0 downto 0);
        signal oVar2S89: std_logic_vector(   0 downto 0);
        signal oVar2S90: std_logic_vector(   0 downto 0);
        signal oVar2S91: std_logic_vector(   0 downto 0);
        signal oVar2S92: std_logic_vector(   0 downto 0);
        signal oVar2S93: std_logic_vector(   0 downto 0);
        signal oVar2S94: std_logic_vector(   0 downto 0);
        signal oVar2S95: std_logic_vector(   0 downto 0);
        signal oVar2S96: std_logic_vector(   0 downto 0);
        signal oVar2S97: std_logic_vector(   0 downto 0);
        signal oVar2S98: std_logic_vector(   0 downto 0);
        signal oVar2S99: std_logic_vector(   0 downto 0);
        signal oVar2S100: std_logic_vector(   0 downto 0);
        signal oVar2S101: std_logic_vector(   0 downto 0);
        signal oVar2S102: std_logic_vector(   0 downto 0);
        signal oVar2S103: std_logic_vector(   0 downto 0);
        signal oVar2S104: std_logic_vector(   0 downto 0);
        signal oVar2S105: std_logic_vector(   0 downto 0);
        signal oVar2S106: std_logic_vector(   0 downto 0);
        signal oVar2S107: std_logic_vector(   0 downto 0);
        signal oVar2S108: std_logic_vector(   0 downto 0);
        signal oVar2S109: std_logic_vector(   0 downto 0);
        signal oVar2S110: std_logic_vector(   0 downto 0);
        signal oVar2S111: std_logic_vector(   0 downto 0);
        signal oVar2S112: std_logic_vector(   0 downto 0);
        signal oVar2S113: std_logic_vector(   0 downto 0);
        signal oVar2S114: std_logic_vector(   0 downto 0);
        signal oVar2S115: std_logic_vector(   0 downto 0);
        signal oVar2S116: std_logic_vector(   0 downto 0);
        signal oVar2S117: std_logic_vector(   0 downto 0);
        signal oVar2S118: std_logic_vector(   0 downto 0);
        signal oVar2S119: std_logic_vector(   0 downto 0);
        signal oVar2S120: std_logic_vector(   0 downto 0);
        signal oVar2S121: std_logic_vector(   0 downto 0);
        signal oVar2S122: std_logic_vector(   0 downto 0);
        signal oVar2S123: std_logic_vector(   0 downto 0);
        signal oVar2S124: std_logic_vector(   0 downto 0);
        signal oVar2S126: std_logic_vector(   0 downto 0);
        signal oVar2S127: std_logic_vector(   0 downto 0);
        signal oVar2S128: std_logic_vector(   0 downto 0);
        signal oVar2S129: std_logic_vector(   0 downto 0);
        signal oVar2S130: std_logic_vector(   0 downto 0);
        signal oVar2S131: std_logic_vector(   0 downto 0);
        signal oVar2S132: std_logic_vector(   0 downto 0);
        signal oVar2S134: std_logic_vector(   0 downto 0);
        signal oVar2S136: std_logic_vector(   0 downto 0);
        signal oVar2S137: std_logic_vector(   0 downto 0);
        signal oVar2S138: std_logic_vector(   0 downto 0);
        signal oVar2S140: std_logic_vector(   0 downto 0);
        signal oVar2S142: std_logic_vector(   0 downto 0);
        signal oVar2S144: std_logic_vector(   0 downto 0);
        signal oVar2S146: std_logic_vector(   0 downto 0);
        signal oVar2S148: std_logic_vector(   0 downto 0);
        signal oVar2S149: std_logic_vector(   0 downto 0);
        signal oVar2S150: std_logic_vector(   0 downto 0);
        signal oVar2S151: std_logic_vector(   0 downto 0);
        signal oVar2S152: std_logic_vector(   0 downto 0);
        signal oVar2S153: std_logic_vector(   0 downto 0);
        signal oVar2S154: std_logic_vector(   0 downto 0);
        signal oVar2S155: std_logic_vector(   0 downto 0);
        signal oVar2S156: std_logic_vector(   0 downto 0);
        signal oVar2S157: std_logic_vector(   0 downto 0);
        signal oVar2S159: std_logic_vector(   0 downto 0);
        signal oVar2S160: std_logic_vector(   0 downto 0);
        signal oVar2S161: std_logic_vector(   0 downto 0);
        signal oVar2S162: std_logic_vector(   0 downto 0);
        signal oVar2S164: std_logic_vector(   0 downto 0);
        signal oVar2S165: std_logic_vector(   0 downto 0);
        signal oVar2S166: std_logic_vector(   0 downto 0);
        signal oVar2S167: std_logic_vector(   0 downto 0);
        signal oVar2S168: std_logic_vector(   0 downto 0);
        signal oVar2S169: std_logic_vector(   0 downto 0);
        signal oVar2S170: std_logic_vector(   0 downto 0);
        signal oVar2S171: std_logic_vector(   0 downto 0);
        signal oVar2S172: std_logic_vector(   0 downto 0);
        signal oVar2S173: std_logic_vector(   0 downto 0);
        signal oVar2S174: std_logic_vector(   0 downto 0);
        signal oVar2S175: std_logic_vector(   0 downto 0);
        signal oVar2S176: std_logic_vector(   0 downto 0);
        signal oVar2S177: std_logic_vector(   0 downto 0);
        signal oVar2S178: std_logic_vector(   0 downto 0);
        signal oVar2S179: std_logic_vector(   0 downto 0);
        signal oVar2S180: std_logic_vector(   0 downto 0);
        signal oVar2S181: std_logic_vector(   0 downto 0);
        signal oVar2S182: std_logic_vector(   0 downto 0);
        signal oVar2S184: std_logic_vector(   0 downto 0);
        signal oVar2S185: std_logic_vector(   0 downto 0);
        signal oVar2S186: std_logic_vector(   0 downto 0);
        signal oVar2S187: std_logic_vector(   0 downto 0);
        signal oVar2S188: std_logic_vector(   0 downto 0);
        signal oVar2S189: std_logic_vector(   0 downto 0);
        signal oVar2S190: std_logic_vector(   0 downto 0);
        signal oVar2S191: std_logic_vector(   0 downto 0);
        signal oVar2S192: std_logic_vector(   0 downto 0);
        signal oVar2S193: std_logic_vector(   0 downto 0);
        signal oVar2S194: std_logic_vector(   0 downto 0);
        signal oVar2S196: std_logic_vector(   0 downto 0);
        signal oVar2S197: std_logic_vector(   0 downto 0);
        signal oVar2S198: std_logic_vector(   0 downto 0);
        signal oVar2S199: std_logic_vector(   0 downto 0);
        signal oVar2S200: std_logic_vector(   0 downto 0);
        signal oVar2S201: std_logic_vector(   0 downto 0);
        signal oVar2S202: std_logic_vector(   0 downto 0);
        signal oVar2S204: std_logic_vector(   0 downto 0);
        signal oVar2S205: std_logic_vector(   0 downto 0);
        signal oVar2S206: std_logic_vector(   0 downto 0);
        signal oVar2S208: std_logic_vector(   0 downto 0);
        signal oVar2S209: std_logic_vector(   0 downto 0);
        signal oVar2S210: std_logic_vector(   0 downto 0);
        signal oVar2S212: std_logic_vector(   0 downto 0);
        signal oVar2S214: std_logic_vector(   0 downto 0);
        signal oVar2S216: std_logic_vector(   0 downto 0);
        signal oVar2S217: std_logic_vector(   0 downto 0);
        signal oVar2S218: std_logic_vector(   0 downto 0);
        signal oVar2S219: std_logic_vector(   0 downto 0);
        signal oVar2S221: std_logic_vector(   0 downto 0);
        signal oVar2S223: std_logic_vector(   0 downto 0);
        signal oVar2S225: std_logic_vector(   0 downto 0);
        signal oVar2S227: std_logic_vector(   0 downto 0);
        signal oVar2S228: std_logic_vector(   0 downto 0);
        signal oVar2S229: std_logic_vector(   0 downto 0);
        signal oVar2S231: std_logic_vector(   0 downto 0);
        signal oVar2S232: std_logic_vector(   0 downto 0);
        signal oVar2S233: std_logic_vector(   0 downto 0);
        signal oVar2S235: std_logic_vector(   0 downto 0);
        signal oVar2S237: std_logic_vector(   0 downto 0);
        signal oVar2S238: std_logic_vector(   0 downto 0);
        signal oVar2S239: std_logic_vector(   0 downto 0);
        signal oVar2S241: std_logic_vector(   0 downto 0);
        signal oVar2S243: std_logic_vector(   0 downto 0);
        signal oVar2S245: std_logic_vector(   0 downto 0);
        signal oVar2S246: std_logic_vector(   0 downto 0);
        signal oVar2S247: std_logic_vector(   0 downto 0);
        signal oVar2S248: std_logic_vector(   0 downto 0);
        signal oVar2S249: std_logic_vector(   0 downto 0);
        signal oVar2S250: std_logic_vector(   0 downto 0);
        signal oVar2S251: std_logic_vector(   0 downto 0);
        signal oVar2S252: std_logic_vector(   0 downto 0);
        signal oVar3S0: std_logic_vector(   0 downto 0);
        signal oVar3S1: std_logic_vector(   0 downto 0);
        signal oVar3S2: std_logic_vector(   0 downto 0);
        signal oVar3S3: std_logic_vector(   0 downto 0);
        signal oVar3S4: std_logic_vector(   0 downto 0);
        signal oVar3S5: std_logic_vector(   0 downto 0);
        signal oVar3S6: std_logic_vector(   0 downto 0);
        signal oVar3S7: std_logic_vector(   0 downto 0);
        signal oVar3S8: std_logic_vector(   0 downto 0);
        signal oVar3S9: std_logic_vector(   0 downto 0);
        signal oVar3S10: std_logic_vector(   0 downto 0);
        signal oVar3S11: std_logic_vector(   0 downto 0);
        signal oVar3S12: std_logic_vector(   0 downto 0);
        signal oVar3S13: std_logic_vector(   0 downto 0);
        signal oVar3S14: std_logic_vector(   0 downto 0);
        signal oVar3S15: std_logic_vector(   0 downto 0);
        signal oVar3S16: std_logic_vector(   0 downto 0);
        signal oVar3S17: std_logic_vector(   0 downto 0);
        signal oVar3S18: std_logic_vector(   0 downto 0);
        signal oVar3S19: std_logic_vector(   0 downto 0);
        signal oVar3S20: std_logic_vector(   0 downto 0);
        signal oVar3S21: std_logic_vector(   0 downto 0);
        signal oVar3S22: std_logic_vector(   0 downto 0);
        signal oVar3S23: std_logic_vector(   0 downto 0);
        signal oVar3S24: std_logic_vector(   0 downto 0);
        signal oVar3S25: std_logic_vector(   0 downto 0);
        signal oVar3S26: std_logic_vector(   0 downto 0);
        signal oVar3S27: std_logic_vector(   0 downto 0);
        signal oVar3S28: std_logic_vector(   0 downto 0);
        signal oVar3S29: std_logic_vector(   0 downto 0);
        signal oVar3S30: std_logic_vector(   0 downto 0);
        signal oVar3S31: std_logic_vector(   0 downto 0);
        signal oVar3S32: std_logic_vector(   0 downto 0);
        signal oVar3S33: std_logic_vector(   0 downto 0);
        signal oVar3S34: std_logic_vector(   0 downto 0);
        signal oVar3S35: std_logic_vector(   0 downto 0);
        signal oVar3S36: std_logic_vector(   0 downto 0);
        signal oVar3S37: std_logic_vector(   0 downto 0);
        signal oVar3S38: std_logic_vector(   0 downto 0);
        signal oVar3S39: std_logic_vector(   0 downto 0);
        signal oVar3S40: std_logic_vector(   0 downto 0);
        signal oVar3S41: std_logic_vector(   0 downto 0);
        signal oVar3S42: std_logic_vector(   0 downto 0);
        signal oVar3S43: std_logic_vector(   0 downto 0);
        signal oVar3S44: std_logic_vector(   0 downto 0);
        signal oVar3S45: std_logic_vector(   0 downto 0);
        signal oVar3S46: std_logic_vector(   0 downto 0);
        signal oVar3S47: std_logic_vector(   0 downto 0);
        signal oVar3S48: std_logic_vector(   0 downto 0);
        signal oVar3S49: std_logic_vector(   0 downto 0);
        signal oVar3S50: std_logic_vector(   0 downto 0);
        signal oVar3S51: std_logic_vector(   0 downto 0);
        signal oVar3S52: std_logic_vector(   0 downto 0);
        signal oVar3S53: std_logic_vector(   0 downto 0);
        signal oVar3S54: std_logic_vector(   0 downto 0);
        signal oVar3S55: std_logic_vector(   0 downto 0);
        signal oVar3S56: std_logic_vector(   0 downto 0);
        signal oVar3S57: std_logic_vector(   0 downto 0);
        signal oVar3S58: std_logic_vector(   0 downto 0);
        signal oVar3S59: std_logic_vector(   0 downto 0);
        signal oVar3S60: std_logic_vector(   0 downto 0);
        signal oVar3S61: std_logic_vector(   0 downto 0);
        signal oVar3S62: std_logic_vector(   0 downto 0);
        signal oVar3S63: std_logic_vector(   0 downto 0);
        signal oVar3S64: std_logic_vector(   0 downto 0);
        signal oVar3S65: std_logic_vector(   0 downto 0);
        signal oVar3S66: std_logic_vector(   0 downto 0);
        signal oVar3S67: std_logic_vector(   0 downto 0);
        signal oVar3S68: std_logic_vector(   0 downto 0);
        signal oVar3S69: std_logic_vector(   0 downto 0);
        signal oVar3S70: std_logic_vector(   0 downto 0);
        signal oVar3S71: std_logic_vector(   0 downto 0);
        signal oVar3S72: std_logic_vector(   0 downto 0);
        signal oVar3S73: std_logic_vector(   0 downto 0);
        signal oVar3S74: std_logic_vector(   0 downto 0);
        signal oVar3S75: std_logic_vector(   0 downto 0);
        signal oVar3S76: std_logic_vector(   0 downto 0);
        signal oVar3S77: std_logic_vector(   0 downto 0);
        signal oVar3S78: std_logic_vector(   0 downto 0);
        signal oVar3S79: std_logic_vector(   0 downto 0);
        signal oVar3S80: std_logic_vector(   0 downto 0);
        signal oVar3S81: std_logic_vector(   0 downto 0);
        signal oVar3S82: std_logic_vector(   0 downto 0);
        signal oVar3S83: std_logic_vector(   0 downto 0);
        signal oVar3S84: std_logic_vector(   0 downto 0);
        signal oVar3S85: std_logic_vector(   0 downto 0);
        signal oVar3S86: std_logic_vector(   0 downto 0);
        signal oVar3S87: std_logic_vector(   0 downto 0);
        signal oVar3S88: std_logic_vector(   0 downto 0);
        signal oVar3S89: std_logic_vector(   0 downto 0);
        signal oVar3S90: std_logic_vector(   0 downto 0);
        signal oVar3S91: std_logic_vector(   0 downto 0);
        signal oVar3S92: std_logic_vector(   0 downto 0);
        signal oVar3S93: std_logic_vector(   0 downto 0);
        signal oVar3S94: std_logic_vector(   0 downto 0);
        signal oVar3S95: std_logic_vector(   0 downto 0);
        signal oVar3S96: std_logic_vector(   0 downto 0);
        signal oVar3S97: std_logic_vector(   0 downto 0);
        signal oVar3S98: std_logic_vector(   0 downto 0);
        signal oVar3S99: std_logic_vector(   0 downto 0);
        signal oVar3S100: std_logic_vector(   0 downto 0);
        signal oVar3S101: std_logic_vector(   0 downto 0);
        signal oVar3S102: std_logic_vector(   0 downto 0);
        signal oVar3S103: std_logic_vector(   0 downto 0);
        signal oVar3S104: std_logic_vector(   0 downto 0);
        signal oVar3S105: std_logic_vector(   0 downto 0);
        signal oVar3S106: std_logic_vector(   0 downto 0);
        signal oVar3S107: std_logic_vector(   0 downto 0);
        signal oVar3S108: std_logic_vector(   0 downto 0);
        signal oVar3S109: std_logic_vector(   0 downto 0);
        signal oVar3S110: std_logic_vector(   0 downto 0);
        signal oVar3S111: std_logic_vector(   0 downto 0);
        signal oVar3S112: std_logic_vector(   0 downto 0);
        signal oVar3S113: std_logic_vector(   0 downto 0);
        signal oVar3S114: std_logic_vector(   0 downto 0);
        signal oVar3S115: std_logic_vector(   0 downto 0);
        signal oVar3S116: std_logic_vector(   0 downto 0);
        signal oVar3S117: std_logic_vector(   0 downto 0);
        signal oVar3S118: std_logic_vector(   0 downto 0);
        signal oVar3S119: std_logic_vector(   0 downto 0);
        signal oVar3S120: std_logic_vector(   0 downto 0);
        signal oVar3S121: std_logic_vector(   0 downto 0);
        signal aVar3S0: std_logic_vector(   15 downto 0);
        signal aVar3S1: std_logic_vector(   15 downto 0);
        signal aVar3S2: std_logic_vector(   15 downto 0);
        signal aVar3S3: std_logic_vector(   15 downto 0);
        signal aVar3S4: std_logic_vector(   15 downto 0);
        signal aVar3S5: std_logic_vector(   15 downto 0);
        signal aVar3S6: std_logic_vector(   15 downto 0);
        signal aVar3S7: std_logic_vector(   15 downto 0);
        signal aVar3S8: std_logic_vector(   15 downto 0);
        signal aVar3S9: std_logic_vector(   15 downto 0);
        signal aVar3S10: std_logic_vector(   15 downto 0);
        signal aVar3S11: std_logic_vector(   15 downto 0);
        signal aVar3S12: std_logic_vector(   15 downto 0);
        signal aVar3S13: std_logic_vector(   15 downto 0);
        signal aVar3S14: std_logic_vector(   15 downto 0);
        signal aVar3S15: std_logic_vector(   15 downto 0);
        signal aVar4S0: std_logic_vector(   15 downto 0);
        signal aVar4S1: std_logic_vector(   15 downto 0);
        signal aVar4S2: std_logic_vector(   15 downto 0);
        signal aVar4S3: std_logic_vector(   15 downto 0);
        signal aVar4S4: std_logic_vector(   15 downto 0);
        signal aVar4S5: std_logic_vector(   15 downto 0);
        signal aVar4S6: std_logic_vector(   15 downto 0);
        signal aVar4S7: std_logic_vector(   15 downto 0);
        signal aVar5S0: std_logic_vector(   15 downto 0);
        signal aVar5S1: std_logic_vector(   15 downto 0);
        signal aVar5S2: std_logic_vector(   15 downto 0);
        signal aVar5S3: std_logic_vector(   15 downto 0);
        signal aVar6S0: std_logic_vector(   15 downto 0);
        signal aVar6S1: std_logic_vector(   15 downto 0);
        signal aVar7S0: std_logic_vector(   15 downto 0);
signal ADDM4K3S1: std_logic_vector(   7 downto 0);
signal ADDM4K3S0: std_logic_vector(   7 downto 0);
signal ADDM4K3S3: std_logic_vector(   7 downto 0);
signal ADDM4K3S2: std_logic_vector(   7 downto 0);
signal ADDM4K3S5: std_logic_vector(   7 downto 0);
signal ADDM4K3S4: std_logic_vector(   7 downto 0);
signal ADDM4K3S7: std_logic_vector(   7 downto 0);
signal ADDM4K3S6: std_logic_vector(   7 downto 0);
signal ADDM4K3S9: std_logic_vector(   7 downto 0);
signal ADDM4K3S8: std_logic_vector(   7 downto 0);
signal ADDM4K3S11: std_logic_vector(   7 downto 0);
signal ADDM4K3S10: std_logic_vector(   7 downto 0);
signal ADDM4K3S13: std_logic_vector(   7 downto 0);
signal ADDM4K3S12: std_logic_vector(   7 downto 0);
signal ADDM4K3S15: std_logic_vector(   7 downto 0);
signal ADDM4K3S14: std_logic_vector(   7 downto 0);
BEGIN
	A (19 downto 0) <= A_DIN_L (19 downto 0);
	B (8 downto 0) <= A_DIN_L (28 downto 20);
	B (17 downto 9) <= B_DIN_L (8 downto 0);
	D (15 downto 0) <= B_DIN_L (24 downto 9);
	E (15 downto 0) <= D_DIN_L (31 downto 16);
	C_DOUT_L (15 downto 0) <= output (15 downto 0);
lookuptable_LV1 : process(c1)
begin
 if c1'event and c1='1' then
        if(E( 8)='1' AND E(16)='1' AND A(23)='0' AND A(25)='0' )then
          cVar1S0S0P068P069P012P008(0) <='1';
          else
          cVar1S0S0P068P069P012P008(0) <='0';
          end if;
        if(E( 8)='1' AND E(16)='1' AND A(23)='0' AND A(25)='0' )then
          cVar1S1S0P068P069P012P008(0) <='1';
          else
          cVar1S1S0P068P069P012P008(0) <='0';
          end if;
        if(E( 8)='1' AND E(16)='0' AND E(17)='1' AND A(23)='0' )then
          cVar1S2S0P068N069P065P012(0) <='1';
          else
          cVar1S2S0P068N069P065P012(0) <='0';
          end if;
        if(E( 8)='1' AND E(16)='0' AND E(17)='0' AND D(19)='1' )then
          cVar1S3S0P068N069N065P055(0) <='1';
          else
          cVar1S3S0P068N069N065P055(0) <='0';
          end if;
        if(E( 8)='1' AND E(16)='0' AND E(17)='0' AND D(19)='1' )then
          cVar1S4S0P068N069N065P055(0) <='1';
          else
          cVar1S4S0P068N069N065P055(0) <='0';
          end if;
        if(E( 8)='1' AND E(16)='0' AND E(17)='0' AND D(19)='0' )then
          cVar1S5S0P068N069N065N055(0) <='1';
          else
          cVar1S5S0P068N069N065N055(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='1' AND E(17)='1' )then
          cVar1S6S0N068P064P063P065(0) <='1';
          else
          cVar1S6S0N068P064P063P065(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='0' AND B(11)='1' )then
          cVar1S7S0N068P064N063P035(0) <='1';
          else
          cVar1S7S0N068P064N063P035(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='0' AND B(11)='1' )then
          cVar1S8S0N068P064N063P035(0) <='1';
          else
          cVar1S8S0N068P064N063P035(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='0' AND B(11)='1' )then
          cVar1S9S0N068P064N063P035(0) <='1';
          else
          cVar1S9S0N068P064N063P035(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='0' AND B(11)='0' )then
          cVar1S10S0N068P064N063N035(0) <='1';
          else
          cVar1S10S0N068P064N063N035(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='1' AND D(17)='0' AND B(11)='0' )then
          cVar1S11S0N068P064N063N035(0) <='1';
          else
          cVar1S11S0N068P064N063N035(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='1' AND A(22)='0' )then
          cVar1S12S0N068N064P067P014(0) <='1';
          else
          cVar1S12S0N068N064P067P014(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='1' AND A(22)='1' )then
          cVar1S13S0N068N064P067P014(0) <='1';
          else
          cVar1S13S0N068N064P067P014(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='0' AND D(18)='1' )then
          cVar1S14S0N068N064N067P059(0) <='1';
          else
          cVar1S14S0N068N064N067P059(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='0' AND D(18)='1' )then
          cVar1S15S0N068N064N067P059(0) <='1';
          else
          cVar1S15S0N068N064N067P059(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='0' AND D(18)='0' )then
          cVar1S16S0N068N064N067N059(0) <='1';
          else
          cVar1S16S0N068N064N067N059(0) <='0';
          end if;
        if(E( 8)='0' AND E( 9)='0' AND D(16)='0' AND D(18)='0' )then
          cVar1S17S0N068N064N067N059(0) <='1';
          else
          cVar1S17S0N068N064N067N059(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='0' AND E(16)='1' )then
          cVar1S0S1P067P010P068P069(0) <='1';
          else
          cVar1S0S1P067P010P068P069(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='0' AND E(16)='1' )then
          cVar1S1S1P067P010P068P069(0) <='1';
          else
          cVar1S1S1P067P010P068P069(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='0' AND E(16)='0' )then
          cVar1S2S1P067P010P068N069(0) <='1';
          else
          cVar1S2S1P067P010P068N069(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='0' AND E(16)='0' )then
          cVar1S3S1P067P010P068N069(0) <='1';
          else
          cVar1S3S1P067P010P068N069(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='1' AND A(23)='1' )then
          cVar1S4S1P067P010P068P012(0) <='1';
          else
          cVar1S4S1P067P010P068P012(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='1' AND A(23)='0' )then
          cVar1S5S1P067P010P068N012(0) <='1';
          else
          cVar1S5S1P067P010P068N012(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='0' AND E( 8)='1' AND A(23)='0' )then
          cVar1S6S1P067P010P068N012(0) <='1';
          else
          cVar1S6S1P067P010P068N012(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='1' AND B(26)='0' AND B(24)='1' )then
          cVar1S7S1P067P010P024P028nsss(0) <='1';
          else
          cVar1S7S1P067P010P024P028nsss(0) <='0';
          end if;
        if(D(16)='1' AND A(24)='1' AND B(26)='0' AND B(24)='0' )then
          cVar1S8S1P067P010P024N028(0) <='1';
          else
          cVar1S8S1P067P010P024N028(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='0' AND D(17)='0' )then
          cVar1S9S1N067P068P014P063(0) <='1';
          else
          cVar1S9S1N067P068P014P063(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='0' AND D(17)='1' )then
          cVar1S10S1N067P068P014P063(0) <='1';
          else
          cVar1S10S1N067P068P014P063(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='0' AND D(17)='1' )then
          cVar1S11S1N067P068P014P063(0) <='1';
          else
          cVar1S11S1N067P068P014P063(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='0' AND D(17)='1' )then
          cVar1S12S1N067P068P014P063(0) <='1';
          else
          cVar1S12S1N067P068P014P063(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='1' AND D( 8)='1' )then
          cVar1S13S1N067P068P014P066(0) <='1';
          else
          cVar1S13S1N067P068P014P066(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='1' AND D( 8)='1' )then
          cVar1S14S1N067P068P014P066(0) <='1';
          else
          cVar1S14S1N067P068P014P066(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='1' AND D( 8)='1' )then
          cVar1S15S1N067P068P014P066(0) <='1';
          else
          cVar1S15S1N067P068P014P066(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='1' AND A(22)='1' AND D( 8)='0' )then
          cVar1S16S1N067P068P014N066(0) <='1';
          else
          cVar1S16S1N067P068P014N066(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='1' AND B(23)='1' )then
          cVar1S17S1N067N068P055P030nsss(0) <='1';
          else
          cVar1S17S1N067N068P055P030nsss(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='1' AND B(23)='0' )then
          cVar1S18S1N067N068P055N030(0) <='1';
          else
          cVar1S18S1N067N068P055N030(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='1' AND B(23)='0' )then
          cVar1S19S1N067N068P055N030(0) <='1';
          else
          cVar1S19S1N067N068P055N030(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='1' AND B(23)='0' )then
          cVar1S20S1N067N068P055N030(0) <='1';
          else
          cVar1S20S1N067N068P055N030(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='1' )then
          cVar1S21S1N067N068N055P052(0) <='1';
          else
          cVar1S21S1N067N068N055P052(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='1' )then
          cVar1S22S1N067N068N055P052(0) <='1';
          else
          cVar1S22S1N067N068N055P052(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='1' )then
          cVar1S23S1N067N068N055P052(0) <='1';
          else
          cVar1S23S1N067N068N055P052(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='0' )then
          cVar1S24S1N067N068N055N052(0) <='1';
          else
          cVar1S24S1N067N068N055N052(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='0' )then
          cVar1S25S1N067N068N055N052(0) <='1';
          else
          cVar1S25S1N067N068N055N052(0) <='0';
          end if;
        if(D(16)='0' AND E( 8)='0' AND D(19)='0' AND E(12)='0' )then
          cVar1S26S1N067N068N055N052(0) <='1';
          else
          cVar1S26S1N067N068N055N052(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='1' AND A(29)='0' AND E(21)='1' )then
          cVar1S0S2P016P047P000P049nsss(0) <='1';
          else
          cVar1S0S2P016P047P000P049nsss(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='1' AND A(29)='0' AND E(21)='0' )then
          cVar1S1S2P016P047P000N049(0) <='1';
          else
          cVar1S1S2P016P047P000N049(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='1' AND A(29)='0' AND E(21)='0' )then
          cVar1S2S2P016P047P000N049(0) <='1';
          else
          cVar1S2S2P016P047P000N049(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='1' AND B(14)='1' )then
          cVar1S3S2P016N047P052P029nsss(0) <='1';
          else
          cVar1S3S2P016N047P052P029nsss(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='1' AND B(14)='0' )then
          cVar1S4S2P016N047P052N029(0) <='1';
          else
          cVar1S4S2P016N047P052N029(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='1' )then
          cVar1S5S2P016N047N052P060(0) <='1';
          else
          cVar1S5S2P016N047N052P060(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='1' )then
          cVar1S6S2P016N047N052P060(0) <='1';
          else
          cVar1S6S2P016N047N052P060(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='1' )then
          cVar1S7S2P016N047N052P060(0) <='1';
          else
          cVar1S7S2P016N047N052P060(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='0' )then
          cVar1S8S2P016N047N052N060(0) <='1';
          else
          cVar1S8S2P016N047N052N060(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='0' )then
          cVar1S9S2P016N047N052N060(0) <='1';
          else
          cVar1S9S2P016N047N052N060(0) <='0';
          end if;
        if(A(21)='0' AND D(21)='0' AND E(12)='0' AND E(10)='0' )then
          cVar1S10S2P016N047N052N060(0) <='1';
          else
          cVar1S10S2P016N047N052N060(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='1' AND A(20)='0' )then
          cVar1S11S2P016P014P063P018(0) <='1';
          else
          cVar1S11S2P016P014P063P018(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='1' AND A(20)='0' )then
          cVar1S12S2P016P014P063P018(0) <='1';
          else
          cVar1S12S2P016P014P063P018(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='1' AND A(20)='1' )then
          cVar1S13S2P016P014P063P018(0) <='1';
          else
          cVar1S13S2P016P014P063P018(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='1' AND A(20)='1' )then
          cVar1S14S2P016P014P063P018(0) <='1';
          else
          cVar1S14S2P016P014P063P018(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='1' AND A(20)='1' )then
          cVar1S15S2P016P014P063P018(0) <='1';
          else
          cVar1S15S2P016P014P063P018(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='0' AND E(10)='1' )then
          cVar1S16S2P016P014N063P060(0) <='1';
          else
          cVar1S16S2P016P014N063P060(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='0' AND E(10)='1' )then
          cVar1S17S2P016P014N063P060(0) <='1';
          else
          cVar1S17S2P016P014N063P060(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='0' AND E(10)='0' )then
          cVar1S18S2P016P014N063N060(0) <='1';
          else
          cVar1S18S2P016P014N063N060(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='0' AND D(17)='0' AND E(10)='0' )then
          cVar1S19S2P016P014N063N060(0) <='1';
          else
          cVar1S19S2P016P014N063N060(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='1' AND A(25)='0' AND A(24)='0' )then
          cVar1S20S2P016P014P008P010(0) <='1';
          else
          cVar1S20S2P016P014P008P010(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='1' AND A(25)='0' AND A(24)='0' )then
          cVar1S21S2P016P014P008P010(0) <='1';
          else
          cVar1S21S2P016P014P008P010(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='1' AND A(25)='0' AND A(24)='0' )then
          cVar1S22S2P016P014P008P010(0) <='1';
          else
          cVar1S22S2P016P014P008P010(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='1' AND A(25)='0' AND A(24)='1' )then
          cVar1S23S2P016P014P008P010(0) <='1';
          else
          cVar1S23S2P016P014P008P010(0) <='0';
          end if;
        if(A(21)='1' AND A(22)='1' AND A(25)='1' AND A(27)='0' )then
          cVar1S24S2P016P014P008P004(0) <='1';
          else
          cVar1S24S2P016P014P008P004(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='1' AND E( 9)='0' AND A(22)='0' )then
          cVar1S0S3P047P049P064P014nsss(0) <='1';
          else
          cVar1S0S3P047P049P064P014nsss(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='1' AND E( 9)='0' AND A(22)='1' )then
          cVar1S1S3P047P049P064P014(0) <='1';
          else
          cVar1S1S3P047P049P064P014(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='1' AND E( 9)='1' )then
          cVar1S2S3P047P049P064psss(0) <='1';
          else
          cVar1S2S3P047P049P064psss(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='0' AND B(21)='0' AND D(17)='0' )then
          cVar1S3S3P047N049P034P063nsss(0) <='1';
          else
          cVar1S3S3P047N049P034P063nsss(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='1' AND B(14)='1' )then
          cVar1S4S3N047P052P029nsss(0) <='1';
          else
          cVar1S4S3N047P052P029nsss(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='1' AND B(14)='0' AND B(15)='1' )then
          cVar1S5S3N047P052N029P027nsss(0) <='1';
          else
          cVar1S5S3N047P052N029P027nsss(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S6S3N047P052N029N027(0) <='1';
          else
          cVar1S6S3N047P052N029N027(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S7S3N047P052N029N027(0) <='1';
          else
          cVar1S7S3N047P052N029N027(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='1' AND B(14)='0' AND B(15)='0' )then
          cVar1S8S3N047P052N029N027(0) <='1';
          else
          cVar1S8S3N047P052N029N027(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='1' AND E(17)='0' )then
          cVar1S9S3N047N052P060P065(0) <='1';
          else
          cVar1S9S3N047N052P060P065(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='1' AND E(17)='0' )then
          cVar1S10S3N047N052P060P065(0) <='1';
          else
          cVar1S10S3N047N052P060P065(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='1' AND E(17)='1' )then
          cVar1S11S3N047N052P060P065(0) <='1';
          else
          cVar1S11S3N047N052P060P065(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='0' )then
          cVar1S12S3N047N052N060P014(0) <='1';
          else
          cVar1S12S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='0' )then
          cVar1S13S3N047N052N060P014(0) <='1';
          else
          cVar1S13S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='0' )then
          cVar1S14S3N047N052N060P014(0) <='1';
          else
          cVar1S14S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='0' )then
          cVar1S15S3N047N052N060P014(0) <='1';
          else
          cVar1S15S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='1' )then
          cVar1S16S3N047N052N060P014(0) <='1';
          else
          cVar1S16S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='1' )then
          cVar1S17S3N047N052N060P014(0) <='1';
          else
          cVar1S17S3N047N052N060P014(0) <='0';
          end if;
        if(D(21)='0' AND E(12)='0' AND E(10)='0' AND A(22)='1' )then
          cVar1S18S3N047N052N060P014(0) <='1';
          else
          cVar1S18S3N047N052N060P014(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='1' AND A(26)='0' AND A(24)='0' )then
          cVar1S0S4P014P069P006P010(0) <='1';
          else
          cVar1S0S4P014P069P006P010(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='1' AND A(26)='0' AND A(24)='0' )then
          cVar1S1S4P014P069P006P010(0) <='1';
          else
          cVar1S1S4P014P069P006P010(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='1' AND A(26)='0' AND A(24)='1' )then
          cVar1S2S4P014P069P006P010(0) <='1';
          else
          cVar1S2S4P014P069P006P010(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='1' AND A(26)='0' AND A(24)='1' )then
          cVar1S3S4P014P069P006P010(0) <='1';
          else
          cVar1S3S4P014P069P006P010(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='1' AND A(26)='1' AND A(13)='0' )then
          cVar1S4S4P014P069P006P013(0) <='1';
          else
          cVar1S4S4P014P069P006P013(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='1' AND D(20)='1' )then
          cVar1S5S4P014N069P053P051(0) <='1';
          else
          cVar1S5S4P014N069P053P051(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='1' AND D(20)='1' )then
          cVar1S6S4P014N069P053P051(0) <='1';
          else
          cVar1S6S4P014N069P053P051(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='1' AND D(20)='0' )then
          cVar1S7S4P014N069P053N051(0) <='1';
          else
          cVar1S7S4P014N069P053N051(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='1' )then
          cVar1S8S4P014N069N053P045(0) <='1';
          else
          cVar1S8S4P014N069N053P045(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='1' )then
          cVar1S9S4P014N069N053P045(0) <='1';
          else
          cVar1S9S4P014N069N053P045(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='1' )then
          cVar1S10S4P014N069N053P045(0) <='1';
          else
          cVar1S10S4P014N069N053P045(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='0' )then
          cVar1S11S4P014N069N053N045(0) <='1';
          else
          cVar1S11S4P014N069N053N045(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='0' )then
          cVar1S12S4P014N069N053N045(0) <='1';
          else
          cVar1S12S4P014N069N053N045(0) <='0';
          end if;
        if(A(22)='0' AND E(16)='0' AND E(20)='0' AND E(22)='0' )then
          cVar1S13S4P014N069N053N045(0) <='1';
          else
          cVar1S13S4P014N069N053N045(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='1' AND A(24)='0' )then
          cVar1S14S4P014P024P060P010(0) <='1';
          else
          cVar1S14S4P014P024P060P010(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='1' AND A(24)='0' )then
          cVar1S15S4P014P024P060P010(0) <='1';
          else
          cVar1S15S4P014P024P060P010(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='1' AND A(24)='1' )then
          cVar1S16S4P014P024P060P010(0) <='1';
          else
          cVar1S16S4P014P024P060P010(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='1' )then
          cVar1S17S4P014P024N060P029(0) <='1';
          else
          cVar1S17S4P014P024N060P029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='1' )then
          cVar1S18S4P014P024N060P029(0) <='1';
          else
          cVar1S18S4P014P024N060P029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='1' )then
          cVar1S19S4P014P024N060P029(0) <='1';
          else
          cVar1S19S4P014P024N060P029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='0' )then
          cVar1S20S4P014P024N060N029(0) <='1';
          else
          cVar1S20S4P014P024N060N029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='0' )then
          cVar1S21S4P014P024N060N029(0) <='1';
          else
          cVar1S21S4P014P024N060N029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(10)='0' AND B(14)='0' )then
          cVar1S22S4P014P024N060N029(0) <='1';
          else
          cVar1S22S4P014P024N060N029(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND D(21)='1' )then
          cVar1S23S4P014P024P047nsss(0) <='1';
          else
          cVar1S23S4P014P024P047nsss(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND D(21)='0' AND E(22)='1' )then
          cVar1S24S4P014P024N047P045nsss(0) <='1';
          else
          cVar1S24S4P014P024N047P045nsss(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='1' AND B(26)='0' AND B(24)='1' )then
          cVar1S0S5P053P051P024P028nsss(0) <='1';
          else
          cVar1S0S5P053P051P024P028nsss(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='1' AND B(26)='0' AND B(24)='0' )then
          cVar1S1S5P053P051P024N028(0) <='1';
          else
          cVar1S1S5P053P051P024N028(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='1' AND B(26)='0' AND B(24)='0' )then
          cVar1S2S5P053P051P024N028(0) <='1';
          else
          cVar1S2S5P053P051P024N028(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='1' AND B(26)='0' AND B(24)='0' )then
          cVar1S3S5P053P051P024N028(0) <='1';
          else
          cVar1S3S5P053P051P024N028(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='0' AND A(24)='0' AND D(21)='1' )then
          cVar1S4S5P053N051P010P047nsss(0) <='1';
          else
          cVar1S4S5P053N051P010P047nsss(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='0' AND A(24)='0' AND D(21)='0' )then
          cVar1S5S5P053N051P010N047(0) <='1';
          else
          cVar1S5S5P053N051P010N047(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='0' AND A(24)='0' AND D(21)='0' )then
          cVar1S6S5P053N051P010N047(0) <='1';
          else
          cVar1S6S5P053N051P010N047(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='0' AND A(24)='0' AND D(21)='0' )then
          cVar1S7S5P053N051P010N047(0) <='1';
          else
          cVar1S7S5P053N051P010N047(0) <='0';
          end if;
        if(E(20)='1' AND D(20)='0' AND A(24)='1' AND D(19)='1' )then
          cVar1S8S5P053N051P010P055nsss(0) <='1';
          else
          cVar1S8S5P053N051P010P055nsss(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='1' AND A(24)='0' )then
          cVar1S9S5N053P051P069P010(0) <='1';
          else
          cVar1S9S5N053P051P069P010(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='1' AND A(24)='0' )then
          cVar1S10S5N053P051P069P010(0) <='1';
          else
          cVar1S10S5N053P051P069P010(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='1' AND A(24)='0' )then
          cVar1S11S5N053P051P069P010(0) <='1';
          else
          cVar1S11S5N053P051P069P010(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='1' AND A(24)='1' )then
          cVar1S12S5N053P051P069P010(0) <='1';
          else
          cVar1S12S5N053P051P069P010(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='1' AND A(24)='1' )then
          cVar1S13S5N053P051P069P010(0) <='1';
          else
          cVar1S13S5N053P051P069P010(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='0' AND E(22)='1' )then
          cVar1S14S5N053P051N069P045(0) <='1';
          else
          cVar1S14S5N053P051N069P045(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='0' AND E(22)='1' )then
          cVar1S15S5N053P051N069P045(0) <='1';
          else
          cVar1S15S5N053P051N069P045(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='0' AND E(22)='0' )then
          cVar1S16S5N053P051N069N045(0) <='1';
          else
          cVar1S16S5N053P051N069N045(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='0' AND E(22)='0' )then
          cVar1S17S5N053P051N069N045(0) <='1';
          else
          cVar1S17S5N053P051N069N045(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='0' AND E(16)='0' AND E(22)='0' )then
          cVar1S18S5N053P051N069N045(0) <='1';
          else
          cVar1S18S5N053P051N069N045(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='1' AND E(21)='1' AND E(18)='0' )then
          cVar1S19S5N053P051P049P061(0) <='1';
          else
          cVar1S19S5N053P051P049P061(0) <='0';
          end if;
        if(E(20)='0' AND D(20)='1' AND E(21)='0' AND A(12)='0' )then
          cVar1S20S5N053P051N049P015(0) <='1';
          else
          cVar1S20S5N053P051N049P015(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='1' AND E( 9)='0' AND A(23)='0' )then
          cVar1S0S6P047P049P064P012nsss(0) <='1';
          else
          cVar1S0S6P047P049P064P012nsss(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='1' AND E( 9)='0' AND A(23)='1' )then
          cVar1S1S6P047P049P064P012(0) <='1';
          else
          cVar1S1S6P047P049P064P012(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='0' AND B(21)='0' AND B(11)='0' )then
          cVar1S2S6P047N049P034P035(0) <='1';
          else
          cVar1S2S6P047N049P034P035(0) <='0';
          end if;
        if(D(21)='1' AND E(21)='0' AND B(21)='0' AND B(11)='0' )then
          cVar1S3S6P047N049P034P035(0) <='1';
          else
          cVar1S3S6P047N049P034P035(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='1' AND B(23)='1' )then
          cVar1S4S6N047P024P055P030(0) <='1';
          else
          cVar1S4S6N047P024P055P030(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='1' AND B(23)='0' )then
          cVar1S5S6N047P024P055N030(0) <='1';
          else
          cVar1S5S6N047P024P055N030(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='1' AND B(23)='0' )then
          cVar1S6S6N047P024P055N030(0) <='1';
          else
          cVar1S6S6N047P024P055N030(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='0' AND E(20)='1' )then
          cVar1S7S6N047P024N055P053(0) <='1';
          else
          cVar1S7S6N047P024N055P053(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='0' AND E(20)='1' )then
          cVar1S8S6N047P024N055P053(0) <='1';
          else
          cVar1S8S6N047P024N055P053(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='0' AND D(19)='0' AND E(20)='0' )then
          cVar1S9S6N047P024N055N053(0) <='1';
          else
          cVar1S9S6N047P024N055N053(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='1' AND B(22)='0' AND E(22)='1' )then
          cVar1S10S6N047P024P032P045(0) <='1';
          else
          cVar1S10S6N047P024P032P045(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='1' AND B(22)='0' AND E(22)='0' )then
          cVar1S11S6N047P024P032N045(0) <='1';
          else
          cVar1S11S6N047P024P032N045(0) <='0';
          end if;
        if(D(21)='0' AND B(26)='1' AND B(22)='0' AND E(22)='0' )then
          cVar1S12S6N047P024P032N045(0) <='1';
          else
          cVar1S12S6N047P024P032N045(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='1' )then
          cVar1S0S7P053P006P028nsss(0) <='1';
          else
          cVar1S0S7P053P006P028nsss(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='1' )then
          cVar1S1S7P053P006N028P029nsss(0) <='1';
          else
          cVar1S1S7P053P006N028P029nsss(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S2S7P053P006N028N029(0) <='1';
          else
          cVar1S2S7P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S3S7P053P006N028N029(0) <='1';
          else
          cVar1S3S7P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S4S7P053P006N028N029(0) <='1';
          else
          cVar1S4S7P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='1' AND D(17)='0' AND A(11)='0' )then
          cVar1S5S7P053P006P063P017(0) <='1';
          else
          cVar1S5S7P053P006P063P017(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='1' AND B(23)='1' AND E(19)='1' )then
          cVar1S6S7N053P055P030P057(0) <='1';
          else
          cVar1S6S7N053P055P030P057(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='1' AND B(23)='1' AND E(19)='1' )then
          cVar1S7S7N053P055P030P057(0) <='1';
          else
          cVar1S7S7N053P055P030P057(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='1' AND B(23)='0' AND E( 8)='0' )then
          cVar1S8S7N053P055N030P068(0) <='1';
          else
          cVar1S8S7N053P055N030P068(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='1' AND B(23)='0' AND E( 8)='0' )then
          cVar1S9S7N053P055N030P068(0) <='1';
          else
          cVar1S9S7N053P055N030P068(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='1' AND B(23)='0' AND E( 8)='1' )then
          cVar1S10S7N053P055N030P068(0) <='1';
          else
          cVar1S10S7N053P055N030P068(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='1' AND E(21)='1' )then
          cVar1S11S7N053N055P047P049nsss(0) <='1';
          else
          cVar1S11S7N053N055P047P049nsss(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='1' AND E(21)='0' )then
          cVar1S12S7N053N055P047N049(0) <='1';
          else
          cVar1S12S7N053N055P047N049(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='1' AND E(21)='0' )then
          cVar1S13S7N053N055P047N049(0) <='1';
          else
          cVar1S13S7N053N055P047N049(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='1' )then
          cVar1S14S7N053N055N047P033(0) <='1';
          else
          cVar1S14S7N053N055N047P033(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='1' )then
          cVar1S15S7N053N055N047P033(0) <='1';
          else
          cVar1S15S7N053N055N047P033(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='1' )then
          cVar1S16S7N053N055N047P033(0) <='1';
          else
          cVar1S16S7N053N055N047P033(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='0' )then
          cVar1S17S7N053N055N047N033(0) <='1';
          else
          cVar1S17S7N053N055N047N033(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='0' )then
          cVar1S18S7N053N055N047N033(0) <='1';
          else
          cVar1S18S7N053N055N047N033(0) <='0';
          end if;
        if(E(20)='0' AND D(19)='0' AND D(21)='0' AND B(12)='0' )then
          cVar1S19S7N053N055N047N033(0) <='1';
          else
          cVar1S19S7N053N055N047N033(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='1' AND A(29)='0' AND B(24)='1' )then
          cVar1S0S8P036P053P000P028nsss(0) <='1';
          else
          cVar1S0S8P036P053P000P028nsss(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='1' AND A(29)='0' AND B(24)='0' )then
          cVar1S1S8P036P053P000N028(0) <='1';
          else
          cVar1S1S8P036P053P000N028(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='1' AND A(29)='0' AND B(24)='0' )then
          cVar1S2S8P036P053P000N028(0) <='1';
          else
          cVar1S2S8P036P053P000N028(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='1' AND A(29)='0' AND B(24)='0' )then
          cVar1S3S8P036P053P000N028(0) <='1';
          else
          cVar1S3S8P036P053P000N028(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S4S8P036N053P046P025nsss(0) <='1';
          else
          cVar1S4S8P036N053P046P025nsss(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S5S8P036N053P046N025(0) <='1';
          else
          cVar1S5S8P036N053P046N025(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S6S8P036N053P046N025(0) <='1';
          else
          cVar1S6S8P036N053P046N025(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S7S8P036N053P046N025(0) <='1';
          else
          cVar1S7S8P036N053P046N025(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='0' AND D(20)='0' )then
          cVar1S8S8P036N053N046P051(0) <='1';
          else
          cVar1S8S8P036N053N046P051(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='0' AND D(20)='0' )then
          cVar1S9S8P036N053N046P051(0) <='1';
          else
          cVar1S9S8P036N053N046P051(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='0' AND D(20)='0' )then
          cVar1S10S8P036N053N046P051(0) <='1';
          else
          cVar1S10S8P036N053N046P051(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='0' AND D(20)='1' )then
          cVar1S11S8P036N053N046P051(0) <='1';
          else
          cVar1S11S8P036N053N046P051(0) <='0';
          end if;
        if(B(20)='0' AND E(20)='0' AND D(13)='0' AND D(20)='1' )then
          cVar1S12S8P036N053N046P051(0) <='1';
          else
          cVar1S12S8P036N053N046P051(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='1' AND A(25)='0' )then
          cVar1S13S8P036P010P016P008(0) <='1';
          else
          cVar1S13S8P036P010P016P008(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='1' AND A(25)='0' )then
          cVar1S14S8P036P010P016P008(0) <='1';
          else
          cVar1S14S8P036P010P016P008(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='0' AND A(20)='1' )then
          cVar1S15S8P036P010N016P018(0) <='1';
          else
          cVar1S15S8P036P010N016P018(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='0' AND A(20)='1' )then
          cVar1S16S8P036P010N016P018(0) <='1';
          else
          cVar1S16S8P036P010N016P018(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='0' AND A(20)='1' )then
          cVar1S17S8P036P010N016P018(0) <='1';
          else
          cVar1S17S8P036P010N016P018(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='0' AND A(20)='0' )then
          cVar1S18S8P036P010N016N018(0) <='1';
          else
          cVar1S18S8P036P010N016N018(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='0' AND A(21)='0' AND A(20)='0' )then
          cVar1S19S8P036P010N016N018(0) <='1';
          else
          cVar1S19S8P036P010N016N018(0) <='0';
          end if;
        if(B(20)='1' AND A(24)='1' AND B(26)='0' AND A(27)='1' )then
          cVar1S20S8P036P010P024P004(0) <='1';
          else
          cVar1S20S8P036P010P024P004(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='1' )then
          cVar1S0S9P052P029nsss(0) <='1';
          else
          cVar1S0S9P052P029nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B(15)='1' )then
          cVar1S1S9P052N029P027nsss(0) <='1';
          else
          cVar1S1S9P052N029P027nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B(15)='0' AND B(24)='1' )then
          cVar1S2S9P052N029N027P028nsss(0) <='1';
          else
          cVar1S2S9P052N029N027P028nsss(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B(15)='0' AND B(24)='0' )then
          cVar1S3S9P052N029N027N028(0) <='1';
          else
          cVar1S3S9P052N029N027N028(0) <='0';
          end if;
        if(E(12)='1' AND B(14)='0' AND B(15)='0' AND B(24)='0' )then
          cVar1S4S9P052N029N027N028(0) <='1';
          else
          cVar1S4S9P052N029N027N028(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S5S9N052P046P025nsss(0) <='1';
          else
          cVar1S5S9N052P046P025nsss(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='1' AND B(16)='0' AND A(22)='0' )then
          cVar1S6S9N052P046N025P014(0) <='1';
          else
          cVar1S6S9N052P046N025P014(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='1' AND B(16)='0' AND A(22)='0' )then
          cVar1S7S9N052P046N025P014(0) <='1';
          else
          cVar1S7S9N052P046N025P014(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='1' AND B(16)='0' AND A(22)='0' )then
          cVar1S8S9N052P046N025P014(0) <='1';
          else
          cVar1S8S9N052P046N025P014(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S9S9N052N046P041P039(0) <='1';
          else
          cVar1S9S9N052N046P041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S10S9N052N046P041P039(0) <='1';
          else
          cVar1S10S9N052N046P041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S11S9N052N046P041P039(0) <='1';
          else
          cVar1S11S9N052N046P041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='1' AND D(23)='0' )then
          cVar1S12S9N052N046P041N039(0) <='1';
          else
          cVar1S12S9N052N046P041N039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S13S9N052N046N041P039(0) <='1';
          else
          cVar1S13S9N052N046N041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S14S9N052N046N041P039(0) <='1';
          else
          cVar1S14S9N052N046N041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S15S9N052N046N041P039(0) <='1';
          else
          cVar1S15S9N052N046N041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S16S9N052N046N041P039(0) <='1';
          else
          cVar1S16S9N052N046N041P039(0) <='0';
          end if;
        if(E(12)='0' AND D(13)='0' AND E(23)='0' AND D(23)='1' )then
          cVar1S17S9N052N046N041P039(0) <='1';
          else
          cVar1S17S9N052N046N041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='1' AND D(17)='0' AND B(24)='1' )then
          cVar1S0S10P012P053P063P028nsss(0) <='1';
          else
          cVar1S0S10P012P053P063P028nsss(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='1' AND D(17)='0' AND B(24)='0' )then
          cVar1S1S10P012P053P063N028(0) <='1';
          else
          cVar1S1S10P012P053P063N028(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='1' AND D(17)='0' AND B(24)='0' )then
          cVar1S2S10P012P053P063N028(0) <='1';
          else
          cVar1S2S10P012P053P063N028(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='1' AND D(17)='0' AND B(24)='0' )then
          cVar1S3S10P012P053P063N028(0) <='1';
          else
          cVar1S3S10P012P053P063N028(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='1' AND D(17)='1' AND D( 9)='0' )then
          cVar1S4S10P012P053P063P062(0) <='1';
          else
          cVar1S4S10P012P053P063P062(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S5S10P012N053P041P039(0) <='1';
          else
          cVar1S5S10P012N053P041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S6S10P012N053P041P039(0) <='1';
          else
          cVar1S6S10P012N053P041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S7S10P012N053P041P039(0) <='1';
          else
          cVar1S7S10P012N053P041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='1' AND D(23)='0' )then
          cVar1S8S10P012N053P041N039(0) <='1';
          else
          cVar1S8S10P012N053P041N039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S9S10P012N053N041P039(0) <='1';
          else
          cVar1S9S10P012N053N041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S10S10P012N053N041P039(0) <='1';
          else
          cVar1S10S10P012N053N041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S11S10P012N053N041P039(0) <='1';
          else
          cVar1S11S10P012N053N041P039(0) <='0';
          end if;
        if(A(23)='0' AND E(20)='0' AND E(23)='0' AND D(23)='1' )then
          cVar1S12S10P012N053N041P039(0) <='1';
          else
          cVar1S12S10P012N053N041P039(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='1' AND A(26)='0' AND A(22)='0' )then
          cVar1S13S10P012P030P006P014(0) <='1';
          else
          cVar1S13S10P012P030P006P014(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='1' AND A(26)='0' AND A(22)='0' )then
          cVar1S14S10P012P030P006P014(0) <='1';
          else
          cVar1S14S10P012P030P006P014(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='1' AND A(26)='0' AND A(22)='0' )then
          cVar1S15S10P012P030P006P014(0) <='1';
          else
          cVar1S15S10P012P030P006P014(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='1' AND A(26)='0' AND A(22)='1' )then
          cVar1S16S10P012P030P006P014(0) <='1';
          else
          cVar1S16S10P012P030P006P014(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='1' )then
          cVar1S17S10P012N030P008P031(0) <='1';
          else
          cVar1S17S10P012N030P008P031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='1' )then
          cVar1S18S10P012N030P008P031(0) <='1';
          else
          cVar1S18S10P012N030P008P031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='1' )then
          cVar1S19S10P012N030P008P031(0) <='1';
          else
          cVar1S19S10P012N030P008P031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='0' )then
          cVar1S20S10P012N030P008N031(0) <='1';
          else
          cVar1S20S10P012N030P008N031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='0' )then
          cVar1S21S10P012N030P008N031(0) <='1';
          else
          cVar1S21S10P012N030P008N031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='0' AND B(13)='0' )then
          cVar1S22S10P012N030P008N031(0) <='1';
          else
          cVar1S22S10P012N030P008N031(0) <='0';
          end if;
        if(A(23)='1' AND B(23)='0' AND A(25)='1' AND A(14)='0' )then
          cVar1S23S10P012N030P008P011(0) <='1';
          else
          cVar1S23S10P012N030P008P011(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='1' )then
          cVar1S0S11P053P006P028nsss(0) <='1';
          else
          cVar1S0S11P053P006P028nsss(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='1' )then
          cVar1S1S11P053P006N028P029nsss(0) <='1';
          else
          cVar1S1S11P053P006N028P029nsss(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S2S11P053P006N028N029(0) <='1';
          else
          cVar1S2S11P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S3S11P053P006N028N029(0) <='1';
          else
          cVar1S3S11P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='0' AND B(24)='0' AND B(14)='0' )then
          cVar1S4S11P053P006N028N029(0) <='1';
          else
          cVar1S4S11P053P006N028N029(0) <='0';
          end if;
        if(E(20)='1' AND A(26)='1' AND D(17)='0' AND A(11)='0' )then
          cVar1S5S11P053P006P063P017(0) <='1';
          else
          cVar1S5S11P053P006P063P017(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='1' AND B(28)='1' )then
          cVar1S6S11N053P041P020nsss(0) <='1';
          else
          cVar1S6S11N053P041P020nsss(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='1' AND B(28)='0' AND B(18)='1' )then
          cVar1S7S11N053P041N020P021nsss(0) <='1';
          else
          cVar1S7S11N053P041N020P021nsss(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='1' AND B(28)='0' AND B(18)='0' )then
          cVar1S8S11N053P041N020N021(0) <='1';
          else
          cVar1S8S11N053P041N020N021(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='1' )then
          cVar1S9S11N053N041P039P046(0) <='1';
          else
          cVar1S9S11N053N041P039P046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='1' )then
          cVar1S10S11N053N041P039P046(0) <='1';
          else
          cVar1S10S11N053N041P039P046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='1' )then
          cVar1S11S11N053N041P039P046(0) <='1';
          else
          cVar1S11S11N053N041P039P046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='0' )then
          cVar1S12S11N053N041P039N046(0) <='1';
          else
          cVar1S12S11N053N041P039N046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='0' )then
          cVar1S13S11N053N041P039N046(0) <='1';
          else
          cVar1S13S11N053N041P039N046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='0' )then
          cVar1S14S11N053N041P039N046(0) <='1';
          else
          cVar1S14S11N053N041P039N046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='0' AND D(13)='0' )then
          cVar1S15S11N053N041P039N046(0) <='1';
          else
          cVar1S15S11N053N041P039N046(0) <='0';
          end if;
        if(E(20)='0' AND E(23)='0' AND D(23)='1' AND A(25)='0' )then
          cVar1S16S11N053N041P039P008(0) <='1';
          else
          cVar1S16S11N053N041P039P008(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='1' AND A(26)='0' )then
          cVar1S0S12P015P016P037P006(0) <='1';
          else
          cVar1S0S12P015P016P037P006(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='1' AND A(26)='0' )then
          cVar1S1S12P015P016P037P006(0) <='1';
          else
          cVar1S1S12P015P016P037P006(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='1' AND A(26)='1' )then
          cVar1S2S12P015P016P037P006(0) <='1';
          else
          cVar1S2S12P015P016P037P006(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='0' AND D(17)='1' )then
          cVar1S3S12P015P016N037P063(0) <='1';
          else
          cVar1S3S12P015P016N037P063(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='0' AND D(17)='1' )then
          cVar1S4S12P015P016N037P063(0) <='1';
          else
          cVar1S4S12P015P016N037P063(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='0' AND D(17)='0' )then
          cVar1S5S12P015P016N037N063(0) <='1';
          else
          cVar1S5S12P015P016N037N063(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(10)='0' AND D(17)='0' )then
          cVar1S6S12P015P016N037N063(0) <='1';
          else
          cVar1S6S12P015P016N037N063(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='0' AND E(23)='1' )then
          cVar1S7S12P015N016P065P041(0) <='1';
          else
          cVar1S7S12P015N016P065P041(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='0' AND E(23)='1' )then
          cVar1S8S12P015N016P065P041(0) <='1';
          else
          cVar1S8S12P015N016P065P041(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='0' AND E(23)='0' )then
          cVar1S9S12P015N016P065N041(0) <='1';
          else
          cVar1S9S12P015N016P065N041(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='0' AND E(23)='0' )then
          cVar1S10S12P015N016P065N041(0) <='1';
          else
          cVar1S10S12P015N016P065N041(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='0' AND E(23)='0' )then
          cVar1S11S12P015N016P065N041(0) <='1';
          else
          cVar1S11S12P015N016P065N041(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='1' AND A(27)='0' )then
          cVar1S12S12P015N016P065P004(0) <='1';
          else
          cVar1S12S12P015N016P065P004(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='1' AND A(27)='0' )then
          cVar1S13S12P015N016P065P004(0) <='1';
          else
          cVar1S13S12P015N016P065P004(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND E(17)='1' AND A(27)='0' )then
          cVar1S14S12P015N016P065P004(0) <='1';
          else
          cVar1S14S12P015N016P065P004(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='1' AND D(17)='0' )then
          cVar1S15S12P015P016P033P063(0) <='1';
          else
          cVar1S15S12P015P016P033P063(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='1' AND D(17)='0' )then
          cVar1S16S12P015P016P033P063(0) <='1';
          else
          cVar1S16S12P015P016P033P063(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='0' AND B(11)='1' )then
          cVar1S17S12P015P016N033P035(0) <='1';
          else
          cVar1S17S12P015P016N033P035(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='0' AND B(11)='1' )then
          cVar1S18S12P015P016N033P035(0) <='1';
          else
          cVar1S18S12P015P016N033P035(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='0' AND B(11)='0' )then
          cVar1S19S12P015P016N033N035(0) <='1';
          else
          cVar1S19S12P015P016N033N035(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='0' AND B(12)='0' AND B(11)='0' )then
          cVar1S20S12P015P016N033N035(0) <='1';
          else
          cVar1S20S12P015P016N033N035(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='1' AND A(26)='0' AND A(10)='0' )then
          cVar1S21S12P015P016P006P019(0) <='1';
          else
          cVar1S21S12P015P016P006P019(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='1' AND A(26)='0' AND A(10)='0' )then
          cVar1S22S12P015P016P006P019(0) <='1';
          else
          cVar1S22S12P015P016P006P019(0) <='0';
          end if;
        if(A(12)='1' AND A(21)='1' AND A(26)='0' AND A(10)='1' )then
          cVar1S23S12P015P016P006P019(0) <='1';
          else
          cVar1S23S12P015P016P006P019(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar1S0S13P001P066P011P068(0) <='1';
          else
          cVar1S0S13P001P066P011P068(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar1S1S13P001P066P011P068(0) <='1';
          else
          cVar1S1S13P001P066P011P068(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='0' AND E( 8)='1' )then
          cVar1S2S13P001P066P011P068(0) <='1';
          else
          cVar1S2S13P001P066P011P068(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='0' AND E( 8)='0' )then
          cVar1S3S13P001P066P011N068(0) <='1';
          else
          cVar1S3S13P001P066P011N068(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='1' AND A(28)='0' )then
          cVar1S4S13P001P066P011P002(0) <='1';
          else
          cVar1S4S13P001P066P011P002(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='1' AND A(28)='0' )then
          cVar1S5S13P001P066P011P002(0) <='1';
          else
          cVar1S5S13P001P066P011P002(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='1' AND A(14)='1' AND A(28)='0' )then
          cVar1S6S13P001P066P011P002(0) <='1';
          else
          cVar1S6S13P001P066P011P002(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S7S13P001N066P027P009(0) <='1';
          else
          cVar1S7S13P001N066P027P009(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S8S13P001N066P027P009(0) <='1';
          else
          cVar1S8S13P001N066P027P009(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='1' AND A(15)='0' )then
          cVar1S9S13P001N066P027N009(0) <='1';
          else
          cVar1S9S13P001N066P027N009(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='1' AND A(15)='0' )then
          cVar1S10S13P001N066P027N009(0) <='1';
          else
          cVar1S10S13P001N066P027N009(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='1' )then
          cVar1S11S13P001N066N027P053(0) <='1';
          else
          cVar1S11S13P001N066N027P053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='1' )then
          cVar1S12S13P001N066N027P053(0) <='1';
          else
          cVar1S12S13P001N066N027P053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='1' )then
          cVar1S13S13P001N066N027P053(0) <='1';
          else
          cVar1S13S13P001N066N027P053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='0' )then
          cVar1S14S13P001N066N027N053(0) <='1';
          else
          cVar1S14S13P001N066N027N053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='0' )then
          cVar1S15S13P001N066N027N053(0) <='1';
          else
          cVar1S15S13P001N066N027N053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='0' )then
          cVar1S16S13P001N066N027N053(0) <='1';
          else
          cVar1S16S13P001N066N027N053(0) <='0';
          end if;
        if(A(19)='0' AND D( 8)='0' AND B(15)='0' AND E(20)='0' )then
          cVar1S17S13P001N066N027N053(0) <='1';
          else
          cVar1S17S13P001N066N027N053(0) <='0';
          end if;
        if(A(19)='1' AND A(26)='0' AND D(20)='0' AND A(27)='0' )then
          cVar1S18S13P001P006P051P004(0) <='1';
          else
          cVar1S18S13P001P006P051P004(0) <='0';
          end if;
        if(A(19)='1' AND A(26)='0' AND D(20)='0' AND A(27)='0' )then
          cVar1S19S13P001P006P051P004(0) <='1';
          else
          cVar1S19S13P001P006P051P004(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='1' AND D(17)='1' )then
          cVar1S0S14P015P016P034P063nsss(0) <='1';
          else
          cVar1S0S14P015P016P034P063nsss(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='1' AND D(17)='0' )then
          cVar1S1S14P015P016P034N063(0) <='1';
          else
          cVar1S1S14P015P016P034N063(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='0' AND B(10)='1' )then
          cVar1S2S14P015P016N034P037(0) <='1';
          else
          cVar1S2S14P015P016N034P037(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='0' AND B(10)='1' )then
          cVar1S3S14P015P016N034P037(0) <='1';
          else
          cVar1S3S14P015P016N034P037(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='0' AND B(10)='0' )then
          cVar1S4S14P015P016N034N037(0) <='1';
          else
          cVar1S4S14P015P016N034N037(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='0' AND B(10)='0' )then
          cVar1S5S14P015P016N034N037(0) <='1';
          else
          cVar1S5S14P015P016N034N037(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='1' AND B(21)='0' AND B(10)='0' )then
          cVar1S6S14P015P016N034N037(0) <='1';
          else
          cVar1S6S14P015P016N034N037(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S7S14P015N016P046P025nsss(0) <='1';
          else
          cVar1S7S14P015N016P046P025nsss(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S8S14P015N016P046N025(0) <='1';
          else
          cVar1S8S14P015N016P046N025(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S9S14P015N016P046N025(0) <='1';
          else
          cVar1S9S14P015N016P046N025(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='1' )then
          cVar1S10S14P015N016N046P022(0) <='1';
          else
          cVar1S10S14P015N016N046P022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='1' )then
          cVar1S11S14P015N016N046P022(0) <='1';
          else
          cVar1S11S14P015N016N046P022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='1' )then
          cVar1S12S14P015N016N046P022(0) <='1';
          else
          cVar1S12S14P015N016N046P022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='0' )then
          cVar1S13S14P015N016N046N022(0) <='1';
          else
          cVar1S13S14P015N016N046N022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='0' )then
          cVar1S14S14P015N016N046N022(0) <='1';
          else
          cVar1S14S14P015N016N046N022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='0' )then
          cVar1S15S14P015N016N046N022(0) <='1';
          else
          cVar1S15S14P015N016N046N022(0) <='0';
          end if;
        if(A(12)='0' AND A(21)='0' AND D(13)='0' AND B(27)='0' )then
          cVar1S16S14P015N016N046N022(0) <='1';
          else
          cVar1S16S14P015N016N046N022(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='0' AND B(12)='1' )then
          cVar1S17S14P015P009P016P033(0) <='1';
          else
          cVar1S17S14P015P009P016P033(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='0' AND B(12)='1' )then
          cVar1S18S14P015P009P016P033(0) <='1';
          else
          cVar1S18S14P015P009P016P033(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='0' AND B(12)='0' )then
          cVar1S19S14P015P009P016N033(0) <='1';
          else
          cVar1S19S14P015P009P016N033(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='0' AND B(12)='0' )then
          cVar1S20S14P015P009P016N033(0) <='1';
          else
          cVar1S20S14P015P009P016N033(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='1' AND A(10)='0' )then
          cVar1S21S14P015P009P016P019(0) <='1';
          else
          cVar1S21S14P015P009P016P019(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='1' AND A(10)='0' )then
          cVar1S22S14P015P009P016P019(0) <='1';
          else
          cVar1S22S14P015P009P016P019(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='1' AND A(10)='0' )then
          cVar1S23S14P015P009P016P019(0) <='1';
          else
          cVar1S23S14P015P009P016P019(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='1' AND A(10)='1' )then
          cVar1S24S14P015P009P016P019(0) <='1';
          else
          cVar1S24S14P015P009P016P019(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND A(21)='1' AND A(10)='1' )then
          cVar1S25S14P015P009P016P019(0) <='1';
          else
          cVar1S25S14P015P009P016P019(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='1' AND B(15)='1' )then
          cVar1S26S14P015P009P027nsss(0) <='1';
          else
          cVar1S26S14P015P009P027nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='1' )then
          cVar1S0S15P046P025nsss(0) <='1';
          else
          cVar1S0S15P046P025nsss(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(22)='0' AND A(22)='0' )then
          cVar1S1S15P046N025P032P014(0) <='1';
          else
          cVar1S1S15P046N025P032P014(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(22)='0' AND A(22)='0' )then
          cVar1S2S15P046N025P032P014(0) <='1';
          else
          cVar1S2S15P046N025P032P014(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(22)='0' AND A(22)='0' )then
          cVar1S3S15P046N025P032P014(0) <='1';
          else
          cVar1S3S15P046N025P032P014(0) <='0';
          end if;
        if(D(13)='1' AND B(16)='0' AND B(22)='0' AND A(22)='1' )then
          cVar1S4S15P046N025P032P014(0) <='1';
          else
          cVar1S4S15P046N025P032P014(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='0' AND B(21)='1' )then
          cVar1S5S15N046P016P018P034(0) <='1';
          else
          cVar1S5S15N046P016P018P034(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='0' AND B(21)='1' )then
          cVar1S6S15N046P016P018P034(0) <='1';
          else
          cVar1S6S15N046P016P018P034(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='0' AND B(21)='0' )then
          cVar1S7S15N046P016P018N034(0) <='1';
          else
          cVar1S7S15N046P016P018N034(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='0' AND B(21)='0' )then
          cVar1S8S15N046P016P018N034(0) <='1';
          else
          cVar1S8S15N046P016P018N034(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='0' AND B(21)='0' )then
          cVar1S9S15N046P016P018N034(0) <='1';
          else
          cVar1S9S15N046P016P018N034(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='1' AND A(10)='0' )then
          cVar1S10S15N046P016P018P019(0) <='1';
          else
          cVar1S10S15N046P016P018P019(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='1' AND A(10)='0' )then
          cVar1S11S15N046P016P018P019(0) <='1';
          else
          cVar1S11S15N046P016P018P019(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='1' AND A(20)='1' AND A(10)='1' )then
          cVar1S12S15N046P016P018P019(0) <='1';
          else
          cVar1S12S15N046P016P018P019(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='1' AND E(19)='1' )then
          cVar1S13S15N046N016P056P057nsss(0) <='1';
          else
          cVar1S13S15N046N016P056P057nsss(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='1' AND E(19)='0' )then
          cVar1S14S15N046N016P056N057(0) <='1';
          else
          cVar1S14S15N046N016P056N057(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='1' AND E(19)='0' )then
          cVar1S15S15N046N016P056N057(0) <='1';
          else
          cVar1S15S15N046N016P056N057(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='0' AND D(11)='0' )then
          cVar1S16S15N046N016N056P054(0) <='1';
          else
          cVar1S16S15N046N016N056P054(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='0' AND D(11)='0' )then
          cVar1S17S15N046N016N056P054(0) <='1';
          else
          cVar1S17S15N046N016N056P054(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='0' AND D(11)='0' )then
          cVar1S18S15N046N016N056P054(0) <='1';
          else
          cVar1S18S15N046N016N056P054(0) <='0';
          end if;
        if(D(13)='0' AND A(21)='0' AND E(11)='0' AND D(11)='1' )then
          cVar1S19S15N046N016N056P054(0) <='1';
          else
          cVar1S19S15N046N016N056P054(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='1' AND D(14)='1' )then
          cVar1S0S16P016P000P023P042nsss(0) <='1';
          else
          cVar1S0S16P016P000P023P042nsss(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='1' AND D(14)='0' )then
          cVar1S1S16P016P000P023N042(0) <='1';
          else
          cVar1S1S16P016P000P023N042(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='0' AND B(27)='1' )then
          cVar1S2S16P016P000N023P022(0) <='1';
          else
          cVar1S2S16P016P000N023P022(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='0' AND B(27)='1' )then
          cVar1S3S16P016P000N023P022(0) <='1';
          else
          cVar1S3S16P016P000N023P022(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='0' AND B(27)='0' )then
          cVar1S4S16P016P000N023N022(0) <='1';
          else
          cVar1S4S16P016P000N023N022(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND B(17)='0' AND B(27)='0' )then
          cVar1S5S16P016P000N023N022(0) <='1';
          else
          cVar1S5S16P016P000N023N022(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='1' AND E(20)='0' AND D( 9)='0' )then
          cVar1S6S16P016P000P053P062(0) <='1';
          else
          cVar1S6S16P016P000P053P062(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S7S16P016P015P034P063(0) <='1';
          else
          cVar1S7S16P016P015P034P063(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S8S16P016P015P034P063(0) <='1';
          else
          cVar1S8S16P016P015P034P063(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S9S16P016P015P034P063(0) <='1';
          else
          cVar1S9S16P016P015P034P063(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='1' AND D(17)='0' )then
          cVar1S10S16P016P015P034N063(0) <='1';
          else
          cVar1S10S16P016P015P034N063(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='0' AND B(10)='1' )then
          cVar1S11S16P016P015N034P037(0) <='1';
          else
          cVar1S11S16P016P015N034P037(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='0' AND B(10)='0' )then
          cVar1S12S16P016P015N034N037(0) <='1';
          else
          cVar1S12S16P016P015N034N037(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='0' AND B(10)='0' )then
          cVar1S13S16P016P015N034N037(0) <='1';
          else
          cVar1S13S16P016P015N034N037(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='0' AND B(21)='0' AND B(10)='0' )then
          cVar1S14S16P016P015N034N037(0) <='1';
          else
          cVar1S14S16P016P015N034N037(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='1' AND A(26)='0' AND A(10)='0' )then
          cVar1S15S16P016P015P006P019(0) <='1';
          else
          cVar1S15S16P016P015P006P019(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='1' AND A(26)='0' AND A(10)='0' )then
          cVar1S16S16P016P015P006P019(0) <='1';
          else
          cVar1S16S16P016P015P006P019(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='1' AND A(26)='0' AND A(10)='1' )then
          cVar1S17S16P016P015P006P019(0) <='1';
          else
          cVar1S17S16P016P015P006P019(0) <='0';
          end if;
        if(A(21)='1' AND A(12)='1' AND A(26)='1' AND A(14)='0' )then
          cVar1S18S16P016P015P006P011(0) <='1';
          else
          cVar1S18S16P016P015P006P011(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='1' )then
          cVar1S0S17P023P042nsss(0) <='1';
          else
          cVar1S0S17P023P042nsss(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='0' AND A(17)='1' )then
          cVar1S1S17P023N042P005nsss(0) <='1';
          else
          cVar1S1S17P023N042P005nsss(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='0' AND A(17)='0' AND D(16)='0' )then
          cVar1S2S17P023N042N005P067(0) <='1';
          else
          cVar1S2S17P023N042N005P067(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='1' AND A(26)='0' )then
          cVar1S3S17N023P005P053P006(0) <='1';
          else
          cVar1S3S17N023P005P053P006(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='1' AND A(26)='0' )then
          cVar1S4S17N023P005P053P006(0) <='1';
          else
          cVar1S4S17N023P005P053P006(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='1' AND A(26)='1' )then
          cVar1S5S17N023P005P053P006(0) <='1';
          else
          cVar1S5S17N023P005P053P006(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='1' )then
          cVar1S6S17N023P005N053P058(0) <='1';
          else
          cVar1S6S17N023P005N053P058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='1' )then
          cVar1S7S17N023P005N053P058(0) <='1';
          else
          cVar1S7S17N023P005N053P058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='1' )then
          cVar1S8S17N023P005N053P058(0) <='1';
          else
          cVar1S8S17N023P005N053P058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='0' )then
          cVar1S9S17N023P005N053N058(0) <='1';
          else
          cVar1S9S17N023P005N053N058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='0' )then
          cVar1S10S17N023P005N053N058(0) <='1';
          else
          cVar1S10S17N023P005N053N058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='0' )then
          cVar1S11S17N023P005N053N058(0) <='1';
          else
          cVar1S11S17N023P005N053N058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='0' AND E(20)='0' AND D(10)='0' )then
          cVar1S12S17N023P005N053N058(0) <='1';
          else
          cVar1S12S17N023P005N053N058(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='1' AND A(26)='0' AND E(23)='1' )then
          cVar1S13S17N023P005P006P041nsss(0) <='1';
          else
          cVar1S13S17N023P005P006P041nsss(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='1' AND A(26)='0' AND E(23)='0' )then
          cVar1S14S17N023P005P006N041(0) <='1';
          else
          cVar1S14S17N023P005P006N041(0) <='0';
          end if;
        if(B(17)='0' AND A(17)='1' AND A(26)='0' AND E(23)='0' )then
          cVar1S15S17N023P005P006N041(0) <='1';
          else
          cVar1S15S17N023P005P006N041(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='1' AND D(23)='0' AND B(26)='0' )then
          cVar1S0S18P011P058P039P024(0) <='1';
          else
          cVar1S0S18P011P058P039P024(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='1' AND D(23)='0' AND B(26)='0' )then
          cVar1S1S18P011P058P039P024(0) <='1';
          else
          cVar1S1S18P011P058P039P024(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='1' AND D(23)='0' AND B(26)='0' )then
          cVar1S2S18P011P058P039P024(0) <='1';
          else
          cVar1S2S18P011P058P039P024(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='1' AND D(23)='0' AND B(26)='1' )then
          cVar1S3S18P011P058P039P024(0) <='1';
          else
          cVar1S3S18P011P058P039P024(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='1' AND B(16)='1' )then
          cVar1S4S18P011N058P046P025nsss(0) <='1';
          else
          cVar1S4S18P011N058P046P025nsss(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S5S18P011N058P046N025(0) <='1';
          else
          cVar1S5S18P011N058P046N025(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='1' AND B(16)='0' )then
          cVar1S6S18P011N058P046N025(0) <='1';
          else
          cVar1S6S18P011N058P046N025(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='0' AND B(18)='1' )then
          cVar1S7S18P011N058N046P021(0) <='1';
          else
          cVar1S7S18P011N058N046P021(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='0' AND B(18)='1' )then
          cVar1S8S18P011N058N046P021(0) <='1';
          else
          cVar1S8S18P011N058N046P021(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='0' AND B(18)='0' )then
          cVar1S9S18P011N058N046N021(0) <='1';
          else
          cVar1S9S18P011N058N046N021(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='0' AND B(18)='0' )then
          cVar1S10S18P011N058N046N021(0) <='1';
          else
          cVar1S10S18P011N058N046N021(0) <='0';
          end if;
        if(A(14)='0' AND D(10)='0' AND D(13)='0' AND B(18)='0' )then
          cVar1S11S18P011N058N046N021(0) <='1';
          else
          cVar1S11S18P011N058N046N021(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='1' AND D( 8)='0' AND D(11)='1' )then
          cVar1S12S18P011P029P066P054nsss(0) <='1';
          else
          cVar1S12S18P011P029P066P054nsss(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='1' AND D( 8)='0' AND D(11)='0' )then
          cVar1S13S18P011P029P066N054(0) <='1';
          else
          cVar1S13S18P011P029P066N054(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='1' AND D( 8)='0' AND D(11)='0' )then
          cVar1S14S18P011P029P066N054(0) <='1';
          else
          cVar1S14S18P011P029P066N054(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='1' AND D( 8)='0' AND D(11)='0' )then
          cVar1S15S18P011P029P066N054(0) <='1';
          else
          cVar1S15S18P011P029P066N054(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='0' AND A(13)='0' AND B(22)='0' )then
          cVar1S16S18P011N029P013P032(0) <='1';
          else
          cVar1S16S18P011N029P013P032(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='0' AND A(13)='0' AND B(22)='0' )then
          cVar1S17S18P011N029P013P032(0) <='1';
          else
          cVar1S17S18P011N029P013P032(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='0' AND A(13)='0' AND B(22)='0' )then
          cVar1S18S18P011N029P013P032(0) <='1';
          else
          cVar1S18S18P011N029P013P032(0) <='0';
          end if;
        if(A(14)='1' AND B(14)='0' AND A(13)='0' AND B(22)='1' )then
          cVar1S19S18P011N029P013P032(0) <='1';
          else
          cVar1S19S18P011N029P013P032(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' )then
          cVar1S0S19P021P040nsss(0) <='1';
          else
          cVar1S0S19P021P040nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(23)='1' )then
          cVar1S1S19P021N040P041nsss(0) <='1';
          else
          cVar1S1S19P021N040P041nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(23)='0' AND E(11)='0' )then
          cVar1S2S19P021N040N041P056(0) <='1';
          else
          cVar1S2S19P021N040N041P056(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(23)='0' AND E(11)='0' )then
          cVar1S3S19P021N040N041P056(0) <='1';
          else
          cVar1S3S19P021N040N041P056(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='1' AND D(23)='0' )then
          cVar1S4S19N021P001P058P039(0) <='1';
          else
          cVar1S4S19N021P001P058P039(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='1' AND D(23)='0' )then
          cVar1S5S19N021P001P058P039(0) <='1';
          else
          cVar1S5S19N021P001P058P039(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='0' AND B(28)='1' )then
          cVar1S6S19N021P001N058P020(0) <='1';
          else
          cVar1S6S19N021P001N058P020(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='0' AND B(28)='1' )then
          cVar1S7S19N021P001N058P020(0) <='1';
          else
          cVar1S7S19N021P001N058P020(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='0' AND B(28)='1' )then
          cVar1S8S19N021P001N058P020(0) <='1';
          else
          cVar1S8S19N021P001N058P020(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='0' AND D(10)='0' AND B(28)='0' )then
          cVar1S9S19N021P001N058N020(0) <='1';
          else
          cVar1S9S19N021P001N058N020(0) <='0';
          end if;
        if(B(18)='0' AND A(19)='1' AND D(20)='0' AND A(27)='0' )then
          cVar1S10S19N021P001P051P004(0) <='1';
          else
          cVar1S10S19N021P001P051P004(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='1' AND D(14)='1' )then
          cVar1S0S20P032P023P042nsss(0) <='1';
          else
          cVar1S0S20P032P023P042nsss(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='1' AND D(14)='0' AND A(17)='1' )then
          cVar1S1S20P032P023N042P005nsss(0) <='1';
          else
          cVar1S1S20P032P023N042P005nsss(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='1' AND D(14)='0' AND A(17)='0' )then
          cVar1S2S20P032P023N042N005(0) <='1';
          else
          cVar1S2S20P032P023N042N005(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='0' AND E(11)='1' )then
          cVar1S3S20P032N023P005P056(0) <='1';
          else
          cVar1S3S20P032N023P005P056(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='0' AND E(11)='0' )then
          cVar1S4S20P032N023P005N056(0) <='1';
          else
          cVar1S4S20P032N023P005N056(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='0' AND E(11)='0' )then
          cVar1S5S20P032N023P005N056(0) <='1';
          else
          cVar1S5S20P032N023P005N056(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='0' AND E(11)='0' )then
          cVar1S6S20P032N023P005N056(0) <='1';
          else
          cVar1S6S20P032N023P005N056(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='1' AND B(13)='0' )then
          cVar1S7S20P032N023P005P031(0) <='1';
          else
          cVar1S7S20P032N023P005P031(0) <='0';
          end if;
        if(B(22)='0' AND B(17)='0' AND A(17)='1' AND B(13)='0' )then
          cVar1S8S20P032N023P005P031(0) <='1';
          else
          cVar1S8S20P032N023P005P031(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='1' AND D(20)='0' )then
          cVar1S9S20P032P008P014P051(0) <='1';
          else
          cVar1S9S20P032P008P014P051(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='1' AND D(20)='0' )then
          cVar1S10S20P032P008P014P051(0) <='1';
          else
          cVar1S10S20P032P008P014P051(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='0' AND A(23)='1' )then
          cVar1S11S20P032P008N014P012(0) <='1';
          else
          cVar1S11S20P032P008N014P012(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='0' AND A(23)='1' )then
          cVar1S12S20P032P008N014P012(0) <='1';
          else
          cVar1S12S20P032P008N014P012(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='0' AND A(23)='0' )then
          cVar1S13S20P032P008N014N012(0) <='1';
          else
          cVar1S13S20P032P008N014N012(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='0' AND A(22)='0' AND A(23)='0' )then
          cVar1S14S20P032P008N014N012(0) <='1';
          else
          cVar1S14S20P032P008N014N012(0) <='0';
          end if;
        if(B(22)='1' AND A(25)='1' AND A(26)='0' AND E( 8)='1' )then
          cVar1S15S20P032P008P006P068(0) <='1';
          else
          cVar1S15S20P032P008P006P068(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='1' )then
          cVar1S0S21P023P042nsss(0) <='1';
          else
          cVar1S0S21P023P042nsss(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='0' AND B(26)='0' AND A(17)='1' )then
          cVar1S1S21P023N042P024P005nsss(0) <='1';
          else
          cVar1S1S21P023N042P024P005nsss(0) <='0';
          end if;
        if(B(17)='1' AND D(14)='0' AND B(26)='0' AND A(17)='0' )then
          cVar1S2S21P023N042P024N005(0) <='1';
          else
          cVar1S2S21P023N042P024N005(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='1' AND B(26)='1' )then
          cVar1S3S21N023P001P047P024(0) <='1';
          else
          cVar1S3S21N023P001P047P024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='1' AND B(26)='0' )then
          cVar1S4S21N023P001P047N024(0) <='1';
          else
          cVar1S4S21N023P001P047N024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='1' AND B(26)='0' )then
          cVar1S5S21N023P001P047N024(0) <='1';
          else
          cVar1S5S21N023P001P047N024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='1' AND B(26)='0' )then
          cVar1S6S21N023P001P047N024(0) <='1';
          else
          cVar1S6S21N023P001P047N024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='0' AND B(26)='0' )then
          cVar1S7S21N023P001N047P024(0) <='1';
          else
          cVar1S7S21N023P001N047P024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='0' AND B(26)='0' )then
          cVar1S8S21N023P001N047P024(0) <='1';
          else
          cVar1S8S21N023P001N047P024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='0' AND D(21)='0' AND B(26)='1' )then
          cVar1S9S21N023P001N047P024(0) <='1';
          else
          cVar1S9S21N023P001N047P024(0) <='0';
          end if;
        if(B(17)='0' AND A(19)='1' AND A(26)='0' AND B(24)='0' )then
          cVar1S10S21N023P001P006P028(0) <='1';
          else
          cVar1S10S21N023P001P006P028(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='0' AND B(15)='1' )then
          cVar1S0S22P001P010P028P027(0) <='1';
          else
          cVar1S0S22P001P010P028P027(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='0' AND B(15)='1' )then
          cVar1S1S22P001P010P028P027(0) <='1';
          else
          cVar1S1S22P001P010P028P027(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='0' AND B(15)='0' )then
          cVar1S2S22P001P010P028N027(0) <='1';
          else
          cVar1S2S22P001P010P028N027(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='0' AND B(15)='0' )then
          cVar1S3S22P001P010P028N027(0) <='1';
          else
          cVar1S3S22P001P010P028N027(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='0' AND B(15)='0' )then
          cVar1S4S22P001P010P028N027(0) <='1';
          else
          cVar1S4S22P001P010P028N027(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='1' AND A(29)='0' )then
          cVar1S5S22P001P010P028P000(0) <='1';
          else
          cVar1S5S22P001P010P028P000(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='0' AND B(24)='1' AND A(29)='0' )then
          cVar1S6S22P001P010P028P000(0) <='1';
          else
          cVar1S6S22P001P010P028P000(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='1' AND B(24)='1' AND B(21)='0' )then
          cVar1S7S22P001P010P028P034nsss(0) <='1';
          else
          cVar1S7S22P001P010P028P034nsss(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='1' AND B(24)='0' AND E(22)='0' )then
          cVar1S8S22P001P010N028P045(0) <='1';
          else
          cVar1S8S22P001P010N028P045(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='1' AND B(24)='0' AND E(22)='0' )then
          cVar1S9S22P001P010N028P045(0) <='1';
          else
          cVar1S9S22P001P010N028P045(0) <='0';
          end if;
        if(A(19)='0' AND A(24)='1' AND B(24)='0' AND E(22)='1' )then
          cVar1S10S22P001P010N028P045(0) <='1';
          else
          cVar1S10S22P001P010N028P045(0) <='0';
          end if;
        if(A(19)='1' AND A(27)='0' AND D(20)='0' AND B(26)='0' )then
          cVar1S11S22P001P004P051P024(0) <='1';
          else
          cVar1S11S22P001P004P051P024(0) <='0';
          end if;
        if(A(19)='1' AND A(27)='0' AND D(20)='0' AND B(26)='0' )then
          cVar1S12S22P001P004P051P024(0) <='1';
          else
          cVar1S12S22P001P004P051P024(0) <='0';
          end if;
        if(B(15)='1' AND A(29)='0' AND E(13)='1' )then
          cVar1S0S23P027P000P048nsss(0) <='1';
          else
          cVar1S0S23P027P000P048nsss(0) <='0';
          end if;
        if(B(15)='1' AND A(29)='0' AND E(13)='0' AND B(11)='0' )then
          cVar1S1S23P027P000N048P035(0) <='1';
          else
          cVar1S1S23P027P000N048P035(0) <='0';
          end if;
        if(B(15)='1' AND A(29)='0' AND E(13)='0' AND B(11)='0' )then
          cVar1S2S23P027P000N048P035(0) <='1';
          else
          cVar1S2S23P027P000N048P035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='1' AND D(14)='1' )then
          cVar1S3S23N027P009P023P042nsss(0) <='1';
          else
          cVar1S3S23N027P009P023P042nsss(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='1' AND D(14)='0' )then
          cVar1S4S23N027P009P023N042(0) <='1';
          else
          cVar1S4S23N027P009P023N042(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='1' AND D(14)='0' )then
          cVar1S5S23N027P009P023N042(0) <='1';
          else
          cVar1S5S23N027P009P023N042(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='0' AND B(11)='1' )then
          cVar1S6S23N027P009N023P035(0) <='1';
          else
          cVar1S6S23N027P009N023P035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='0' AND B(11)='1' )then
          cVar1S7S23N027P009N023P035(0) <='1';
          else
          cVar1S7S23N027P009N023P035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='0' AND B(11)='0' )then
          cVar1S8S23N027P009N023N035(0) <='1';
          else
          cVar1S8S23N027P009N023N035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='0' AND B(11)='0' )then
          cVar1S9S23N027P009N023N035(0) <='1';
          else
          cVar1S9S23N027P009N023N035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='0' AND B(17)='0' AND B(11)='0' )then
          cVar1S10S23N027P009N023N035(0) <='1';
          else
          cVar1S10S23N027P009N023N035(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='1' AND E( 8)='0' AND D( 9)='0' )then
          cVar1S11S23N027P009P068P062(0) <='1';
          else
          cVar1S11S23N027P009P068P062(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='1' AND E( 8)='0' AND D( 9)='0' )then
          cVar1S12S23N027P009P068P062(0) <='1';
          else
          cVar1S12S23N027P009P068P062(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='1' AND E( 8)='0' AND D( 9)='1' )then
          cVar1S13S23N027P009P068P062(0) <='1';
          else
          cVar1S13S23N027P009P068P062(0) <='0';
          end if;
        if(B(15)='0' AND A(15)='1' AND E( 8)='1' AND A(28)='0' )then
          cVar1S14S23N027P009P068P002(0) <='1';
          else
          cVar1S14S23N027P009P068P002(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S0S24P008P026P055P057(0) <='1';
          else
          cVar1S0S24P008P026P055P057(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S1S24P008P026P055P057(0) <='1';
          else
          cVar1S1S24P008P026P055P057(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S2S24P008P026P055P057(0) <='1';
          else
          cVar1S2S24P008P026P055P057(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='1' AND E(19)='0' )then
          cVar1S3S24P008P026P055N057(0) <='1';
          else
          cVar1S3S24P008P026P055N057(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='1' AND E(19)='0' )then
          cVar1S4S24P008P026P055N057(0) <='1';
          else
          cVar1S4S24P008P026P055N057(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='0' AND E(23)='1' )then
          cVar1S5S24P008P026N055P041(0) <='1';
          else
          cVar1S5S24P008P026N055P041(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='0' AND E(23)='1' )then
          cVar1S6S24P008P026N055P041(0) <='1';
          else
          cVar1S6S24P008P026N055P041(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='0' AND E(23)='1' )then
          cVar1S7S24P008P026N055P041(0) <='1';
          else
          cVar1S7S24P008P026N055P041(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='0' AND D(19)='0' AND E(23)='0' )then
          cVar1S8S24P008P026N055N041(0) <='1';
          else
          cVar1S8S24P008P026N055N041(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='1' AND E(22)='0' AND D(21)='1' )then
          cVar1S9S24P008P026P045P047nsss(0) <='1';
          else
          cVar1S9S24P008P026P045P047nsss(0) <='0';
          end if;
        if(A(25)='0' AND B(25)='1' AND E(22)='0' AND D(21)='0' )then
          cVar1S10S24P008P026P045N047(0) <='1';
          else
          cVar1S10S24P008P026P045N047(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='1' AND A(27)='0' AND D(20)='1' )then
          cVar1S11S24P008P026P004P051nsss(0) <='1';
          else
          cVar1S11S24P008P026P004P051nsss(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='1' AND A(27)='0' AND D(20)='0' )then
          cVar1S12S24P008P026P004N051(0) <='1';
          else
          cVar1S12S24P008P026P004N051(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='1' AND A(27)='0' AND D(20)='0' )then
          cVar1S13S24P008P026P004N051(0) <='1';
          else
          cVar1S13S24P008P026P004N051(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='0' AND B(22)='0' AND D(23)='0' )then
          cVar1S14S24P008N026P032P039(0) <='1';
          else
          cVar1S14S24P008N026P032P039(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='0' AND B(22)='0' AND D(23)='0' )then
          cVar1S15S24P008N026P032P039(0) <='1';
          else
          cVar1S15S24P008N026P032P039(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='0' AND B(22)='0' AND D(23)='0' )then
          cVar1S16S24P008N026P032P039(0) <='1';
          else
          cVar1S16S24P008N026P032P039(0) <='0';
          end if;
        if(A(25)='1' AND B(25)='0' AND B(22)='0' AND D(23)='0' )then
          cVar1S17S24P008N026P032P039(0) <='1';
          else
          cVar1S17S24P008N026P032P039(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND B(23)='1' AND E(19)='1' )then
          cVar1S0S25P055P026P030P057(0) <='1';
          else
          cVar1S0S25P055P026P030P057(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND B(23)='1' AND E(19)='1' )then
          cVar1S1S25P055P026P030P057(0) <='1';
          else
          cVar1S1S25P055P026P030P057(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND B(23)='0' AND B(13)='1' )then
          cVar1S2S25P055P026N030P031(0) <='1';
          else
          cVar1S2S25P055P026N030P031(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND B(23)='0' AND B(13)='0' )then
          cVar1S3S25P055P026N030N031(0) <='1';
          else
          cVar1S3S25P055P026N030N031(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND B(23)='0' AND B(13)='0' )then
          cVar1S4S25P055P026N030N031(0) <='1';
          else
          cVar1S4S25P055P026N030N031(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='1' AND B(28)='1' )then
          cVar1S5S25N055P057P041P020nsss(0) <='1';
          else
          cVar1S5S25N055P057P041P020nsss(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='1' AND B(28)='0' )then
          cVar1S6S25N055P057P041N020(0) <='1';
          else
          cVar1S6S25N055P057P041N020(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='1' AND B(28)='0' )then
          cVar1S7S25N055P057P041N020(0) <='1';
          else
          cVar1S7S25N055P057P041N020(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='0' AND E(20)='1' )then
          cVar1S8S25N055P057N041P053(0) <='1';
          else
          cVar1S8S25N055P057N041P053(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='0' AND E(20)='1' )then
          cVar1S9S25N055P057N041P053(0) <='1';
          else
          cVar1S9S25N055P057N041P053(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='0' AND E(20)='1' )then
          cVar1S10S25N055P057N041P053(0) <='1';
          else
          cVar1S10S25N055P057N041P053(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='0' AND E(20)='0' )then
          cVar1S11S25N055P057N041N053(0) <='1';
          else
          cVar1S11S25N055P057N041N053(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='0' AND E(23)='0' AND E(20)='0' )then
          cVar1S12S25N055P057N041N053(0) <='1';
          else
          cVar1S12S25N055P057N041N053(0) <='0';
          end if;
        if(D(19)='0' AND E(19)='1' AND E(20)='0' AND B(10)='0' )then
          cVar1S13S25N055P057P053P037(0) <='1';
          else
          cVar1S13S25N055P057P053P037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='1' AND A(28)='0' )then
          cVar1S0S26P017P019P037P002(0) <='1';
          else
          cVar1S0S26P017P019P037P002(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='1' AND A(28)='0' )then
          cVar1S1S26P017P019P037P002(0) <='1';
          else
          cVar1S1S26P017P019P037P002(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='1' AND A(28)='0' )then
          cVar1S2S26P017P019P037P002(0) <='1';
          else
          cVar1S2S26P017P019P037P002(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='1' AND A(28)='0' )then
          cVar1S3S26P017P019P037P002(0) <='1';
          else
          cVar1S3S26P017P019P037P002(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='1' AND A(28)='1' )then
          cVar1S4S26P017P019P037P002(0) <='1';
          else
          cVar1S4S26P017P019P037P002(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='0' AND A(20)='0' )then
          cVar1S5S26P017P019N037P018(0) <='1';
          else
          cVar1S5S26P017P019N037P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='0' AND A(20)='0' )then
          cVar1S6S26P017P019N037P018(0) <='1';
          else
          cVar1S6S26P017P019N037P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='0' AND A(20)='0' )then
          cVar1S7S26P017P019N037P018(0) <='1';
          else
          cVar1S7S26P017P019N037P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='0' AND A(20)='1' )then
          cVar1S8S26P017P019N037P018(0) <='1';
          else
          cVar1S8S26P017P019N037P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND B(10)='0' AND A(20)='1' )then
          cVar1S9S26P017P019N037P018(0) <='1';
          else
          cVar1S9S26P017P019N037P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='0' AND E( 9)='0' )then
          cVar1S10S26P017N019P037P064nsss(0) <='1';
          else
          cVar1S10S26P017N019P037P064nsss(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='0' AND E( 9)='1' )then
          cVar1S11S26P017N019P037P064(0) <='1';
          else
          cVar1S11S26P017N019P037P064(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='0' AND E( 9)='1' )then
          cVar1S12S26P017N019P037P064(0) <='1';
          else
          cVar1S12S26P017N019P037P064(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='0' AND E( 9)='1' )then
          cVar1S13S26P017N019P037P064(0) <='1';
          else
          cVar1S13S26P017N019P037P064(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='1' AND A(18)='0' )then
          cVar1S14S26P017N019P037P003(0) <='1';
          else
          cVar1S14S26P017N019P037P003(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='1' AND A(18)='0' )then
          cVar1S15S26P017N019P037P003(0) <='1';
          else
          cVar1S15S26P017N019P037P003(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND B(10)='1' AND A(18)='0' )then
          cVar1S16S26P017N019P037P003(0) <='1';
          else
          cVar1S16S26P017N019P037P003(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='0' AND E( 9)='1' )then
          cVar1S17S26P017P037P019P064(0) <='1';
          else
          cVar1S17S26P017P037P019P064(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='0' AND E( 9)='1' )then
          cVar1S18S26P017P037P019P064(0) <='1';
          else
          cVar1S18S26P017P037P019P064(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='0' AND E( 9)='0' )then
          cVar1S19S26P017P037P019N064(0) <='1';
          else
          cVar1S19S26P017P037P019N064(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='1' AND A(13)='0' )then
          cVar1S20S26P017P037P019P013(0) <='1';
          else
          cVar1S20S26P017P037P019P013(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='1' AND A(13)='0' )then
          cVar1S21S26P017P037P019P013(0) <='1';
          else
          cVar1S21S26P017P037P019P013(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='1' AND A(13)='0' )then
          cVar1S22S26P017P037P019P013(0) <='1';
          else
          cVar1S22S26P017P037P019P013(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='1' AND A(13)='1' )then
          cVar1S23S26P017P037P019P013(0) <='1';
          else
          cVar1S23S26P017P037P019P013(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='1' AND A(10)='1' AND A(13)='1' )then
          cVar1S24S26P017P037P019P013(0) <='1';
          else
          cVar1S24S26P017P037P019P013(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='1' AND A(10)='0' )then
          cVar1S25S26P017N037P035P019(0) <='1';
          else
          cVar1S25S26P017N037P035P019(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='1' AND A(10)='0' )then
          cVar1S26S26P017N037P035P019(0) <='1';
          else
          cVar1S26S26P017N037P035P019(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='1' AND A(10)='0' )then
          cVar1S27S26P017N037P035P019(0) <='1';
          else
          cVar1S27S26P017N037P035P019(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='1' AND A(10)='1' )then
          cVar1S28S26P017N037P035P019(0) <='1';
          else
          cVar1S28S26P017N037P035P019(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='0' AND E( 9)='0' )then
          cVar1S29S26P017N037N035P064(0) <='1';
          else
          cVar1S29S26P017N037N035P064(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='0' AND E( 9)='1' )then
          cVar1S30S26P017N037N035P064(0) <='1';
          else
          cVar1S30S26P017N037N035P064(0) <='0';
          end if;
        if(A(11)='1' AND B(10)='0' AND B(11)='0' AND E( 9)='1' )then
          cVar1S31S26P017N037N035P064(0) <='1';
          else
          cVar1S31S26P017N037N035P064(0) <='0';
          end if;
        if(A(11)='1' AND D(20)='0' AND E(13)='0' AND B(16)='0' )then
          cVar1S0S27P017P051P048P025(0) <='1';
          else
          cVar1S0S27P017P051P048P025(0) <='0';
          end if;
        if(A(11)='1' AND D(20)='0' AND E(13)='1' AND B(25)='1' )then
          cVar1S1S27P017P051P048P026nsss(0) <='1';
          else
          cVar1S1S27P017P051P048P026nsss(0) <='0';
          end if;
        if(A(11)='1' AND D(20)='1' AND D(10)='0' AND E(23)='0' )then
          cVar1S2S27P017P051P058P041(0) <='1';
          else
          cVar1S2S27P017P051P058P041(0) <='0';
          end if;
        if(A(11)='1' AND D(20)='1' AND D(10)='0' AND E(23)='0' )then
          cVar1S3S27P017P051P058P041(0) <='1';
          else
          cVar1S3S27P017P051P058P041(0) <='0';
          end if;
        if(A(11)='1' AND D(20)='1' AND D(10)='0' AND E(23)='0' )then
          cVar1S4S27P017P051P058P041(0) <='1';
          else
          cVar1S4S27P017P051P058P041(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='1' AND B(26)='0' )then
          cVar1S5S27N017P019P067P024(0) <='1';
          else
          cVar1S5S27N017P019P067P024(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='1' AND B(26)='0' )then
          cVar1S6S27N017P019P067P024(0) <='1';
          else
          cVar1S6S27N017P019P067P024(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='0' AND B(10)='1' )then
          cVar1S7S27N017P019N067P037(0) <='1';
          else
          cVar1S7S27N017P019N067P037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='0' AND B(10)='1' )then
          cVar1S8S27N017P019N067P037(0) <='1';
          else
          cVar1S8S27N017P019N067P037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='0' AND B(10)='1' )then
          cVar1S9S27N017P019N067P037(0) <='1';
          else
          cVar1S9S27N017P019N067P037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='0' AND B(10)='1' )then
          cVar1S10S27N017P019N067P037(0) <='1';
          else
          cVar1S10S27N017P019N067P037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='1' AND D(16)='0' AND B(10)='0' )then
          cVar1S11S27N017P019N067N037(0) <='1';
          else
          cVar1S11S27N017P019N067N037(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='1' )then
          cVar1S12S27N017N019P068P027(0) <='1';
          else
          cVar1S12S27N017N019P068P027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='1' )then
          cVar1S13S27N017N019P068P027(0) <='1';
          else
          cVar1S13S27N017N019P068P027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='1' )then
          cVar1S14S27N017N019P068P027(0) <='1';
          else
          cVar1S14S27N017N019P068P027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='0' )then
          cVar1S15S27N017N019P068N027(0) <='1';
          else
          cVar1S15S27N017N019P068N027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='0' )then
          cVar1S16S27N017N019P068N027(0) <='1';
          else
          cVar1S16S27N017N019P068N027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='0' )then
          cVar1S17S27N017N019P068N027(0) <='1';
          else
          cVar1S17S27N017N019P068N027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='0' AND B(15)='0' )then
          cVar1S18S27N017N019P068N027(0) <='1';
          else
          cVar1S18S27N017N019P068N027(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='1' AND A(20)='1' )then
          cVar1S19S27N017N019P068P018(0) <='1';
          else
          cVar1S19S27N017N019P068P018(0) <='0';
          end if;
        if(A(11)='0' AND A(10)='0' AND E( 8)='1' AND A(20)='0' )then
          cVar1S20S27N017N019P068N018(0) <='1';
          else
          cVar1S20S27N017N019P068N018(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='0' AND E(14)='1' )then
          cVar1S0S28P017P068P064P044(0) <='1';
          else
          cVar1S0S28P017P068P064P044(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='0' AND E(14)='1' )then
          cVar1S1S28P017P068P064P044(0) <='1';
          else
          cVar1S1S28P017P068P064P044(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='0' AND E(14)='1' )then
          cVar1S2S28P017P068P064P044(0) <='1';
          else
          cVar1S2S28P017P068P064P044(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='0' AND E(14)='0' )then
          cVar1S3S28P017P068P064N044(0) <='1';
          else
          cVar1S3S28P017P068P064N044(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='0' AND E(14)='0' )then
          cVar1S4S28P017P068P064N044(0) <='1';
          else
          cVar1S4S28P017P068P064N044(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='1' AND D(19)='1' )then
          cVar1S5S28P017P068P064P055nsss(0) <='1';
          else
          cVar1S5S28P017P068P064P055nsss(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='1' AND D(19)='0' )then
          cVar1S6S28P017P068P064N055(0) <='1';
          else
          cVar1S6S28P017P068P064N055(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='0' AND E( 9)='1' AND D(19)='0' )then
          cVar1S7S28P017P068P064N055(0) <='1';
          else
          cVar1S7S28P017P068P064N055(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='1' AND E( 9)='1' )then
          cVar1S8S28P017P068P019P064(0) <='1';
          else
          cVar1S8S28P017P068P019P064(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='1' AND E( 9)='1' )then
          cVar1S9S28P017P068P019P064(0) <='1';
          else
          cVar1S9S28P017P068P019P064(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='1' AND E( 9)='0' )then
          cVar1S10S28P017P068P019N064(0) <='1';
          else
          cVar1S10S28P017P068P019N064(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='0' AND D(16)='0' )then
          cVar1S11S28P017P068N019P067(0) <='1';
          else
          cVar1S11S28P017P068N019P067(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='0' AND D(16)='0' )then
          cVar1S12S28P017P068N019P067(0) <='1';
          else
          cVar1S12S28P017P068N019P067(0) <='0';
          end if;
        if(A(11)='0' AND E( 8)='1' AND A(10)='0' AND D(16)='0' )then
          cVar1S13S28P017P068N019P067(0) <='1';
          else
          cVar1S13S28P017P068N019P067(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='1' AND D(16)='0' )then
          cVar1S14S28P017P019P016P067(0) <='1';
          else
          cVar1S14S28P017P019P016P067(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='1' AND D(16)='0' )then
          cVar1S15S28P017P019P016P067(0) <='1';
          else
          cVar1S15S28P017P019P016P067(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='1' AND D(16)='1' )then
          cVar1S16S28P017P019P016P067(0) <='1';
          else
          cVar1S16S28P017P019P016P067(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='1' AND D(16)='1' )then
          cVar1S17S28P017P019P016P067(0) <='1';
          else
          cVar1S17S28P017P019P016P067(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='0' AND A(24)='1' )then
          cVar1S18S28P017P019N016P010(0) <='1';
          else
          cVar1S18S28P017P019N016P010(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='0' AND A(24)='0' )then
          cVar1S19S28P017P019N016N010(0) <='1';
          else
          cVar1S19S28P017P019N016N010(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='0' AND A(24)='0' )then
          cVar1S20S28P017P019N016N010(0) <='1';
          else
          cVar1S20S28P017P019N016N010(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='0' AND A(21)='0' AND A(24)='0' )then
          cVar1S21S28P017P019N016N010(0) <='1';
          else
          cVar1S21S28P017P019N016N010(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='0' AND E(19)='0' )then
          cVar1S22S28P017P019P064P057(0) <='1';
          else
          cVar1S22S28P017P019P064P057(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='0' AND E(19)='1' )then
          cVar1S23S28P017P019P064P057(0) <='1';
          else
          cVar1S23S28P017P019P064P057(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='1' AND E( 8)='1' )then
          cVar1S24S28P017P019P064P068(0) <='1';
          else
          cVar1S24S28P017P019P064P068(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='1' AND E( 8)='1' )then
          cVar1S25S28P017P019P064P068(0) <='1';
          else
          cVar1S25S28P017P019P064P068(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='1' AND E( 8)='0' )then
          cVar1S26S28P017P019P064N068(0) <='1';
          else
          cVar1S26S28P017P019P064N068(0) <='0';
          end if;
        if(A(11)='1' AND A(10)='1' AND E( 9)='1' AND E( 8)='0' )then
          cVar1S27S28P017P019P064N068(0) <='1';
          else
          cVar1S27S28P017P019P064N068(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='1' AND B(22)='0' )then
          cVar1S0S29P017P013P011P032(0) <='1';
          else
          cVar1S0S29P017P013P011P032(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='1' AND B(22)='0' )then
          cVar1S1S29P017P013P011P032(0) <='1';
          else
          cVar1S1S29P017P013P011P032(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='0' AND B(14)='0' )then
          cVar1S2S29P017P013N011P029(0) <='1';
          else
          cVar1S2S29P017P013N011P029(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='0' AND B(14)='0' )then
          cVar1S3S29P017P013N011P029(0) <='1';
          else
          cVar1S3S29P017P013N011P029(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='0' AND B(14)='0' )then
          cVar1S4S29P017P013N011P029(0) <='1';
          else
          cVar1S4S29P017P013N011P029(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='0' AND A(14)='0' AND B(14)='1' )then
          cVar1S5S29P017P013N011P029(0) <='1';
          else
          cVar1S5S29P017P013N011P029(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='1' AND D(16)='0' AND B(15)='0' )then
          cVar1S6S29P017P013P067P027(0) <='1';
          else
          cVar1S6S29P017P013P067P027(0) <='0';
          end if;
        if(A(11)='1' AND A(13)='1' AND D(16)='1' AND D(20)='0' )then
          cVar1S7S29P017P013P067P051(0) <='1';
          else
          cVar1S7S29P017P013P067P051(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='1' AND B(17)='1' )then
          cVar1S8S29N017P044P023nsss(0) <='1';
          else
          cVar1S8S29N017P044P023nsss(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S9S29N017P044N023P025nsss(0) <='1';
          else
          cVar1S9S29N017P044N023P025nsss(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S10S29N017P044N023N025(0) <='1';
          else
          cVar1S10S29N017P044N023N025(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S11S29N017N044P055P057(0) <='1';
          else
          cVar1S11S29N017N044P055P057(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S12S29N017N044P055P057(0) <='1';
          else
          cVar1S12S29N017N044P055P057(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S13S29N017N044P055P057(0) <='1';
          else
          cVar1S13S29N017N044P055P057(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='1' AND E(19)='1' )then
          cVar1S14S29N017N044P055P057(0) <='1';
          else
          cVar1S14S29N017N044P055P057(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='1' AND E(19)='0' )then
          cVar1S15S29N017N044P055N057(0) <='1';
          else
          cVar1S15S29N017N044P055N057(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='0' AND E(23)='1' )then
          cVar1S16S29N017N044N055P041(0) <='1';
          else
          cVar1S16S29N017N044N055P041(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='0' AND E(23)='1' )then
          cVar1S17S29N017N044N055P041(0) <='1';
          else
          cVar1S17S29N017N044N055P041(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='0' AND E(23)='0' )then
          cVar1S18S29N017N044N055N041(0) <='1';
          else
          cVar1S18S29N017N044N055N041(0) <='0';
          end if;
        if(A(11)='0' AND E(14)='0' AND D(19)='0' AND E(23)='0' )then
          cVar1S19S29N017N044N055N041(0) <='1';
          else
          cVar1S19S29N017N044N055N041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='1' AND B(22)='0' )then
          cVar1S0S30P017P036P044P032(0) <='1';
          else
          cVar1S0S30P017P036P044P032(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='1' AND B(22)='0' )then
          cVar1S1S30P017P036P044P032(0) <='1';
          else
          cVar1S1S30P017P036P044P032(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='1' AND B(22)='0' )then
          cVar1S2S30P017P036P044P032(0) <='1';
          else
          cVar1S2S30P017P036P044P032(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='0' AND E(23)='1' )then
          cVar1S3S30P017P036N044P041(0) <='1';
          else
          cVar1S3S30P017P036N044P041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='0' AND E(23)='1' )then
          cVar1S4S30P017P036N044P041(0) <='1';
          else
          cVar1S4S30P017P036N044P041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='0' AND E(23)='0' )then
          cVar1S5S30P017P036N044N041(0) <='1';
          else
          cVar1S5S30P017P036N044N041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='0' AND E(23)='0' )then
          cVar1S6S30P017P036N044N041(0) <='1';
          else
          cVar1S6S30P017P036N044N041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='0' AND E(14)='0' AND E(23)='0' )then
          cVar1S7S30P017P036N044N041(0) <='1';
          else
          cVar1S7S30P017P036N044N041(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='1' AND A(27)='0' AND A(13)='1' )then
          cVar1S8S30P017P036P004P013(0) <='1';
          else
          cVar1S8S30P017P036P004P013(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='1' AND A(27)='0' AND A(13)='1' )then
          cVar1S9S30P017P036P004P013(0) <='1';
          else
          cVar1S9S30P017P036P004P013(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='1' AND A(27)='0' AND A(13)='0' )then
          cVar1S10S30P017P036P004N013(0) <='1';
          else
          cVar1S10S30P017P036P004N013(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='1' AND A(27)='0' AND A(13)='0' )then
          cVar1S11S30P017P036P004N013(0) <='1';
          else
          cVar1S11S30P017P036P004N013(0) <='0';
          end if;
        if(A(11)='0' AND B(20)='1' AND A(27)='1' AND A(26)='0' )then
          cVar1S12S30P017P036P004P006(0) <='1';
          else
          cVar1S12S30P017P036P004P006(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='1' AND D(22)='0' )then
          cVar1S13S30P017P044P063P043(0) <='1';
          else
          cVar1S13S30P017P044P063P043(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='1' AND D(22)='0' )then
          cVar1S14S30P017P044P063P043(0) <='1';
          else
          cVar1S14S30P017P044P063P043(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='0' AND E(17)='0' )then
          cVar1S15S30P017P044N063P065(0) <='1';
          else
          cVar1S15S30P017P044N063P065(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='0' AND E(17)='0' )then
          cVar1S16S30P017P044N063P065(0) <='1';
          else
          cVar1S16S30P017P044N063P065(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='0' AND E(17)='0' )then
          cVar1S17S30P017P044N063P065(0) <='1';
          else
          cVar1S17S30P017P044N063P065(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='0' AND D(17)='0' AND E(17)='1' )then
          cVar1S18S30P017P044N063P065(0) <='1';
          else
          cVar1S18S30P017P044N063P065(0) <='0';
          end if;
        if(A(11)='1' AND E(14)='1' AND B(21)='0' AND A(22)='0' )then
          cVar1S19S30P017P044P034P014(0) <='1';
          else
          cVar1S19S30P017P044P034P014(0) <='0';
          end if;
        if(B(12)='1' AND D(11)='0' AND E(18)='1' AND B(22)='0' )then
          cVar1S0S31P033P054P061P032(0) <='1';
          else
          cVar1S0S31P033P054P061P032(0) <='0';
          end if;
        if(B(12)='1' AND D(11)='0' AND E(18)='0' AND D(17)='0' )then
          cVar1S1S31P033P054N061P063(0) <='1';
          else
          cVar1S1S31P033P054N061P063(0) <='0';
          end if;
        if(B(12)='1' AND D(11)='0' AND E(18)='0' AND D(17)='1' )then
          cVar1S2S31P033P054N061P063(0) <='1';
          else
          cVar1S2S31P033P054N061P063(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S3S31N033P061P029P011(0) <='1';
          else
          cVar1S3S31N033P061P029P011(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S4S31N033P061P029N011(0) <='1';
          else
          cVar1S4S31N033P061P029N011(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S5S31N033P061P029N011(0) <='1';
          else
          cVar1S5S31N033P061P029N011(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S6S31N033P061P029N011(0) <='1';
          else
          cVar1S6S31N033P061P029N011(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='0' AND E(15)='1' )then
          cVar1S7S31N033P061N029P040(0) <='1';
          else
          cVar1S7S31N033P061N029P040(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='0' AND E(15)='1' )then
          cVar1S8S31N033P061N029P040(0) <='1';
          else
          cVar1S8S31N033P061N029P040(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='0' AND E(15)='1' )then
          cVar1S9S31N033P061N029P040(0) <='1';
          else
          cVar1S9S31N033P061N029P040(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='0' AND E(15)='0' )then
          cVar1S10S31N033P061N029N040(0) <='1';
          else
          cVar1S10S31N033P061N029N040(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='0' AND B(14)='0' AND E(15)='0' )then
          cVar1S11S31N033P061N029N040(0) <='1';
          else
          cVar1S11S31N033P061N029N040(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='1' AND B(22)='0' )then
          cVar1S12S31N033P061P059P032(0) <='1';
          else
          cVar1S12S31N033P061P059P032(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='1' AND B(22)='0' )then
          cVar1S13S31N033P061P059P032(0) <='1';
          else
          cVar1S13S31N033P061P059P032(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='1' AND B(22)='1' )then
          cVar1S14S31N033P061P059P032(0) <='1';
          else
          cVar1S14S31N033P061P059P032(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='1' AND B(22)='1' )then
          cVar1S15S31N033P061P059P032(0) <='1';
          else
          cVar1S15S31N033P061P059P032(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='0' AND A(20)='1' )then
          cVar1S16S31N033P061N059P018(0) <='1';
          else
          cVar1S16S31N033P061N059P018(0) <='0';
          end if;
        if(B(12)='0' AND E(18)='1' AND D(18)='0' AND A(20)='0' )then
          cVar1S17S31N033P061N059N018(0) <='1';
          else
          cVar1S17S31N033P061N059N018(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='0' AND E( 9)='1' )then
          cVar1S0S32P061P033P060P064(0) <='1';
          else
          cVar1S0S32P061P033P060P064(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='0' AND E( 9)='1' )then
          cVar1S1S32P061P033P060P064(0) <='1';
          else
          cVar1S1S32P061P033P060P064(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='0' AND E( 9)='1' )then
          cVar1S2S32P061P033P060P064(0) <='1';
          else
          cVar1S2S32P061P033P060P064(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='0' AND E( 9)='0' )then
          cVar1S3S32P061P033P060N064(0) <='1';
          else
          cVar1S3S32P061P033P060N064(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='0' AND E( 9)='0' )then
          cVar1S4S32P061P033P060N064(0) <='1';
          else
          cVar1S4S32P061P033P060N064(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='1' AND B(22)='1' )then
          cVar1S5S32P061P033P060P032nsss(0) <='1';
          else
          cVar1S5S32P061P033P060P032nsss(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='1' AND B(22)='0' )then
          cVar1S6S32P061P033P060N032(0) <='1';
          else
          cVar1S6S32P061P033P060N032(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='0' AND E(10)='1' AND B(22)='0' )then
          cVar1S7S32P061P033P060N032(0) <='1';
          else
          cVar1S7S32P061P033P060N032(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='1' AND E(17)='0' AND E(10)='1' )then
          cVar1S8S32P061P033P065P060(0) <='1';
          else
          cVar1S8S32P061P033P065P060(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='1' AND E(17)='0' AND E(10)='1' )then
          cVar1S9S32P061P033P065P060(0) <='1';
          else
          cVar1S9S32P061P033P065P060(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='1' AND E(17)='0' AND E(10)='0' )then
          cVar1S10S32P061P033P065N060(0) <='1';
          else
          cVar1S10S32P061P033P065N060(0) <='0';
          end if;
        if(E(18)='0' AND B(12)='1' AND E(17)='1' AND A(10)='0' )then
          cVar1S11S32P061P033P065P019(0) <='1';
          else
          cVar1S11S32P061P033P065P019(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='0' AND E( 9)='0' )then
          cVar1S12S32P061P059P032P064(0) <='1';
          else
          cVar1S12S32P061P059P032P064(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='0' AND E( 9)='0' )then
          cVar1S13S32P061P059P032P064(0) <='1';
          else
          cVar1S13S32P061P059P032P064(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='0' AND E( 9)='0' )then
          cVar1S14S32P061P059P032P064(0) <='1';
          else
          cVar1S14S32P061P059P032P064(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='0' AND E( 9)='1' )then
          cVar1S15S32P061P059P032P064(0) <='1';
          else
          cVar1S15S32P061P059P032P064(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='1' AND D(16)='1' )then
          cVar1S16S32P061P059P032P067(0) <='1';
          else
          cVar1S16S32P061P059P032P067(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='1' AND D(16)='0' )then
          cVar1S17S32P061P059P032N067(0) <='1';
          else
          cVar1S17S32P061P059P032N067(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='1' AND B(22)='1' AND D(16)='0' )then
          cVar1S18S32P061P059P032N067(0) <='1';
          else
          cVar1S18S32P061P059P032N067(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='0' AND A(20)='1' AND B(21)='0' )then
          cVar1S19S32P061N059P018P034(0) <='1';
          else
          cVar1S19S32P061N059P018P034(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='0' AND A(20)='1' AND B(21)='0' )then
          cVar1S20S32P061N059P018P034(0) <='1';
          else
          cVar1S20S32P061N059P018P034(0) <='0';
          end if;
        if(E(18)='1' AND D(18)='0' AND A(20)='0' AND D(17)='1' )then
          cVar1S21S32P061N059N018P063(0) <='1';
          else
          cVar1S21S32P061N059N018P063(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='0' AND D(11)='0' AND B(10)='1' )then
          cVar1S0S33P062P013P054P037(0) <='1';
          else
          cVar1S0S33P062P013P054P037(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='0' AND D(11)='0' AND B(10)='0' )then
          cVar1S1S33P062P013P054N037(0) <='1';
          else
          cVar1S1S33P062P013P054N037(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='0' AND D(11)='0' AND B(10)='0' )then
          cVar1S2S33P062P013P054N037(0) <='1';
          else
          cVar1S2S33P062P013P054N037(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='0' AND D(11)='1' AND E( 8)='0' )then
          cVar1S3S33P062P013P054P068(0) <='1';
          else
          cVar1S3S33P062P013P054P068(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='1' AND D(16)='0' AND D(18)='0' )then
          cVar1S4S33P062P013P067P059(0) <='1';
          else
          cVar1S4S33P062P013P067P059(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='1' AND D(16)='0' AND D(18)='0' )then
          cVar1S5S33P062P013P067P059(0) <='1';
          else
          cVar1S5S33P062P013P067P059(0) <='0';
          end if;
        if(D( 9)='1' AND A(13)='1' AND D(16)='1' AND A(14)='0' )then
          cVar1S6S33P062P013P067P011(0) <='1';
          else
          cVar1S6S33P062P013P067P011(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='1' AND B(28)='1' )then
          cVar1S7S33N062P041P020nsss(0) <='1';
          else
          cVar1S7S33N062P041P020nsss(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='1' AND B(28)='0' AND B(11)='0' )then
          cVar1S8S33N062P041N020P035(0) <='1';
          else
          cVar1S8S33N062P041N020P035(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='1' AND B(28)='0' AND B(11)='0' )then
          cVar1S9S33N062P041N020P035(0) <='1';
          else
          cVar1S9S33N062P041N020P035(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='1' AND E(18)='1' )then
          cVar1S10S33N062N041P033P061(0) <='1';
          else
          cVar1S10S33N062N041P033P061(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='1' AND E(18)='1' )then
          cVar1S11S33N062N041P033P061(0) <='1';
          else
          cVar1S11S33N062N041P033P061(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='1' AND E(18)='0' )then
          cVar1S12S33N062N041P033N061(0) <='1';
          else
          cVar1S12S33N062N041P033N061(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='1' AND E(18)='0' )then
          cVar1S13S33N062N041P033N061(0) <='1';
          else
          cVar1S13S33N062N041P033N061(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='1' AND E(18)='0' )then
          cVar1S14S33N062N041P033N061(0) <='1';
          else
          cVar1S14S33N062N041P033N061(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='0' AND D(23)='0' )then
          cVar1S15S33N062N041N033P039(0) <='1';
          else
          cVar1S15S33N062N041N033P039(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='0' AND D(23)='0' )then
          cVar1S16S33N062N041N033P039(0) <='1';
          else
          cVar1S16S33N062N041N033P039(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='0' AND D(23)='0' )then
          cVar1S17S33N062N041N033P039(0) <='1';
          else
          cVar1S17S33N062N041N033P039(0) <='0';
          end if;
        if(D( 9)='0' AND E(23)='0' AND B(12)='0' AND D(23)='1' )then
          cVar1S18S33N062N041N033P039(0) <='1';
          else
          cVar1S18S33N062N041N033P039(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='1' AND A(18)='0' )then
          cVar1S0S34P011P029P062P003(0) <='1';
          else
          cVar1S0S34P011P029P062P003(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='1' AND A(18)='0' )then
          cVar1S1S34P011P029P062P003(0) <='1';
          else
          cVar1S1S34P011P029P062P003(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='1' AND A(18)='1' )then
          cVar1S2S34P011P029P062P003(0) <='1';
          else
          cVar1S2S34P011P029P062P003(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='1' )then
          cVar1S3S34P011P029N062P059(0) <='1';
          else
          cVar1S3S34P011P029N062P059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='1' )then
          cVar1S4S34P011P029N062P059(0) <='1';
          else
          cVar1S4S34P011P029N062P059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='1' )then
          cVar1S5S34P011P029N062P059(0) <='1';
          else
          cVar1S5S34P011P029N062P059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='0' )then
          cVar1S6S34P011P029N062N059(0) <='1';
          else
          cVar1S6S34P011P029N062N059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='0' )then
          cVar1S7S34P011P029N062N059(0) <='1';
          else
          cVar1S7S34P011P029N062N059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='0' AND D( 9)='0' AND D(18)='0' )then
          cVar1S8S34P011P029N062N059(0) <='1';
          else
          cVar1S8S34P011P029N062N059(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='1' AND E(12)='1' )then
          cVar1S9S34P011P029P052nsss(0) <='1';
          else
          cVar1S9S34P011P029P052nsss(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='1' AND E(12)='0' AND A(27)='0' )then
          cVar1S10S34P011P029N052P004(0) <='1';
          else
          cVar1S10S34P011P029N052P004(0) <='0';
          end if;
        if(A(14)='0' AND B(14)='1' AND E(12)='0' AND A(27)='0' )then
          cVar1S11S34P011P029N052P004(0) <='1';
          else
          cVar1S11S34P011P029N052P004(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='0' AND B(22)='0' AND B(14)='1' )then
          cVar1S12S34P011P013P032P029(0) <='1';
          else
          cVar1S12S34P011P013P032P029(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='0' AND B(22)='0' AND B(14)='0' )then
          cVar1S13S34P011P013P032N029(0) <='1';
          else
          cVar1S13S34P011P013P032N029(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='0' AND B(22)='0' AND B(14)='0' )then
          cVar1S14S34P011P013P032N029(0) <='1';
          else
          cVar1S14S34P011P013P032N029(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='0' AND B(22)='0' AND B(14)='0' )then
          cVar1S15S34P011P013P032N029(0) <='1';
          else
          cVar1S15S34P011P013P032N029(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='1' AND A(27)='0' AND A(25)='0' )then
          cVar1S16S34P011P013P004P008(0) <='1';
          else
          cVar1S16S34P011P013P004P008(0) <='0';
          end if;
        if(A(14)='1' AND A(13)='1' AND A(27)='0' AND A(25)='1' )then
          cVar1S17S34P011P013P004P008(0) <='1';
          else
          cVar1S17S34P011P013P004P008(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='0' AND B(21)='0' AND D(11)='0' )then
          cVar1S0S35P015P022P034P054(0) <='1';
          else
          cVar1S0S35P015P022P034P054(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='0' AND B(21)='0' AND D(11)='0' )then
          cVar1S1S35P015P022P034P054(0) <='1';
          else
          cVar1S1S35P015P022P034P054(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='0' AND B(21)='0' AND D(11)='0' )then
          cVar1S2S35P015P022P034P054(0) <='1';
          else
          cVar1S2S35P015P022P034P054(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='0' AND B(21)='0' AND D(11)='1' )then
          cVar1S3S35P015P022P034P054(0) <='1';
          else
          cVar1S3S35P015P022P034P054(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='0' AND B(21)='1' AND E(14)='0' )then
          cVar1S4S35P015P022P034P044(0) <='1';
          else
          cVar1S4S35P015P022P034P044(0) <='0';
          end if;
        if(A(12)='1' AND B(27)='1' AND A(23)='1' AND A(22)='0' )then
          cVar1S5S35P015P022P012P014nsss(0) <='1';
          else
          cVar1S5S35P015P022P012P014nsss(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='1' AND D(22)='0' AND B(12)='0' )then
          cVar1S6S35N015P064P043P033(0) <='1';
          else
          cVar1S6S35N015P064P043P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='1' AND D(22)='0' AND B(12)='0' )then
          cVar1S7S35N015P064P043P033(0) <='1';
          else
          cVar1S7S35N015P064P043P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='1' AND D(22)='0' AND B(12)='0' )then
          cVar1S8S35N015P064P043P033(0) <='1';
          else
          cVar1S8S35N015P064P043P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='1' AND D(22)='0' AND B(12)='1' )then
          cVar1S9S35N015P064P043P033(0) <='1';
          else
          cVar1S9S35N015P064P043P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='1' )then
          cVar1S10S35N015N064P068P034(0) <='1';
          else
          cVar1S10S35N015N064P068P034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='1' )then
          cVar1S11S35N015N064P068P034(0) <='1';
          else
          cVar1S11S35N015N064P068P034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='1' )then
          cVar1S12S35N015N064P068P034(0) <='1';
          else
          cVar1S12S35N015N064P068P034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='0' )then
          cVar1S13S35N015N064P068N034(0) <='1';
          else
          cVar1S13S35N015N064P068N034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='0' )then
          cVar1S14S35N015N064P068N034(0) <='1';
          else
          cVar1S14S35N015N064P068N034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='0' )then
          cVar1S15S35N015N064P068N034(0) <='1';
          else
          cVar1S15S35N015N064P068N034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='0' AND B(21)='0' )then
          cVar1S16S35N015N064P068N034(0) <='1';
          else
          cVar1S16S35N015N064P068N034(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='1' AND A(14)='0' )then
          cVar1S17S35N015N064P068P011(0) <='1';
          else
          cVar1S17S35N015N064P068P011(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='1' AND A(14)='0' )then
          cVar1S18S35N015N064P068P011(0) <='1';
          else
          cVar1S18S35N015N064P068P011(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='1' AND A(14)='0' )then
          cVar1S19S35N015N064P068P011(0) <='1';
          else
          cVar1S19S35N015N064P068P011(0) <='0';
          end if;
        if(A(12)='0' AND E( 9)='0' AND E( 8)='1' AND A(14)='1' )then
          cVar1S20S35N015N064P068P011(0) <='1';
          else
          cVar1S20S35N015N064P068P011(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='1' )then
          cVar1S0S36P011P015P065P063(0) <='1';
          else
          cVar1S0S36P011P015P065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='1' )then
          cVar1S1S36P011P015P065P063(0) <='1';
          else
          cVar1S1S36P011P015P065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='1' )then
          cVar1S2S36P011P015P065P063(0) <='1';
          else
          cVar1S2S36P011P015P065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='0' )then
          cVar1S3S36P011P015P065N063(0) <='1';
          else
          cVar1S3S36P011P015P065N063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='0' )then
          cVar1S4S36P011P015P065N063(0) <='1';
          else
          cVar1S4S36P011P015P065N063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='1' AND D(17)='0' )then
          cVar1S5S36P011P015P065N063(0) <='1';
          else
          cVar1S5S36P011P015P065N063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='0' )then
          cVar1S6S36P011P015N065P063(0) <='1';
          else
          cVar1S6S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='0' )then
          cVar1S7S36P011P015N065P063(0) <='1';
          else
          cVar1S7S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='0' )then
          cVar1S8S36P011P015N065P063(0) <='1';
          else
          cVar1S8S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='0' )then
          cVar1S9S36P011P015N065P063(0) <='1';
          else
          cVar1S9S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='1' )then
          cVar1S10S36P011P015N065P063(0) <='1';
          else
          cVar1S10S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='0' AND E(17)='0' AND D(17)='1' )then
          cVar1S11S36P011P015N065P063(0) <='1';
          else
          cVar1S11S36P011P015N065P063(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='1' AND B(27)='0' AND D(18)='1' )then
          cVar1S12S36P011P015P022P059(0) <='1';
          else
          cVar1S12S36P011P015P022P059(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='1' AND B(27)='0' AND D(18)='0' )then
          cVar1S13S36P011P015P022N059(0) <='1';
          else
          cVar1S13S36P011P015P022N059(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='1' AND B(27)='0' AND D(18)='0' )then
          cVar1S14S36P011P015P022N059(0) <='1';
          else
          cVar1S14S36P011P015P022N059(0) <='0';
          end if;
        if(A(14)='0' AND A(12)='1' AND B(27)='0' AND D(18)='0' )then
          cVar1S15S36P011P015P022N059(0) <='1';
          else
          cVar1S15S36P011P015P022N059(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='0' AND B(14)='1' AND D(11)='1' )then
          cVar1S16S36P011P004P029P054nsss(0) <='1';
          else
          cVar1S16S36P011P004P029P054nsss(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='0' AND B(14)='1' AND D(11)='0' )then
          cVar1S17S36P011P004P029N054(0) <='1';
          else
          cVar1S17S36P011P004P029N054(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='0' AND B(14)='1' AND D(11)='0' )then
          cVar1S18S36P011P004P029N054(0) <='1';
          else
          cVar1S18S36P011P004P029N054(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='0' AND B(14)='0' AND A(28)='0' )then
          cVar1S19S36P011P004N029P002(0) <='1';
          else
          cVar1S19S36P011P004N029P002(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='0' AND B(14)='0' AND A(28)='1' )then
          cVar1S20S36P011P004N029P002(0) <='1';
          else
          cVar1S20S36P011P004N029P002(0) <='0';
          end if;
        if(A(14)='1' AND A(27)='1' AND A(29)='0' AND E(11)='0' )then
          cVar1S21S36P011P004P000P056(0) <='1';
          else
          cVar1S21S36P011P004P000P056(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='0' AND B(27)='0' AND A(26)='0' )then
          cVar1S0S37P015P031P022P006(0) <='1';
          else
          cVar1S0S37P015P031P022P006(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='0' AND B(27)='0' AND A(26)='0' )then
          cVar1S1S37P015P031P022P006(0) <='1';
          else
          cVar1S1S37P015P031P022P006(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='0' AND B(27)='0' AND A(26)='0' )then
          cVar1S2S37P015P031P022P006(0) <='1';
          else
          cVar1S2S37P015P031P022P006(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='0' AND B(27)='0' AND A(26)='1' )then
          cVar1S3S37P015P031P022P006(0) <='1';
          else
          cVar1S3S37P015P031P022P006(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='0' AND B(27)='1' AND A(23)='1' )then
          cVar1S4S37P015P031P022P012nsss(0) <='1';
          else
          cVar1S4S37P015P031P022P012nsss(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='1' AND A(27)='0' AND B(23)='0' )then
          cVar1S5S37P015P031P004P030(0) <='1';
          else
          cVar1S5S37P015P031P004P030(0) <='0';
          end if;
        if(A(12)='1' AND B(13)='1' AND A(27)='0' AND B(23)='0' )then
          cVar1S6S37P015P031P004P030(0) <='1';
          else
          cVar1S6S37P015P031P004P030(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='1' AND A(16)='0' AND E(12)='1' )then
          cVar1S7S37N015P065P007P052nsss(0) <='1';
          else
          cVar1S7S37N015P065P007P052nsss(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='1' AND A(16)='0' AND E(12)='0' )then
          cVar1S8S37N015P065P007N052(0) <='1';
          else
          cVar1S8S37N015P065P007N052(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='1' AND A(16)='0' AND E(12)='0' )then
          cVar1S9S37N015P065P007N052(0) <='1';
          else
          cVar1S9S37N015P065P007N052(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='1' AND A(16)='1' AND A(15)='0' )then
          cVar1S10S37N015P065P007P009(0) <='1';
          else
          cVar1S10S37N015P065P007P009(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='1' AND D(22)='1' )then
          cVar1S11S37N015N065P022P043nsss(0) <='1';
          else
          cVar1S11S37N015N065P022P043nsss(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='1' AND D(22)='0' )then
          cVar1S12S37N015N065P022N043(0) <='1';
          else
          cVar1S12S37N015N065P022N043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='0' )then
          cVar1S13S37N015N065N022P043(0) <='1';
          else
          cVar1S13S37N015N065N022P043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='0' )then
          cVar1S14S37N015N065N022P043(0) <='1';
          else
          cVar1S14S37N015N065N022P043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='0' )then
          cVar1S15S37N015N065N022P043(0) <='1';
          else
          cVar1S15S37N015N065N022P043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='1' )then
          cVar1S16S37N015N065N022P043(0) <='1';
          else
          cVar1S16S37N015N065N022P043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='1' )then
          cVar1S17S37N015N065N022P043(0) <='1';
          else
          cVar1S17S37N015N065N022P043(0) <='0';
          end if;
        if(A(12)='0' AND E(17)='0' AND B(27)='0' AND D(22)='1' )then
          cVar1S18S37N015N065N022P043(0) <='1';
          else
          cVar1S18S37N015N065N022P043(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='1' )then
          cVar1S0S38P006P024P015P014(0) <='1';
          else
          cVar1S0S38P006P024P015P014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='1' )then
          cVar1S1S38P006P024P015P014(0) <='1';
          else
          cVar1S1S38P006P024P015P014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='1' )then
          cVar1S2S38P006P024P015P014(0) <='1';
          else
          cVar1S2S38P006P024P015P014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S3S38P006P024P015N014(0) <='1';
          else
          cVar1S3S38P006P024P015N014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S4S38P006P024P015N014(0) <='1';
          else
          cVar1S4S38P006P024P015N014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S5S38P006P024P015N014(0) <='1';
          else
          cVar1S5S38P006P024P015N014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S6S38P006P024P015N014(0) <='1';
          else
          cVar1S6S38P006P024P015N014(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='1' AND E(20)='1' )then
          cVar1S7S38P006P024P015P053(0) <='1';
          else
          cVar1S7S38P006P024P015P053(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='1' AND E(20)='0' )then
          cVar1S8S38P006P024P015N053(0) <='1';
          else
          cVar1S8S38P006P024P015N053(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND A(12)='1' AND E(20)='0' )then
          cVar1S9S38P006P024P015N053(0) <='1';
          else
          cVar1S9S38P006P024P015N053(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(22)='0' AND D(21)='1' )then
          cVar1S10S38P006P024P014P047nsss(0) <='1';
          else
          cVar1S10S38P006P024P014P047nsss(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(22)='0' AND D(21)='0' )then
          cVar1S11S38P006P024P014N047(0) <='1';
          else
          cVar1S11S38P006P024P014N047(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(22)='0' AND D(21)='0' )then
          cVar1S12S38P006P024P014N047(0) <='1';
          else
          cVar1S12S38P006P024P014N047(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(22)='1' AND D(16)='0' )then
          cVar1S13S38P006P024P014P067(0) <='1';
          else
          cVar1S13S38P006P024P014P067(0) <='0';
          end if;
        if(A(26)='1' AND B(21)='0' AND B(26)='1' AND D(20)='0' )then
          cVar1S14S38P006P034P024P051(0) <='1';
          else
          cVar1S14S38P006P034P024P051(0) <='0';
          end if;
        if(A(26)='1' AND B(21)='0' AND B(26)='0' AND E(17)='0' )then
          cVar1S15S38P006P034N024P065(0) <='1';
          else
          cVar1S15S38P006P034N024P065(0) <='0';
          end if;
        if(A(26)='1' AND B(21)='0' AND B(26)='0' AND E(17)='0' )then
          cVar1S16S38P006P034N024P065(0) <='1';
          else
          cVar1S16S38P006P034N024P065(0) <='0';
          end if;
        if(A(26)='1' AND B(21)='0' AND B(26)='0' AND E(17)='1' )then
          cVar1S17S38P006P034N024P065(0) <='1';
          else
          cVar1S17S38P006P034N024P065(0) <='0';
          end if;
        if(A(26)='1' AND B(21)='1' AND B(20)='0' AND A(14)='0' )then
          cVar1S18S38P006P034P036P011(0) <='1';
          else
          cVar1S18S38P006P034P036P011(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='0' AND D(22)='0' )then
          cVar1S0S39P006P067P024P043(0) <='1';
          else
          cVar1S0S39P006P067P024P043(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='0' AND D(22)='0' )then
          cVar1S1S39P006P067P024P043(0) <='1';
          else
          cVar1S1S39P006P067P024P043(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='0' AND D(22)='0' )then
          cVar1S2S39P006P067P024P043(0) <='1';
          else
          cVar1S2S39P006P067P024P043(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='0' AND D(22)='0' )then
          cVar1S3S39P006P067P024P043(0) <='1';
          else
          cVar1S3S39P006P067P024P043(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='0' AND D(22)='1' )then
          cVar1S4S39P006P067P024P043(0) <='1';
          else
          cVar1S4S39P006P067P024P043(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='1' AND B(26)='1' AND A(22)='0' )then
          cVar1S5S39P006P067P024P014(0) <='1';
          else
          cVar1S5S39P006P067P024P014(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='1' AND E(22)='0' )then
          cVar1S6S39P006N067P015P045(0) <='1';
          else
          cVar1S6S39P006N067P015P045(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='1' AND E(22)='0' )then
          cVar1S7S39P006N067P015P045(0) <='1';
          else
          cVar1S7S39P006N067P015P045(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='1' AND E(22)='0' )then
          cVar1S8S39P006N067P015P045(0) <='1';
          else
          cVar1S8S39P006N067P015P045(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='1' AND E(22)='1' )then
          cVar1S9S39P006N067P015P045(0) <='1';
          else
          cVar1S9S39P006N067P015P045(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='0' AND A(22)='1' )then
          cVar1S10S39P006N067N015P014(0) <='1';
          else
          cVar1S10S39P006N067N015P014(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='0' AND A(22)='1' )then
          cVar1S11S39P006N067N015P014(0) <='1';
          else
          cVar1S11S39P006N067N015P014(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S12S39P006N067N015N014(0) <='1';
          else
          cVar1S12S39P006N067N015N014(0) <='0';
          end if;
        if(A(26)='0' AND D(16)='0' AND A(12)='0' AND A(22)='0' )then
          cVar1S13S39P006N067N015N014(0) <='1';
          else
          cVar1S13S39P006N067N015N014(0) <='0';
          end if;
        if(A(26)='1' AND D(20)='0' AND B(26)='1' AND A(14)='0' )then
          cVar1S14S39P006P051P024P011(0) <='1';
          else
          cVar1S14S39P006P051P024P011(0) <='0';
          end if;
        if(A(26)='1' AND D(20)='0' AND B(26)='1' AND A(14)='0' )then
          cVar1S15S39P006P051P024P011(0) <='1';
          else
          cVar1S15S39P006P051P024P011(0) <='0';
          end if;
        if(A(26)='1' AND D(20)='0' AND B(26)='0' AND E(17)='0' )then
          cVar1S16S39P006P051N024P065(0) <='1';
          else
          cVar1S16S39P006P051N024P065(0) <='0';
          end if;
        if(A(26)='1' AND D(20)='0' AND B(26)='0' AND E(17)='1' )then
          cVar1S17S39P006P051N024P065(0) <='1';
          else
          cVar1S17S39P006P051N024P065(0) <='0';
          end if;
        if(A(26)='1' AND D(20)='1' AND D(16)='0' AND A(22)='0' )then
          cVar1S18S39P006P051P067P014(0) <='1';
          else
          cVar1S18S39P006P051P067P014(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='1' )then
          cVar1S0S40P014P032P030P012(0) <='1';
          else
          cVar1S0S40P014P032P030P012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='1' )then
          cVar1S1S40P014P032P030P012(0) <='1';
          else
          cVar1S1S40P014P032P030P012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='1' )then
          cVar1S2S40P014P032P030P012(0) <='1';
          else
          cVar1S2S40P014P032P030P012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S3S40P014P032P030N012(0) <='1';
          else
          cVar1S3S40P014P032P030N012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S4S40P014P032P030N012(0) <='1';
          else
          cVar1S4S40P014P032P030N012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S5S40P014P032P030N012(0) <='1';
          else
          cVar1S5S40P014P032P030N012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='0' AND E(19)='0' )then
          cVar1S6S40P014P032N030P057(0) <='1';
          else
          cVar1S6S40P014P032N030P057(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='0' AND E(19)='0' )then
          cVar1S7S40P014P032N030P057(0) <='1';
          else
          cVar1S7S40P014P032N030P057(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='0' AND E(19)='0' )then
          cVar1S8S40P014P032N030P057(0) <='1';
          else
          cVar1S8S40P014P032N030P057(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='0' AND E(19)='1' )then
          cVar1S9S40P014P032N030P057(0) <='1';
          else
          cVar1S9S40P014P032N030P057(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='0' AND B(23)='0' AND E(19)='1' )then
          cVar1S10S40P014P032N030P057(0) <='1';
          else
          cVar1S10S40P014P032N030P057(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='1' AND A(24)='0' AND A(23)='1' )then
          cVar1S11S40P014P032P010P012(0) <='1';
          else
          cVar1S11S40P014P032P010P012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='1' AND A(24)='0' AND A(23)='1' )then
          cVar1S12S40P014P032P010P012(0) <='1';
          else
          cVar1S12S40P014P032P010P012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='1' AND A(24)='0' AND A(23)='0' )then
          cVar1S13S40P014P032P010N012(0) <='1';
          else
          cVar1S13S40P014P032P010N012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='1' AND A(24)='0' AND A(23)='0' )then
          cVar1S14S40P014P032P010N012(0) <='1';
          else
          cVar1S14S40P014P032P010N012(0) <='0';
          end if;
        if(A(22)='0' AND B(22)='1' AND A(24)='1' AND A(11)='1' )then
          cVar1S15S40P014P032P010P017(0) <='1';
          else
          cVar1S15S40P014P032P010P017(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(22)='1' )then
          cVar1S16S40P014P024P044P032(0) <='1';
          else
          cVar1S16S40P014P024P044P032(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(22)='1' )then
          cVar1S17S40P014P024P044P032(0) <='1';
          else
          cVar1S17S40P014P024P044P032(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(22)='0' )then
          cVar1S18S40P014P024P044N032(0) <='1';
          else
          cVar1S18S40P014P024P044N032(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(22)='0' )then
          cVar1S19S40P014P024P044N032(0) <='1';
          else
          cVar1S19S40P014P024P044N032(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(22)='0' )then
          cVar1S20S40P014P024P044N032(0) <='1';
          else
          cVar1S20S40P014P024P044N032(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='1' AND D( 9)='0' )then
          cVar1S21S40P014P024P044P062(0) <='1';
          else
          cVar1S21S40P014P024P044P062(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND D(11)='0' AND B(20)='0' )then
          cVar1S22S40P014P024P054P036(0) <='1';
          else
          cVar1S22S40P014P024P054P036(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='1' AND D(12)='1' )then
          cVar1S0S41P035P015P027P050nsss(0) <='1';
          else
          cVar1S0S41P035P015P027P050nsss(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S1S41P035P015P027N050(0) <='1';
          else
          cVar1S1S41P035P015P027N050(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='1' )then
          cVar1S2S41P035P015N027P022(0) <='1';
          else
          cVar1S2S41P035P015N027P022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='1' )then
          cVar1S3S41P035P015N027P022(0) <='1';
          else
          cVar1S3S41P035P015N027P022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='0' )then
          cVar1S4S41P035P015N027N022(0) <='1';
          else
          cVar1S4S41P035P015N027N022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='0' )then
          cVar1S5S41P035P015N027N022(0) <='1';
          else
          cVar1S5S41P035P015N027N022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='0' )then
          cVar1S6S41P035P015N027N022(0) <='1';
          else
          cVar1S6S41P035P015N027N022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='0' AND B(15)='0' AND B(27)='0' )then
          cVar1S7S41P035P015N027N022(0) <='1';
          else
          cVar1S7S41P035P015N027N022(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='1' AND E(18)='0' )then
          cVar1S8S41P035P015P026P061(0) <='1';
          else
          cVar1S8S41P035P015P026P061(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='1' AND E(18)='0' )then
          cVar1S9S41P035P015P026P061(0) <='1';
          else
          cVar1S9S41P035P015P026P061(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S10S41P035P015N026P062(0) <='1';
          else
          cVar1S10S41P035P015N026P062(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S11S41P035P015N026P062(0) <='1';
          else
          cVar1S11S41P035P015N026P062(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S12S41P035P015N026P062(0) <='1';
          else
          cVar1S12S41P035P015N026P062(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S13S41P035P015N026P062(0) <='1';
          else
          cVar1S13S41P035P015N026P062(0) <='0';
          end if;
        if(B(11)='0' AND A(12)='1' AND B(25)='0' AND D( 9)='1' )then
          cVar1S14S41P035P015N026P062(0) <='1';
          else
          cVar1S14S41P035P015N026P062(0) <='0';
          end if;
        if(B(11)='1' AND E(22)='0' AND A(26)='0' AND D(17)='1' )then
          cVar1S15S41P035P045P006P063(0) <='1';
          else
          cVar1S15S41P035P045P006P063(0) <='0';
          end if;
        if(B(11)='1' AND E(22)='0' AND A(26)='0' AND D(17)='1' )then
          cVar1S16S41P035P045P006P063(0) <='1';
          else
          cVar1S16S41P035P045P006P063(0) <='0';
          end if;
        if(B(11)='1' AND E(22)='0' AND A(26)='0' AND D(17)='0' )then
          cVar1S17S41P035P045P006N063(0) <='1';
          else
          cVar1S17S41P035P045P006N063(0) <='0';
          end if;
        if(B(11)='1' AND E(22)='0' AND A(26)='0' AND D(17)='0' )then
          cVar1S18S41P035P045P006N063(0) <='1';
          else
          cVar1S18S41P035P045P006N063(0) <='0';
          end if;
        if(B(11)='1' AND E(22)='0' AND A(26)='1' AND B(21)='0' )then
          cVar1S19S41P035P045P006P034(0) <='1';
          else
          cVar1S19S41P035P045P006P034(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='0' )then
          cVar1S0S42P015P035P001P002(0) <='1';
          else
          cVar1S0S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='0' )then
          cVar1S1S42P015P035P001P002(0) <='1';
          else
          cVar1S1S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='0' )then
          cVar1S2S42P015P035P001P002(0) <='1';
          else
          cVar1S2S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='0' )then
          cVar1S3S42P015P035P001P002(0) <='1';
          else
          cVar1S3S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='1' )then
          cVar1S4S42P015P035P001P002(0) <='1';
          else
          cVar1S4S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='0' AND A(28)='1' )then
          cVar1S5S42P015P035P001P002(0) <='1';
          else
          cVar1S5S42P015P035P001P002(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='0' AND A(19)='1' AND A(13)='0' )then
          cVar1S6S42P015P035P001P013(0) <='1';
          else
          cVar1S6S42P015P035P001P013(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='1' AND B(28)='0' AND E(22)='0' )then
          cVar1S7S42P015P035P020P045(0) <='1';
          else
          cVar1S7S42P015P035P020P045(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='1' AND B(28)='0' AND E(22)='0' )then
          cVar1S8S42P015P035P020P045(0) <='1';
          else
          cVar1S8S42P015P035P020P045(0) <='0';
          end if;
        if(A(12)='0' AND B(11)='1' AND B(28)='0' AND E(22)='0' )then
          cVar1S9S42P015P035P020P045(0) <='1';
          else
          cVar1S9S42P015P035P020P045(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='1' )then
          cVar1S10S42P015P009P034P055(0) <='1';
          else
          cVar1S10S42P015P009P034P055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='1' )then
          cVar1S11S42P015P009P034P055(0) <='1';
          else
          cVar1S11S42P015P009P034P055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='1' )then
          cVar1S12S42P015P009P034P055(0) <='1';
          else
          cVar1S12S42P015P009P034P055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='0' )then
          cVar1S13S42P015P009P034N055(0) <='1';
          else
          cVar1S13S42P015P009P034N055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='0' )then
          cVar1S14S42P015P009P034N055(0) <='1';
          else
          cVar1S14S42P015P009P034N055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='0' AND D(19)='0' )then
          cVar1S15S42P015P009P034N055(0) <='1';
          else
          cVar1S15S42P015P009P034N055(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S16S42P015P009P034P063(0) <='1';
          else
          cVar1S16S42P015P009P034P063(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S17S42P015P009P034P063(0) <='1';
          else
          cVar1S17S42P015P009P034P063(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='1' AND D(17)='1' )then
          cVar1S18S42P015P009P034P063(0) <='1';
          else
          cVar1S18S42P015P009P034P063(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='0' AND B(21)='1' AND D(17)='0' )then
          cVar1S19S42P015P009P034N063(0) <='1';
          else
          cVar1S19S42P015P009P034N063(0) <='0';
          end if;
        if(A(12)='1' AND A(15)='1' AND E(23)='0' AND A(27)='0' )then
          cVar1S20S42P015P009P041P004(0) <='1';
          else
          cVar1S20S42P015P009P041P004(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='0' AND A(21)='0' )then
          cVar1S0S43P015P034P022P016(0) <='1';
          else
          cVar1S0S43P015P034P022P016(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='0' AND A(21)='0' )then
          cVar1S1S43P015P034P022P016(0) <='1';
          else
          cVar1S1S43P015P034P022P016(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='0' AND A(21)='0' )then
          cVar1S2S43P015P034P022P016(0) <='1';
          else
          cVar1S2S43P015P034P022P016(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='0' AND A(21)='1' )then
          cVar1S3S43P015P034P022P016(0) <='1';
          else
          cVar1S3S43P015P034P022P016(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='0' AND A(21)='1' )then
          cVar1S4S43P015P034P022P016(0) <='1';
          else
          cVar1S4S43P015P034P022P016(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='0' AND B(27)='1' AND A(15)='0' )then
          cVar1S5S43P015P034P022P009(0) <='1';
          else
          cVar1S5S43P015P034P022P009(0) <='0';
          end if;
        if(A(12)='1' AND B(21)='1' AND D(22)='0' AND E(14)='0' )then
          cVar1S6S43P015P034P043P044(0) <='1';
          else
          cVar1S6S43P015P034P043P044(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='1' AND E(13)='1' )then
          cVar1S7S43N015P027P048nsss(0) <='1';
          else
          cVar1S7S43N015P027P048nsss(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='1' AND E(13)='0' AND A(17)='0' )then
          cVar1S8S43N015P027N048P005(0) <='1';
          else
          cVar1S8S43N015P027N048P005(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='1' AND E(13)='0' AND A(17)='0' )then
          cVar1S9S43N015P027N048P005(0) <='1';
          else
          cVar1S9S43N015P027N048P005(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='1' AND A(23)='1' )then
          cVar1S10S43N015N027P030P012(0) <='1';
          else
          cVar1S10S43N015N027P030P012(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S11S43N015N027P030N012(0) <='1';
          else
          cVar1S11S43N015N027P030N012(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S12S43N015N027P030N012(0) <='1';
          else
          cVar1S12S43N015N027P030N012(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='1' AND A(23)='0' )then
          cVar1S13S43N015N027P030N012(0) <='1';
          else
          cVar1S13S43N015N027P030N012(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='0' AND E(15)='1' )then
          cVar1S14S43N015N027N030P040(0) <='1';
          else
          cVar1S14S43N015N027N030P040(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='0' AND E(15)='1' )then
          cVar1S15S43N015N027N030P040(0) <='1';
          else
          cVar1S15S43N015N027N030P040(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='0' AND E(15)='1' )then
          cVar1S16S43N015N027N030P040(0) <='1';
          else
          cVar1S16S43N015N027N030P040(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND B(23)='0' AND E(15)='0' )then
          cVar1S17S43N015N027N030N040(0) <='1';
          else
          cVar1S17S43N015N027N030N040(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='1' AND A(29)='0' AND E(13)='1' )then
          cVar1S0S44P015P027P000P048nsss(0) <='1';
          else
          cVar1S0S44P015P027P000P048nsss(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='1' AND A(29)='0' AND E(13)='0' )then
          cVar1S1S44P015P027P000N048(0) <='1';
          else
          cVar1S1S44P015P027P000N048(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='0' )then
          cVar1S2S44P015N027P018P068(0) <='1';
          else
          cVar1S2S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='0' )then
          cVar1S3S44P015N027P018P068(0) <='1';
          else
          cVar1S3S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='0' )then
          cVar1S4S44P015N027P018P068(0) <='1';
          else
          cVar1S4S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='1' )then
          cVar1S5S44P015N027P018P068(0) <='1';
          else
          cVar1S5S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='1' )then
          cVar1S6S44P015N027P018P068(0) <='1';
          else
          cVar1S6S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='0' AND E( 8)='1' )then
          cVar1S7S44P015N027P018P068(0) <='1';
          else
          cVar1S7S44P015N027P018P068(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='1' )then
          cVar1S8S44P015N027P018P013(0) <='1';
          else
          cVar1S8S44P015N027P018P013(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='1' )then
          cVar1S9S44P015N027P018P013(0) <='1';
          else
          cVar1S9S44P015N027P018P013(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='1' )then
          cVar1S10S44P015N027P018P013(0) <='1';
          else
          cVar1S10S44P015N027P018P013(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='0' )then
          cVar1S11S44P015N027P018N013(0) <='1';
          else
          cVar1S11S44P015N027P018N013(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='0' )then
          cVar1S12S44P015N027P018N013(0) <='1';
          else
          cVar1S12S44P015N027P018N013(0) <='0';
          end if;
        if(A(12)='0' AND B(15)='0' AND A(20)='1' AND A(13)='0' )then
          cVar1S13S44P015N027P018N013(0) <='1';
          else
          cVar1S13S44P015N027P018N013(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(20)='0' )then
          cVar1S14S44P015P051P068P036(0) <='1';
          else
          cVar1S14S44P015P051P068P036(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(20)='0' )then
          cVar1S15S44P015P051P068P036(0) <='1';
          else
          cVar1S15S44P015P051P068P036(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(20)='0' )then
          cVar1S16S44P015P051P068P036(0) <='1';
          else
          cVar1S16S44P015P051P068P036(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(20)='1' )then
          cVar1S17S44P015P051P068P036(0) <='1';
          else
          cVar1S17S44P015P051P068P036(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='1' AND A(20)='1' )then
          cVar1S18S44P015P051P068P018(0) <='1';
          else
          cVar1S18S44P015P051P068P018(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='1' AND A(20)='0' )then
          cVar1S19S44P015P051P068N018(0) <='1';
          else
          cVar1S19S44P015P051P068N018(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='1' AND A(20)='0' )then
          cVar1S20S44P015P051P068N018(0) <='1';
          else
          cVar1S20S44P015P051P068N018(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='1' AND A(29)='0' )then
          cVar1S21S44P015P051P053P000(0) <='1';
          else
          cVar1S21S44P015P051P053P000(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='0' AND E(21)='1' )then
          cVar1S22S44P015P051N053P049(0) <='1';
          else
          cVar1S22S44P015P051N053P049(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='0' )then
          cVar1S0S45P015P018P030P056(0) <='1';
          else
          cVar1S0S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='0' )then
          cVar1S1S45P015P018P030P056(0) <='1';
          else
          cVar1S1S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='0' )then
          cVar1S2S45P015P018P030P056(0) <='1';
          else
          cVar1S2S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='0' )then
          cVar1S3S45P015P018P030P056(0) <='1';
          else
          cVar1S3S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='1' )then
          cVar1S4S45P015P018P030P056(0) <='1';
          else
          cVar1S4S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='0' AND E(11)='1' )then
          cVar1S5S45P015P018P030P056(0) <='1';
          else
          cVar1S5S45P015P018P030P056(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='1' AND E(16)='1' )then
          cVar1S6S45P015P018P030P069nsss(0) <='1';
          else
          cVar1S6S45P015P018P030P069nsss(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='1' AND B(23)='1' AND E(16)='0' )then
          cVar1S7S45P015P018P030N069(0) <='1';
          else
          cVar1S7S45P015P018P030N069(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S8S45P015N018P019P017(0) <='1';
          else
          cVar1S8S45P015N018P019P017(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S9S45P015N018P019P017(0) <='1';
          else
          cVar1S9S45P015N018P019P017(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='1' AND A(11)='0' )then
          cVar1S10S45P015N018P019P017(0) <='1';
          else
          cVar1S10S45P015N018P019P017(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='1' AND A(11)='1' )then
          cVar1S11S45P015N018P019P017(0) <='1';
          else
          cVar1S11S45P015N018P019P017(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='1' AND A(11)='1' )then
          cVar1S12S45P015N018P019P017(0) <='1';
          else
          cVar1S12S45P015N018P019P017(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='0' AND D(16)='0' )then
          cVar1S13S45P015N018N019P067(0) <='1';
          else
          cVar1S13S45P015N018N019P067(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='0' AND D(16)='0' )then
          cVar1S14S45P015N018N019P067(0) <='1';
          else
          cVar1S14S45P015N018N019P067(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='0' AND D(16)='0' )then
          cVar1S15S45P015N018N019P067(0) <='1';
          else
          cVar1S15S45P015N018N019P067(0) <='0';
          end if;
        if(A(12)='0' AND A(20)='0' AND A(10)='0' AND D(16)='0' )then
          cVar1S16S45P015N018N019P067(0) <='1';
          else
          cVar1S16S45P015N018N019P067(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(27)='0' )then
          cVar1S17S45P015P051P068P022(0) <='1';
          else
          cVar1S17S45P015P051P068P022(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='0' AND B(27)='1' )then
          cVar1S18S45P015P051P068P022(0) <='1';
          else
          cVar1S18S45P015P051P068P022(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='1' AND A(20)='1' )then
          cVar1S19S45P015P051P068P018(0) <='1';
          else
          cVar1S19S45P015P051P068P018(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND E( 8)='1' AND A(20)='0' )then
          cVar1S20S45P015P051P068N018(0) <='1';
          else
          cVar1S20S45P015P051P068N018(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='1' AND A(29)='0' )then
          cVar1S21S45P015P051P053P000(0) <='1';
          else
          cVar1S21S45P015P051P053P000(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='0' AND E(21)='1' )then
          cVar1S22S45P015P051N053P049(0) <='1';
          else
          cVar1S22S45P015P051N053P049(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='1' AND B(23)='1' )then
          cVar1S0S46P068P019P057P030(0) <='1';
          else
          cVar1S0S46P068P019P057P030(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='1' AND B(23)='0' )then
          cVar1S1S46P068P019P057N030(0) <='1';
          else
          cVar1S1S46P068P019P057N030(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='1' AND B(23)='0' )then
          cVar1S2S46P068P019P057N030(0) <='1';
          else
          cVar1S2S46P068P019P057N030(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='1' )then
          cVar1S3S46P068P019N057P005(0) <='1';
          else
          cVar1S3S46P068P019N057P005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='1' )then
          cVar1S4S46P068P019N057P005(0) <='1';
          else
          cVar1S4S46P068P019N057P005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='0' )then
          cVar1S5S46P068P019N057N005(0) <='1';
          else
          cVar1S5S46P068P019N057N005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='0' )then
          cVar1S6S46P068P019N057N005(0) <='1';
          else
          cVar1S6S46P068P019N057N005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='0' )then
          cVar1S7S46P068P019N057N005(0) <='1';
          else
          cVar1S7S46P068P019N057N005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='0' AND E(19)='0' AND A(17)='0' )then
          cVar1S8S46P068P019N057N005(0) <='1';
          else
          cVar1S8S46P068P019N057N005(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND A(26)='0' AND D(22)='0' )then
          cVar1S9S46P068P019P006P043(0) <='1';
          else
          cVar1S9S46P068P019P006P043(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND A(26)='0' AND D(22)='0' )then
          cVar1S10S46P068P019P006P043(0) <='1';
          else
          cVar1S10S46P068P019P006P043(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND A(26)='0' AND D(22)='1' )then
          cVar1S11S46P068P019P006P043(0) <='1';
          else
          cVar1S11S46P068P019P006P043(0) <='0';
          end if;
        if(E( 8)='0' AND A(10)='1' AND A(26)='1' AND E(10)='0' )then
          cVar1S12S46P068P019P006P060(0) <='1';
          else
          cVar1S12S46P068P019P006P060(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='1' AND E(20)='0' )then
          cVar1S13S46P068P009P064P053(0) <='1';
          else
          cVar1S13S46P068P009P064P053(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='1' AND E(20)='0' )then
          cVar1S14S46P068P009P064P053(0) <='1';
          else
          cVar1S14S46P068P009P064P053(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='1' AND E(20)='0' )then
          cVar1S15S46P068P009P064P053(0) <='1';
          else
          cVar1S15S46P068P009P064P053(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='0' AND E(11)='1' )then
          cVar1S16S46P068P009N064P056(0) <='1';
          else
          cVar1S16S46P068P009N064P056(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='0' AND E(11)='1' )then
          cVar1S17S46P068P009N064P056(0) <='1';
          else
          cVar1S17S46P068P009N064P056(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='0' AND E(11)='0' )then
          cVar1S18S46P068P009N064N056(0) <='1';
          else
          cVar1S18S46P068P009N064N056(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND E( 9)='0' AND E(11)='0' )then
          cVar1S19S46P068P009N064N056(0) <='1';
          else
          cVar1S19S46P068P009N064N056(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='1' AND A(28)='0' AND D( 8)='1' )then
          cVar1S20S46P068P009P002P066(0) <='1';
          else
          cVar1S20S46P068P009P002P066(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='1' AND A(28)='0' AND D( 8)='1' )then
          cVar1S21S46P068P009P002P066(0) <='1';
          else
          cVar1S21S46P068P009P002P066(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND A(26)='0' AND D(22)='0' )then
          cVar1S0S47P019P033P006P043(0) <='1';
          else
          cVar1S0S47P019P033P006P043(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND A(26)='0' AND D(22)='0' )then
          cVar1S1S47P019P033P006P043(0) <='1';
          else
          cVar1S1S47P019P033P006P043(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND A(26)='0' AND D(22)='1' )then
          cVar1S2S47P019P033P006P043(0) <='1';
          else
          cVar1S2S47P019P033P006P043(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND A(26)='1' AND A(24)='0' )then
          cVar1S3S47P019P033P006P010(0) <='1';
          else
          cVar1S3S47P019P033P006P010(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND A(26)='1' AND A(24)='1' )then
          cVar1S4S47P019P033P006P010(0) <='1';
          else
          cVar1S4S47P019P033P006P010(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S5S47P019P033P016P065(0) <='1';
          else
          cVar1S5S47P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S6S47P019P033P016P065(0) <='1';
          else
          cVar1S6S47P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='1' )then
          cVar1S7S47P019P033P016P067(0) <='1';
          else
          cVar1S7S47P019P033P016P067(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='0' )then
          cVar1S8S47P019P033P016N067(0) <='1';
          else
          cVar1S8S47P019P033P016N067(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='1' AND E(23)='0' AND A(29)='0' )then
          cVar1S9S47N019P057P041P000(0) <='1';
          else
          cVar1S9S47N019P057P041P000(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='1' AND E(23)='0' AND A(29)='0' )then
          cVar1S10S47N019P057P041P000(0) <='1';
          else
          cVar1S10S47N019P057P041P000(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='1' AND E(23)='0' AND A(29)='0' )then
          cVar1S11S47N019P057P041P000(0) <='1';
          else
          cVar1S11S47N019P057P041P000(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='1' AND E(23)='0' AND A(29)='0' )then
          cVar1S12S47N019P057P041P000(0) <='1';
          else
          cVar1S12S47N019P057P041P000(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='0' )then
          cVar1S13S47N019N057P069P030(0) <='1';
          else
          cVar1S13S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='0' )then
          cVar1S14S47N019N057P069P030(0) <='1';
          else
          cVar1S14S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='0' )then
          cVar1S15S47N019N057P069P030(0) <='1';
          else
          cVar1S15S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='1' )then
          cVar1S16S47N019N057P069P030(0) <='1';
          else
          cVar1S16S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='1' )then
          cVar1S17S47N019N057P069P030(0) <='1';
          else
          cVar1S17S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='0' AND B(23)='1' )then
          cVar1S18S47N019N057P069P030(0) <='1';
          else
          cVar1S18S47N019N057P069P030(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='1' AND B(14)='1' )then
          cVar1S19S47N019N057P069P029(0) <='1';
          else
          cVar1S19S47N019N057P069P029(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='1' AND B(14)='0' )then
          cVar1S20S47N019N057P069N029(0) <='1';
          else
          cVar1S20S47N019N057P069N029(0) <='0';
          end if;
        if(A(10)='0' AND E(19)='0' AND E(16)='1' AND B(14)='0' )then
          cVar1S21S47N019N057P069N029(0) <='1';
          else
          cVar1S21S47N019N057P069N029(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='1' )then
          cVar1S0S48P019P069P061P007(0) <='1';
          else
          cVar1S0S48P019P069P061P007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='1' )then
          cVar1S1S48P019P069P061P007(0) <='1';
          else
          cVar1S1S48P019P069P061P007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='1' )then
          cVar1S2S48P019P069P061P007(0) <='1';
          else
          cVar1S2S48P019P069P061P007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='0' )then
          cVar1S3S48P019P069P061N007(0) <='1';
          else
          cVar1S3S48P019P069P061N007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='0' )then
          cVar1S4S48P019P069P061N007(0) <='1';
          else
          cVar1S4S48P019P069P061N007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='0' AND A(16)='0' )then
          cVar1S5S48P019P069P061N007(0) <='1';
          else
          cVar1S5S48P019P069P061N007(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='1' AND B(12)='1' )then
          cVar1S6S48P019P069P061P033(0) <='1';
          else
          cVar1S6S48P019P069P061P033(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='1' AND B(12)='0' )then
          cVar1S7S48P019P069P061N033(0) <='1';
          else
          cVar1S7S48P019P069P061N033(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='0' AND E(18)='1' AND B(12)='0' )then
          cVar1S8S48P019P069P061N033(0) <='1';
          else
          cVar1S8S48P019P069P061N033(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='1' AND E(22)='0' AND D(22)='0' )then
          cVar1S9S48P019P069P045P043(0) <='1';
          else
          cVar1S9S48P019P069P045P043(0) <='0';
          end if;
        if(A(10)='0' AND E(16)='1' AND E(22)='0' AND D(22)='0' )then
          cVar1S10S48P019P069P045P043(0) <='1';
          else
          cVar1S10S48P019P069P045P043(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='1' AND E(23)='0' AND A(18)='0' )then
          cVar1S11S48P019P059P041P003(0) <='1';
          else
          cVar1S11S48P019P059P041P003(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='0' AND B(12)='0' )then
          cVar1S12S48P019N059P061P033(0) <='1';
          else
          cVar1S12S48P019N059P061P033(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='0' AND B(12)='0' )then
          cVar1S13S48P019N059P061P033(0) <='1';
          else
          cVar1S13S48P019N059P061P033(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='0' AND B(12)='1' )then
          cVar1S14S48P019N059P061P033(0) <='1';
          else
          cVar1S14S48P019N059P061P033(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='0' AND B(12)='1' )then
          cVar1S15S48P019N059P061P033(0) <='1';
          else
          cVar1S15S48P019N059P061P033(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='1' AND A(20)='1' )then
          cVar1S16S48P019N059P061P018(0) <='1';
          else
          cVar1S16S48P019N059P061P018(0) <='0';
          end if;
        if(A(10)='1' AND D(18)='0' AND E(18)='1' AND A(20)='1' )then
          cVar1S17S48P019N059P061P018(0) <='1';
          else
          cVar1S17S48P019N059P061P018(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='0' AND A(13)='0' )then
          cVar1S0S49P019P033P057P013(0) <='1';
          else
          cVar1S0S49P019P033P057P013(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='0' AND A(13)='0' )then
          cVar1S1S49P019P033P057P013(0) <='1';
          else
          cVar1S1S49P019P033P057P013(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='0' AND A(13)='0' )then
          cVar1S2S49P019P033P057P013(0) <='1';
          else
          cVar1S2S49P019P033P057P013(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='0' AND A(13)='1' )then
          cVar1S3S49P019P033P057P013(0) <='1';
          else
          cVar1S3S49P019P033P057P013(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='1' AND B(23)='1' )then
          cVar1S4S49P019P033P057P030(0) <='1';
          else
          cVar1S4S49P019P033P057P030(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(19)='1' AND B(23)='0' )then
          cVar1S5S49P019P033P057N030(0) <='1';
          else
          cVar1S5S49P019P033P057N030(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S6S49P019P033P016P065(0) <='1';
          else
          cVar1S6S49P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S7S49P019P033P016P065(0) <='1';
          else
          cVar1S7S49P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='1' )then
          cVar1S8S49P019P033P016P067(0) <='1';
          else
          cVar1S8S49P019P033P016P067(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='0' )then
          cVar1S9S49P019P033P016N067(0) <='1';
          else
          cVar1S9S49P019P033P016N067(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='1' AND B(16)='1' )then
          cVar1S10S49N019P007P025nsss(0) <='1';
          else
          cVar1S10S49N019P007P025nsss(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='1' AND B(16)='0' AND D(18)='0' )then
          cVar1S11S49N019P007N025P059(0) <='1';
          else
          cVar1S11S49N019P007N025P059(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='1' AND B(16)='0' AND D(18)='0' )then
          cVar1S12S49N019P007N025P059(0) <='1';
          else
          cVar1S12S49N019P007N025P059(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='1' AND A(27)='0' )then
          cVar1S13S49N019N007P060P004(0) <='1';
          else
          cVar1S13S49N019N007P060P004(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='1' AND A(27)='0' )then
          cVar1S14S49N019N007P060P004(0) <='1';
          else
          cVar1S14S49N019N007P060P004(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='1' )then
          cVar1S15S49N019N007N060P057(0) <='1';
          else
          cVar1S15S49N019N007N060P057(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='1' )then
          cVar1S16S49N019N007N060P057(0) <='1';
          else
          cVar1S16S49N019N007N060P057(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='1' )then
          cVar1S17S49N019N007N060P057(0) <='1';
          else
          cVar1S17S49N019N007N060P057(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='1' )then
          cVar1S18S49N019N007N060P057(0) <='1';
          else
          cVar1S18S49N019N007N060P057(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='0' )then
          cVar1S19S49N019N007N060N057(0) <='1';
          else
          cVar1S19S49N019N007N060N057(0) <='0';
          end if;
        if(A(10)='0' AND A(16)='0' AND E(10)='0' AND E(19)='0' )then
          cVar1S20S49N019N007N060N057(0) <='1';
          else
          cVar1S20S49N019N007N060N057(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S0S50P019P014P027P009nsss(0) <='1';
          else
          cVar1S0S50P019P014P027P009nsss(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='1' AND A(15)='0' )then
          cVar1S1S50P019P014P027N009(0) <='1';
          else
          cVar1S1S50P019P014P027N009(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S2S50P019P014N027P050(0) <='1';
          else
          cVar1S2S50P019P014N027P050(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S3S50P019P014N027P050(0) <='1';
          else
          cVar1S3S50P019P014N027P050(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S4S50P019P014N027P050(0) <='1';
          else
          cVar1S4S50P019P014N027P050(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='0' AND B(15)='0' AND D(12)='1' )then
          cVar1S5S50P019P014N027P050(0) <='1';
          else
          cVar1S5S50P019P014N027P050(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='1' AND B(23)='0' AND D(17)='0' )then
          cVar1S6S50P019P014P030P063(0) <='1';
          else
          cVar1S6S50P019P014P030P063(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='1' AND B(23)='0' AND D(17)='0' )then
          cVar1S7S50P019P014P030P063(0) <='1';
          else
          cVar1S7S50P019P014P030P063(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='1' AND B(23)='0' AND D(17)='0' )then
          cVar1S8S50P019P014P030P063(0) <='1';
          else
          cVar1S8S50P019P014P030P063(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='1' AND B(23)='0' AND D(17)='1' )then
          cVar1S9S50P019P014P030P063(0) <='1';
          else
          cVar1S9S50P019P014P030P063(0) <='0';
          end if;
        if(A(10)='0' AND A(22)='1' AND B(23)='1' AND B(11)='1' )then
          cVar1S10S50P019P014P030P035nsss(0) <='1';
          else
          cVar1S10S50P019P014P030P035nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND A(13)='1' )then
          cVar1S11S50P019P002P020P013(0) <='1';
          else
          cVar1S11S50P019P002P020P013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND A(13)='1' )then
          cVar1S12S50P019P002P020P013(0) <='1';
          else
          cVar1S12S50P019P002P020P013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND A(13)='0' )then
          cVar1S13S50P019P002P020N013(0) <='1';
          else
          cVar1S13S50P019P002P020N013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND A(13)='0' )then
          cVar1S14S50P019P002P020N013(0) <='1';
          else
          cVar1S14S50P019P002P020N013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='1' AND A(13)='0' )then
          cVar1S15S50P019P002P020P013(0) <='1';
          else
          cVar1S15S50P019P002P020P013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='1' AND D(11)='0' AND A(15)='0' )then
          cVar1S16S50P019P002P054P009(0) <='1';
          else
          cVar1S16S50P019P002P054P009(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='1' AND D(11)='0' AND A(15)='0' )then
          cVar1S17S50P019P002P054P009(0) <='1';
          else
          cVar1S17S50P019P002P054P009(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND D(23)='0' )then
          cVar1S0S51P019P002P020P039(0) <='1';
          else
          cVar1S0S51P019P002P020P039(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND D(23)='0' )then
          cVar1S1S51P019P002P020P039(0) <='1';
          else
          cVar1S1S51P019P002P020P039(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='0' AND D(23)='1' )then
          cVar1S2S51P019P002P020P039(0) <='1';
          else
          cVar1S2S51P019P002P020P039(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='0' AND B(28)='1' AND A(13)='0' )then
          cVar1S3S51P019P002P020P013(0) <='1';
          else
          cVar1S3S51P019P002P020P013(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='1' AND D(11)='0' AND A(29)='0' )then
          cVar1S4S51P019P002P054P000(0) <='1';
          else
          cVar1S4S51P019P002P054P000(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='1' AND D(11)='0' AND A(29)='0' )then
          cVar1S5S51P019P002P054P000(0) <='1';
          else
          cVar1S5S51P019P002P054P000(0) <='0';
          end if;
        if(A(10)='1' AND A(28)='1' AND D(11)='0' AND A(29)='0' )then
          cVar1S6S51P019P002P054P000(0) <='1';
          else
          cVar1S6S51P019P002P054P000(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='1' AND D(14)='0' AND A(12)='0' )then
          cVar1S7S51N019P017P042P015(0) <='1';
          else
          cVar1S7S51N019P017P042P015(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='1' AND D(14)='0' AND A(12)='0' )then
          cVar1S8S51N019P017P042P015(0) <='1';
          else
          cVar1S8S51N019P017P042P015(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='1' AND D(14)='0' AND A(12)='0' )then
          cVar1S9S51N019P017P042P015(0) <='1';
          else
          cVar1S9S51N019P017P042P015(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='1' AND D(14)='0' AND A(12)='1' )then
          cVar1S10S51N019P017P042P015(0) <='1';
          else
          cVar1S10S51N019P017P042P015(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='1' AND B(17)='1' )then
          cVar1S11S51N019N017P005P023nsss(0) <='1';
          else
          cVar1S11S51N019N017P005P023nsss(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='1' AND B(17)='0' )then
          cVar1S12S51N019N017P005N023(0) <='1';
          else
          cVar1S12S51N019N017P005N023(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='1' AND B(17)='0' )then
          cVar1S13S51N019N017P005N023(0) <='1';
          else
          cVar1S13S51N019N017P005N023(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='0' )then
          cVar1S14S51N019N017N005P012(0) <='1';
          else
          cVar1S14S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='0' )then
          cVar1S15S51N019N017N005P012(0) <='1';
          else
          cVar1S15S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='0' )then
          cVar1S16S51N019N017N005P012(0) <='1';
          else
          cVar1S16S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='0' )then
          cVar1S17S51N019N017N005P012(0) <='1';
          else
          cVar1S17S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='1' )then
          cVar1S18S51N019N017N005P012(0) <='1';
          else
          cVar1S18S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='1' )then
          cVar1S19S51N019N017N005P012(0) <='1';
          else
          cVar1S19S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(11)='0' AND A(17)='0' AND A(23)='1' )then
          cVar1S20S51N019N017N005P012(0) <='1';
          else
          cVar1S20S51N019N017N005P012(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='1' )then
          cVar1S0S52P019P012P030P050(0) <='1';
          else
          cVar1S0S52P019P012P030P050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='1' )then
          cVar1S1S52P019P012P030P050(0) <='1';
          else
          cVar1S1S52P019P012P030P050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='0' )then
          cVar1S2S52P019P012P030N050(0) <='1';
          else
          cVar1S2S52P019P012P030N050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='0' )then
          cVar1S3S52P019P012P030N050(0) <='1';
          else
          cVar1S3S52P019P012P030N050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='0' )then
          cVar1S4S52P019P012P030N050(0) <='1';
          else
          cVar1S4S52P019P012P030N050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='0' AND D(12)='0' )then
          cVar1S5S52P019P012P030N050(0) <='1';
          else
          cVar1S5S52P019P012P030N050(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='1' AND A(24)='1' )then
          cVar1S6S52P019P012P030P010(0) <='1';
          else
          cVar1S6S52P019P012P030P010(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='1' AND A(24)='0' )then
          cVar1S7S52P019P012P030N010(0) <='1';
          else
          cVar1S7S52P019P012P030N010(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='0' AND B(23)='1' AND A(24)='0' )then
          cVar1S8S52P019P012P030N010(0) <='1';
          else
          cVar1S8S52P019P012P030N010(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='0' AND B(13)='1' )then
          cVar1S9S52P019P012P008P031(0) <='1';
          else
          cVar1S9S52P019P012P008P031(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='0' AND B(13)='1' )then
          cVar1S10S52P019P012P008P031(0) <='1';
          else
          cVar1S10S52P019P012P008P031(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='0' AND B(13)='0' )then
          cVar1S11S52P019P012P008N031(0) <='1';
          else
          cVar1S11S52P019P012P008N031(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='0' AND B(13)='0' )then
          cVar1S12S52P019P012P008N031(0) <='1';
          else
          cVar1S12S52P019P012P008N031(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='0' AND B(13)='0' )then
          cVar1S13S52P019P012P008N031(0) <='1';
          else
          cVar1S13S52P019P012P008N031(0) <='0';
          end if;
        if(A(10)='0' AND A(23)='1' AND A(25)='1' AND A(14)='0' )then
          cVar1S14S52P019P012P008P011(0) <='1';
          else
          cVar1S14S52P019P012P008P011(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND B(24)='1' )then
          cVar1S15S52P019P033P049P028(0) <='1';
          else
          cVar1S15S52P019P033P049P028(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND B(24)='1' )then
          cVar1S16S52P019P033P049P028(0) <='1';
          else
          cVar1S16S52P019P033P049P028(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='1' AND E( 8)='1' )then
          cVar1S17S52P019P033P049P068(0) <='1';
          else
          cVar1S17S52P019P033P049P068(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S18S52P019P033P016P065(0) <='1';
          else
          cVar1S18S52P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S19S52P019P033P016P065(0) <='1';
          else
          cVar1S19S52P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='1' )then
          cVar1S20S52P019P033P016P067(0) <='1';
          else
          cVar1S20S52P019P033P016P067(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND E(13)='0' )then
          cVar1S0S53P019P033P049P048(0) <='1';
          else
          cVar1S0S53P019P033P049P048(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND E(13)='0' )then
          cVar1S1S53P019P033P049P048(0) <='1';
          else
          cVar1S1S53P019P033P049P048(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND E(13)='1' )then
          cVar1S2S53P019P033P049P048(0) <='1';
          else
          cVar1S2S53P019P033P049P048(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='0' AND E(13)='1' )then
          cVar1S3S53P019P033P049P048(0) <='1';
          else
          cVar1S3S53P019P033P049P048(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='1' AND E( 8)='1' )then
          cVar1S4S53P019P033P049P068(0) <='1';
          else
          cVar1S4S53P019P033P049P068(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(21)='1' AND E( 8)='1' )then
          cVar1S5S53P019P033P049P068(0) <='1';
          else
          cVar1S5S53P019P033P049P068(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S6S53P019P033P016P065(0) <='1';
          else
          cVar1S6S53P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S7S53P019P033P016P065(0) <='1';
          else
          cVar1S7S53P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='1' )then
          cVar1S8S53P019P033P016P067(0) <='1';
          else
          cVar1S8S53P019P033P016P067(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='1' AND B(18)='0' AND B(15)='1' )then
          cVar1S9S53N019P050P021P027nsss(0) <='1';
          else
          cVar1S9S53N019P050P021P027nsss(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='1' AND B(18)='0' AND B(15)='0' )then
          cVar1S10S53N019P050P021N027(0) <='1';
          else
          cVar1S10S53N019P050P021N027(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='1' AND A(25)='0' )then
          cVar1S11S53N019N050P032P008(0) <='1';
          else
          cVar1S11S53N019N050P032P008(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='1' AND A(25)='0' )then
          cVar1S12S53N019N050P032P008(0) <='1';
          else
          cVar1S12S53N019N050P032P008(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='1' AND A(25)='0' )then
          cVar1S13S53N019N050P032P008(0) <='1';
          else
          cVar1S13S53N019N050P032P008(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='0' AND B(17)='1' )then
          cVar1S14S53N019N050N032P023(0) <='1';
          else
          cVar1S14S53N019N050N032P023(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='0' AND B(17)='1' )then
          cVar1S15S53N019N050N032P023(0) <='1';
          else
          cVar1S15S53N019N050N032P023(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='0' AND B(17)='0' )then
          cVar1S16S53N019N050N032N023(0) <='1';
          else
          cVar1S16S53N019N050N032N023(0) <='0';
          end if;
        if(A(10)='0' AND D(12)='0' AND B(22)='0' AND B(17)='0' )then
          cVar1S17S53N019N050N032N023(0) <='1';
          else
          cVar1S17S53N019N050N032N023(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='1' AND A(23)='1' )then
          cVar1S0S54P019P015P017P012(0) <='1';
          else
          cVar1S0S54P019P015P017P012(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='1' AND A(23)='0' )then
          cVar1S1S54P019P015P017N012(0) <='1';
          else
          cVar1S1S54P019P015P017N012(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='1' AND A(23)='0' )then
          cVar1S2S54P019P015P017N012(0) <='1';
          else
          cVar1S2S54P019P015P017N012(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='0' AND D(17)='0' )then
          cVar1S3S54P019P015N017P063(0) <='1';
          else
          cVar1S3S54P019P015N017P063(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='0' AND D(17)='0' )then
          cVar1S4S54P019P015N017P063(0) <='1';
          else
          cVar1S4S54P019P015N017P063(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='0' AND A(11)='0' AND D(17)='1' )then
          cVar1S5S54P019P015N017P063(0) <='1';
          else
          cVar1S5S54P019P015N017P063(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='0' AND E(18)='1' )then
          cVar1S6S54P019P015P017P061(0) <='1';
          else
          cVar1S6S54P019P015P017P061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='0' AND E(18)='1' )then
          cVar1S7S54P019P015P017P061(0) <='1';
          else
          cVar1S7S54P019P015P017P061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='0' AND E(18)='0' )then
          cVar1S8S54P019P015P017N061(0) <='1';
          else
          cVar1S8S54P019P015P017N061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='0' AND E(18)='0' )then
          cVar1S9S54P019P015P017N061(0) <='1';
          else
          cVar1S9S54P019P015P017N061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='0' AND E(18)='0' )then
          cVar1S10S54P019P015P017N061(0) <='1';
          else
          cVar1S10S54P019P015P017N061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='1' AND E(18)='0' )then
          cVar1S11S54P019P015P017P061(0) <='1';
          else
          cVar1S11S54P019P015P017P061(0) <='0';
          end if;
        if(A(10)='0' AND A(12)='1' AND A(11)='1' AND E(18)='1' )then
          cVar1S12S54P019P015P017P061(0) <='1';
          else
          cVar1S12S54P019P015P017P061(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='1' )then
          cVar1S13S54P019P033P060P017(0) <='1';
          else
          cVar1S13S54P019P033P060P017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='1' )then
          cVar1S14S54P019P033P060P017(0) <='1';
          else
          cVar1S14S54P019P033P060P017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='1' )then
          cVar1S15S54P019P033P060P017(0) <='1';
          else
          cVar1S15S54P019P033P060P017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='0' )then
          cVar1S16S54P019P033P060N017(0) <='1';
          else
          cVar1S16S54P019P033P060N017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='0' )then
          cVar1S17S54P019P033P060N017(0) <='1';
          else
          cVar1S17S54P019P033P060N017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='0' AND A(11)='0' )then
          cVar1S18S54P019P033P060N017(0) <='1';
          else
          cVar1S18S54P019P033P060N017(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='1' AND A(15)='0' )then
          cVar1S19S54P019P033P060P009(0) <='1';
          else
          cVar1S19S54P019P033P060P009(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='0' AND E(10)='1' AND A(15)='0' )then
          cVar1S20S54P019P033P060P009(0) <='1';
          else
          cVar1S20S54P019P033P060P009(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S21S54P019P033P016P065(0) <='1';
          else
          cVar1S21S54P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='0' AND E(17)='0' )then
          cVar1S22S54P019P033P016P065(0) <='1';
          else
          cVar1S22S54P019P033P016P065(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='1' )then
          cVar1S23S54P019P033P016P067(0) <='1';
          else
          cVar1S23S54P019P033P016P067(0) <='0';
          end if;
        if(A(10)='1' AND B(12)='1' AND A(21)='1' AND D(16)='0' )then
          cVar1S24S54P019P033P016N067(0) <='1';
          else
          cVar1S24S54P019P033P016N067(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='0' AND B(27)='0' )then
          cVar1S0S55P015P068P051P022(0) <='1';
          else
          cVar1S0S55P015P068P051P022(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='0' AND B(27)='0' )then
          cVar1S1S55P015P068P051P022(0) <='1';
          else
          cVar1S1S55P015P068P051P022(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='0' AND B(27)='0' )then
          cVar1S2S55P015P068P051P022(0) <='1';
          else
          cVar1S2S55P015P068P051P022(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='0' AND B(27)='0' )then
          cVar1S3S55P015P068P051P022(0) <='1';
          else
          cVar1S3S55P015P068P051P022(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='0' AND B(27)='1' )then
          cVar1S4S55P015P068P051P022(0) <='1';
          else
          cVar1S4S55P015P068P051P022(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='1' AND E(20)='1' )then
          cVar1S5S55P015P068P051P053(0) <='1';
          else
          cVar1S5S55P015P068P051P053(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='1' AND E(20)='1' )then
          cVar1S6S55P015P068P051P053(0) <='1';
          else
          cVar1S6S55P015P068P051P053(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='0' AND D(20)='1' AND E(20)='0' )then
          cVar1S7S55P015P068P051N053(0) <='1';
          else
          cVar1S7S55P015P068P051N053(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='1' AND A(15)='0' AND A(24)='1' )then
          cVar1S8S55P015P068P009P010(0) <='1';
          else
          cVar1S8S55P015P068P009P010(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='1' AND A(15)='0' AND A(24)='0' )then
          cVar1S9S55P015P068P009N010(0) <='1';
          else
          cVar1S9S55P015P068P009N010(0) <='0';
          end if;
        if(A(12)='1' AND E( 8)='1' AND A(15)='1' AND D( 8)='1' )then
          cVar1S10S55P015P068P009P066(0) <='1';
          else
          cVar1S10S55P015P068P009P066(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S11S55N015P068P003P033(0) <='1';
          else
          cVar1S11S55N015P068P003P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='1' AND A(18)='0' AND B(12)='0' )then
          cVar1S12S55N015P068P003P033(0) <='1';
          else
          cVar1S12S55N015P068P003P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='1' AND A(18)='0' AND B(12)='1' )then
          cVar1S13S55N015P068P003P033(0) <='1';
          else
          cVar1S13S55N015P068P003P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='1' AND A(18)='0' AND B(12)='1' )then
          cVar1S14S55N015P068P003P033(0) <='1';
          else
          cVar1S14S55N015P068P003P033(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='1' AND A(18)='1' AND E(17)='0' )then
          cVar1S15S55N015P068P003P065(0) <='1';
          else
          cVar1S15S55N015P068P003P065(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='1' AND A(25)='0' )then
          cVar1S16S55N015N068P069P008(0) <='1';
          else
          cVar1S16S55N015N068P069P008(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='1' AND A(25)='0' )then
          cVar1S17S55N015N068P069P008(0) <='1';
          else
          cVar1S17S55N015N068P069P008(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='1' AND A(25)='0' )then
          cVar1S18S55N015N068P069P008(0) <='1';
          else
          cVar1S18S55N015N068P069P008(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='1' AND A(25)='1' )then
          cVar1S19S55N015N068P069P008(0) <='1';
          else
          cVar1S19S55N015N068P069P008(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='0' AND A(27)='1' )then
          cVar1S20S55N015N068N069P004(0) <='1';
          else
          cVar1S20S55N015N068N069P004(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='0' AND A(27)='1' )then
          cVar1S21S55N015N068N069P004(0) <='1';
          else
          cVar1S21S55N015N068N069P004(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='0' AND A(27)='0' )then
          cVar1S22S55N015N068N069N004(0) <='1';
          else
          cVar1S22S55N015N068N069N004(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='0' AND A(27)='0' )then
          cVar1S23S55N015N068N069N004(0) <='1';
          else
          cVar1S23S55N015N068N069N004(0) <='0';
          end if;
        if(A(12)='0' AND E( 8)='0' AND E(16)='0' AND A(27)='0' )then
          cVar1S24S55N015N068N069N004(0) <='1';
          else
          cVar1S24S55N015N068N069N004(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='1' )then
          cVar1S0S56P068P015P066P034(0) <='1';
          else
          cVar1S0S56P068P015P066P034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='1' )then
          cVar1S1S56P068P015P066P034(0) <='1';
          else
          cVar1S1S56P068P015P066P034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='1' )then
          cVar1S2S56P068P015P066P034(0) <='1';
          else
          cVar1S2S56P068P015P066P034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='0' )then
          cVar1S3S56P068P015P066N034(0) <='1';
          else
          cVar1S3S56P068P015P066N034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='0' )then
          cVar1S4S56P068P015P066N034(0) <='1';
          else
          cVar1S4S56P068P015P066N034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='0' )then
          cVar1S5S56P068P015P066N034(0) <='1';
          else
          cVar1S5S56P068P015P066N034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='0' AND B(21)='0' )then
          cVar1S6S56P068P015P066N034(0) <='1';
          else
          cVar1S6S56P068P015P066N034(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='0' AND D( 8)='1' AND A(25)='0' )then
          cVar1S7S56P068P015P066P008(0) <='1';
          else
          cVar1S7S56P068P015P066P008(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='0' AND B(27)='0' )then
          cVar1S8S56P068P015P051P022(0) <='1';
          else
          cVar1S8S56P068P015P051P022(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='0' AND B(27)='0' )then
          cVar1S9S56P068P015P051P022(0) <='1';
          else
          cVar1S9S56P068P015P051P022(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='0' AND B(27)='0' )then
          cVar1S10S56P068P015P051P022(0) <='1';
          else
          cVar1S10S56P068P015P051P022(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='0' AND B(27)='1' )then
          cVar1S11S56P068P015P051P022(0) <='1';
          else
          cVar1S11S56P068P015P051P022(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='1' AND E(20)='1' )then
          cVar1S12S56P068P015P051P053(0) <='1';
          else
          cVar1S12S56P068P015P051P053(0) <='0';
          end if;
        if(E( 8)='0' AND A(12)='1' AND D(20)='1' AND E(20)='0' )then
          cVar1S13S56P068P015P051N053(0) <='1';
          else
          cVar1S13S56P068P015P051N053(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='0' AND E(12)='1' )then
          cVar1S14S56P068P009P024P052(0) <='1';
          else
          cVar1S14S56P068P009P024P052(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='0' AND E(12)='1' )then
          cVar1S15S56P068P009P024P052(0) <='1';
          else
          cVar1S15S56P068P009P024P052(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='0' AND E(12)='0' )then
          cVar1S16S56P068P009P024N052(0) <='1';
          else
          cVar1S16S56P068P009P024N052(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='0' AND E(12)='0' )then
          cVar1S17S56P068P009P024N052(0) <='1';
          else
          cVar1S17S56P068P009P024N052(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='1' AND A(26)='1' )then
          cVar1S18S56P068P009P024P006nsss(0) <='1';
          else
          cVar1S18S56P068P009P024P006nsss(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='0' AND B(26)='1' AND A(26)='0' )then
          cVar1S19S56P068P009P024N006(0) <='1';
          else
          cVar1S19S56P068P009P024N006(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='1' AND A(28)='0' AND D( 8)='1' )then
          cVar1S20S56P068P009P002P066(0) <='1';
          else
          cVar1S20S56P068P009P002P066(0) <='0';
          end if;
        if(E( 8)='1' AND A(15)='1' AND A(28)='0' AND D( 8)='1' )then
          cVar1S21S56P068P009P002P066(0) <='1';
          else
          cVar1S21S56P068P009P002P066(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='0' )then
          cVar1S0S57P015P051P009P037(0) <='1';
          else
          cVar1S0S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='0' )then
          cVar1S1S57P015P051P009P037(0) <='1';
          else
          cVar1S1S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='0' )then
          cVar1S2S57P015P051P009P037(0) <='1';
          else
          cVar1S2S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='1' )then
          cVar1S3S57P015P051P009P037(0) <='1';
          else
          cVar1S3S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='1' )then
          cVar1S4S57P015P051P009P037(0) <='1';
          else
          cVar1S4S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='1' )then
          cVar1S5S57P015P051P009P037(0) <='1';
          else
          cVar1S5S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='0' AND B(10)='1' )then
          cVar1S6S57P015P051P009P037(0) <='1';
          else
          cVar1S6S57P015P051P009P037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='1' AND E( 8)='0' )then
          cVar1S7S57P015P051P009P068(0) <='1';
          else
          cVar1S7S57P015P051P009P068(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='1' AND E( 8)='0' )then
          cVar1S8S57P015P051P009P068(0) <='1';
          else
          cVar1S8S57P015P051P009P068(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='1' AND E( 8)='0' )then
          cVar1S9S57P015P051P009P068(0) <='1';
          else
          cVar1S9S57P015P051P009P068(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(15)='1' AND E( 8)='1' )then
          cVar1S10S57P015P051P009P068(0) <='1';
          else
          cVar1S10S57P015P051P009P068(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='1' AND A(29)='0' )then
          cVar1S11S57P015P051P053P000(0) <='1';
          else
          cVar1S11S57P015P051P053P000(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='0' AND A(22)='0' )then
          cVar1S12S57P015P051N053P014(0) <='1';
          else
          cVar1S12S57P015P051N053P014(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='1' AND A(26)='0' )then
          cVar1S13S57N015P033P034P006(0) <='1';
          else
          cVar1S13S57N015P033P034P006(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='1' AND A(26)='1' )then
          cVar1S14S57N015P033P034P006(0) <='1';
          else
          cVar1S14S57N015P033P034P006(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='0' AND B(15)='1' )then
          cVar1S15S57N015P033N034P027(0) <='1';
          else
          cVar1S15S57N015P033N034P027(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='0' AND B(15)='1' )then
          cVar1S16S57N015P033N034P027(0) <='1';
          else
          cVar1S16S57N015P033N034P027(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='0' AND B(15)='0' )then
          cVar1S17S57N015P033N034N027(0) <='1';
          else
          cVar1S17S57N015P033N034N027(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='0' AND B(15)='0' )then
          cVar1S18S57N015P033N034N027(0) <='1';
          else
          cVar1S18S57N015P033N034N027(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='0' AND B(21)='0' AND B(15)='0' )then
          cVar1S19S57N015P033N034N027(0) <='1';
          else
          cVar1S19S57N015P033N034N027(0) <='0';
          end if;
        if(A(12)='0' AND B(12)='1' AND E( 9)='0' AND E(11)='0' )then
          cVar1S20S57N015P033P064P056(0) <='1';
          else
          cVar1S20S57N015P033P064P056(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='0' )then
          cVar1S0S58P066P015P033P018(0) <='1';
          else
          cVar1S0S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='0' )then
          cVar1S1S58P066P015P033P018(0) <='1';
          else
          cVar1S1S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='0' )then
          cVar1S2S58P066P015P033P018(0) <='1';
          else
          cVar1S2S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='0' )then
          cVar1S3S58P066P015P033P018(0) <='1';
          else
          cVar1S3S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='1' )then
          cVar1S4S58P066P015P033P018(0) <='1';
          else
          cVar1S4S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='1' )then
          cVar1S5S58P066P015P033P018(0) <='1';
          else
          cVar1S5S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='0' AND A(20)='1' )then
          cVar1S6S58P066P015P033P018(0) <='1';
          else
          cVar1S6S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='1' AND A(20)='1' )then
          cVar1S7S58P066P015P033P018(0) <='1';
          else
          cVar1S7S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='1' AND A(20)='1' )then
          cVar1S8S58P066P015P033P018(0) <='1';
          else
          cVar1S8S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='1' AND A(20)='1' )then
          cVar1S9S58P066P015P033P018(0) <='1';
          else
          cVar1S9S58P066P015P033P018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='0' AND B(12)='1' AND A(20)='0' )then
          cVar1S10S58P066P015P033N018(0) <='1';
          else
          cVar1S10S58P066P015P033N018(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='1' AND A(16)='0' AND E( 8)='0' )then
          cVar1S11S58P066P015P007P068(0) <='1';
          else
          cVar1S11S58P066P015P007P068(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='1' AND A(16)='0' AND E( 8)='0' )then
          cVar1S12S58P066P015P007P068(0) <='1';
          else
          cVar1S12S58P066P015P007P068(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='1' AND A(16)='0' AND E( 8)='0' )then
          cVar1S13S58P066P015P007P068(0) <='1';
          else
          cVar1S13S58P066P015P007P068(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='1' AND A(16)='0' AND E( 8)='1' )then
          cVar1S14S58P066P015P007P068(0) <='1';
          else
          cVar1S14S58P066P015P007P068(0) <='0';
          end if;
        if(D( 8)='0' AND A(12)='1' AND A(16)='1' AND D(18)='0' )then
          cVar1S15S58P066P015P007P059(0) <='1';
          else
          cVar1S15S58P066P015P007P059(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='0' AND B(26)='0' AND E(22)='0' )then
          cVar1S16S58P066P009P024P045(0) <='1';
          else
          cVar1S16S58P066P009P024P045(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='0' AND B(26)='0' AND E(22)='0' )then
          cVar1S17S58P066P009P024P045(0) <='1';
          else
          cVar1S17S58P066P009P024P045(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='0' AND B(26)='0' AND E(22)='1' )then
          cVar1S18S58P066P009P024P045(0) <='1';
          else
          cVar1S18S58P066P009P024P045(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='0' AND B(26)='1' AND E(20)='0' )then
          cVar1S19S58P066P009P024P053(0) <='1';
          else
          cVar1S19S58P066P009P024P053(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='1' AND A(28)='0' AND B(10)='1' )then
          cVar1S20S58P066P009P002P037(0) <='1';
          else
          cVar1S20S58P066P009P002P037(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='1' AND A(28)='0' AND B(10)='1' )then
          cVar1S21S58P066P009P002P037(0) <='1';
          else
          cVar1S21S58P066P009P002P037(0) <='0';
          end if;
        if(D( 8)='1' AND A(15)='1' AND A(28)='0' AND B(10)='0' )then
          cVar1S22S58P066P009P002N037(0) <='1';
          else
          cVar1S22S58P066P009P002N037(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='0' AND D(16)='1' )then
          cVar1S0S59P018P008P050P067(0) <='1';
          else
          cVar1S0S59P018P008P050P067(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='0' AND D(16)='1' )then
          cVar1S1S59P018P008P050P067(0) <='1';
          else
          cVar1S1S59P018P008P050P067(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='0' AND D(16)='1' )then
          cVar1S2S59P018P008P050P067(0) <='1';
          else
          cVar1S2S59P018P008P050P067(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='0' AND D(16)='0' )then
          cVar1S3S59P018P008P050N067(0) <='1';
          else
          cVar1S3S59P018P008P050N067(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='0' AND D(16)='0' )then
          cVar1S4S59P018P008P050N067(0) <='1';
          else
          cVar1S4S59P018P008P050N067(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='1' AND A(15)='1' )then
          cVar1S5S59P018P008P050P009(0) <='1';
          else
          cVar1S5S59P018P008P050P009(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND D(12)='1' AND A(15)='0' )then
          cVar1S6S59P018P008P050N009(0) <='1';
          else
          cVar1S6S59P018P008P050N009(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND A(12)='0' )then
          cVar1S7S59P018P008P054P015(0) <='1';
          else
          cVar1S7S59P018P008P054P015(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND A(12)='0' )then
          cVar1S8S59P018P008P054P015(0) <='1';
          else
          cVar1S8S59P018P008P054P015(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND A(12)='1' )then
          cVar1S9S59P018P008P054P015(0) <='1';
          else
          cVar1S9S59P018P008P054P015(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND A(12)='1' )then
          cVar1S10S59P018P008P054P015(0) <='1';
          else
          cVar1S10S59P018P008P054P015(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='1' AND B(25)='1' )then
          cVar1S11S59N018P061P008P026(0) <='1';
          else
          cVar1S11S59N018P061P008P026(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='1' AND B(25)='0' )then
          cVar1S12S59N018P061P008N026(0) <='1';
          else
          cVar1S12S59N018P061P008N026(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='1' AND B(25)='0' )then
          cVar1S13S59N018P061P008N026(0) <='1';
          else
          cVar1S13S59N018P061P008N026(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='0' AND D(23)='1' )then
          cVar1S14S59N018P061N008P039(0) <='1';
          else
          cVar1S14S59N018P061N008P039(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='0' AND D(23)='1' )then
          cVar1S15S59N018P061N008P039(0) <='1';
          else
          cVar1S15S59N018P061N008P039(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='0' AND D(23)='0' )then
          cVar1S16S59N018P061N008N039(0) <='1';
          else
          cVar1S16S59N018P061N008N039(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND A(25)='0' AND D(23)='0' )then
          cVar1S17S59N018P061N008N039(0) <='1';
          else
          cVar1S17S59N018P061N008N039(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S18S59N018P061P059P000(0) <='1';
          else
          cVar1S18S59N018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='1' )then
          cVar1S19S59N018P061N059P063(0) <='1';
          else
          cVar1S19S59N018P061N059P063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='0' )then
          cVar1S20S59N018P061N059N063(0) <='1';
          else
          cVar1S20S59N018P061N059N063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='1' )then
          cVar1S0S60P018P061P067P010(0) <='1';
          else
          cVar1S0S60P018P061P067P010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='1' )then
          cVar1S1S60P018P061P067P010(0) <='1';
          else
          cVar1S1S60P018P061P067P010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='1' )then
          cVar1S2S60P018P061P067P010(0) <='1';
          else
          cVar1S2S60P018P061P067P010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='0' )then
          cVar1S3S60P018P061P067N010(0) <='1';
          else
          cVar1S3S60P018P061P067N010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='0' )then
          cVar1S4S60P018P061P067N010(0) <='1';
          else
          cVar1S4S60P018P061P067N010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='0' AND A(24)='0' )then
          cVar1S5S60P018P061P067N010(0) <='1';
          else
          cVar1S5S60P018P061P067N010(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='1' AND A(13)='0' )then
          cVar1S6S60P018P061P067P013(0) <='1';
          else
          cVar1S6S60P018P061P067P013(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(16)='1' AND A(13)='1' )then
          cVar1S7S60P018P061P067P013(0) <='1';
          else
          cVar1S7S60P018P061P067P013(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S8S60P018P061P059P000(0) <='1';
          else
          cVar1S8S60P018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='1' )then
          cVar1S9S60P018P061N059P063(0) <='1';
          else
          cVar1S9S60P018P061N059P063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='1' )then
          cVar1S10S60P018P061N059P063(0) <='1';
          else
          cVar1S10S60P018P061N059P063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='0' )then
          cVar1S11S60P018P061N059N063(0) <='1';
          else
          cVar1S11S60P018P061N059N063(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='0' AND E(11)='1' )then
          cVar1S12S60P018P067P019P056nsss(0) <='1';
          else
          cVar1S12S60P018P067P019P056nsss(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='0' AND E(11)='0' )then
          cVar1S13S60P018P067P019N056(0) <='1';
          else
          cVar1S13S60P018P067P019N056(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='0' AND E(11)='0' )then
          cVar1S14S60P018P067P019N056(0) <='1';
          else
          cVar1S14S60P018P067P019N056(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='0' AND E(11)='0' )then
          cVar1S15S60P018P067P019N056(0) <='1';
          else
          cVar1S15S60P018P067P019N056(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='1' AND B(26)='0' )then
          cVar1S16S60P018P067P019P024(0) <='1';
          else
          cVar1S16S60P018P067P019P024(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='1' AND B(26)='0' )then
          cVar1S17S60P018P067P019P024(0) <='1';
          else
          cVar1S17S60P018P067P019P024(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='1' AND A(10)='1' AND B(26)='0' )then
          cVar1S18S60P018P067P019P024(0) <='1';
          else
          cVar1S18S60P018P067P019P024(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='0' AND E(16)='0' AND B(23)='0' )then
          cVar1S19S60P018N067P069P030(0) <='1';
          else
          cVar1S19S60P018N067P069P030(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='0' AND E(16)='0' AND B(23)='0' )then
          cVar1S20S60P018N067P069P030(0) <='1';
          else
          cVar1S20S60P018N067P069P030(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='0' AND E(16)='0' AND B(23)='1' )then
          cVar1S21S60P018N067P069P030(0) <='1';
          else
          cVar1S21S60P018N067P069P030(0) <='0';
          end if;
        if(A(20)='1' AND D(16)='0' AND E(16)='1' AND A(22)='0' )then
          cVar1S22S60P018N067P069P014(0) <='1';
          else
          cVar1S22S60P018N067P069P014(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='0' AND B(21)='0' )then
          cVar1S0S61P018P008P024P034(0) <='1';
          else
          cVar1S0S61P018P008P024P034(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='0' AND B(21)='0' )then
          cVar1S1S61P018P008P024P034(0) <='1';
          else
          cVar1S1S61P018P008P024P034(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='0' AND B(21)='0' )then
          cVar1S2S61P018P008P024P034(0) <='1';
          else
          cVar1S2S61P018P008P024P034(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='0' AND B(21)='0' )then
          cVar1S3S61P018P008P024P034(0) <='1';
          else
          cVar1S3S61P018P008P024P034(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='0' AND B(21)='1' )then
          cVar1S4S61P018P008P024P034(0) <='1';
          else
          cVar1S4S61P018P008P024P034(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='1' AND E(22)='1' )then
          cVar1S5S61P018P008P024P045nsss(0) <='1';
          else
          cVar1S5S61P018P008P024P045nsss(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='1' AND E(22)='0' )then
          cVar1S6S61P018P008P024N045(0) <='1';
          else
          cVar1S6S61P018P008P024N045(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='0' AND B(26)='1' AND E(22)='0' )then
          cVar1S7S61P018P008P024N045(0) <='1';
          else
          cVar1S7S61P018P008P024N045(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND B(27)='0' )then
          cVar1S8S61P018P008P054P022(0) <='1';
          else
          cVar1S8S61P018P008P054P022(0) <='0';
          end if;
        if(A(20)='1' AND A(25)='1' AND D(11)='0' AND B(27)='0' )then
          cVar1S9S61P018P008P054P022(0) <='1';
          else
          cVar1S9S61P018P008P054P022(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='1' AND B(12)='0' )then
          cVar1S10S61N018P061P050P033(0) <='1';
          else
          cVar1S10S61N018P061P050P033(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='1' AND B(12)='0' )then
          cVar1S11S61N018P061P050P033(0) <='1';
          else
          cVar1S11S61N018P061P050P033(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='0' AND A(27)='1' )then
          cVar1S12S61N018P061N050P004(0) <='1';
          else
          cVar1S12S61N018P061N050P004(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='0' AND A(27)='1' )then
          cVar1S13S61N018P061N050P004(0) <='1';
          else
          cVar1S13S61N018P061N050P004(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='0' AND A(27)='1' )then
          cVar1S14S61N018P061N050P004(0) <='1';
          else
          cVar1S14S61N018P061N050P004(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='0' AND A(27)='0' )then
          cVar1S15S61N018P061N050N004(0) <='1';
          else
          cVar1S15S61N018P061N050N004(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(12)='0' AND A(27)='0' )then
          cVar1S16S61N018P061N050N004(0) <='1';
          else
          cVar1S16S61N018P061N050N004(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S17S61N018P061P059P000(0) <='1';
          else
          cVar1S17S61N018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S18S61N018P061P059P000(0) <='1';
          else
          cVar1S18S61N018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='1' )then
          cVar1S19S61N018P061N059P063(0) <='1';
          else
          cVar1S19S61N018P061N059P063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='0' )then
          cVar1S20S61N018P061N059N063(0) <='1';
          else
          cVar1S20S61N018P061N059N063(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='0' AND B(24)='1' )then
          cVar1S0S62P000P018P061P028(0) <='1';
          else
          cVar1S0S62P000P018P061P028(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='0' AND B(24)='1' )then
          cVar1S1S62P000P018P061P028(0) <='1';
          else
          cVar1S1S62P000P018P061P028(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='0' AND B(24)='0' )then
          cVar1S2S62P000P018P061N028(0) <='1';
          else
          cVar1S2S62P000P018P061N028(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='0' AND B(24)='0' )then
          cVar1S3S62P000P018P061N028(0) <='1';
          else
          cVar1S3S62P000P018P061N028(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='0' AND B(24)='0' )then
          cVar1S4S62P000P018P061N028(0) <='1';
          else
          cVar1S4S62P000P018P061N028(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='1' AND D(18)='1' )then
          cVar1S5S62P000P018P061P059(0) <='1';
          else
          cVar1S5S62P000P018P061P059(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='1' AND D(18)='0' )then
          cVar1S6S62P000P018P061N059(0) <='1';
          else
          cVar1S6S62P000P018P061N059(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND E(18)='1' AND D(18)='0' )then
          cVar1S7S62P000P018P061N059(0) <='1';
          else
          cVar1S7S62P000P018P061N059(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND D(22)='0' AND B(26)='0' )then
          cVar1S8S62P000P018P043P024(0) <='1';
          else
          cVar1S8S62P000P018P043P024(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND D(22)='0' AND B(26)='0' )then
          cVar1S9S62P000P018P043P024(0) <='1';
          else
          cVar1S9S62P000P018P043P024(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND D(22)='0' AND B(26)='0' )then
          cVar1S10S62P000P018P043P024(0) <='1';
          else
          cVar1S10S62P000P018P043P024(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND D(22)='1' AND E(22)='1' )then
          cVar1S11S62P000P018P043P045(0) <='1';
          else
          cVar1S11S62P000P018P043P045(0) <='0';
          end if;
        if(A(29)='1' AND B(23)='0' AND B(15)='0' AND E(11)='0' )then
          cVar1S12S62P000P030P027P056(0) <='1';
          else
          cVar1S12S62P000P030P027P056(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='1' AND A(24)='1' )then
          cVar1S0S63P000P018P028P010(0) <='1';
          else
          cVar1S0S63P000P018P028P010(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='1' AND A(24)='0' )then
          cVar1S1S63P000P018P028N010(0) <='1';
          else
          cVar1S1S63P000P018P028N010(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='1' )then
          cVar1S2S63P000P018N028P030(0) <='1';
          else
          cVar1S2S63P000P018N028P030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='1' )then
          cVar1S3S63P000P018N028P030(0) <='1';
          else
          cVar1S3S63P000P018N028P030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='1' )then
          cVar1S4S63P000P018N028P030(0) <='1';
          else
          cVar1S4S63P000P018N028P030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='1' )then
          cVar1S5S63P000P018N028P030(0) <='1';
          else
          cVar1S5S63P000P018N028P030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='0' )then
          cVar1S6S63P000P018N028N030(0) <='1';
          else
          cVar1S6S63P000P018N028N030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='0' )then
          cVar1S7S63P000P018N028N030(0) <='1';
          else
          cVar1S7S63P000P018N028N030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='0' AND B(24)='0' AND B(23)='0' )then
          cVar1S8S63P000P018N028N030(0) <='1';
          else
          cVar1S8S63P000P018N028N030(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='1' AND A(27)='0' )then
          cVar1S9S63P000P018P036P004(0) <='1';
          else
          cVar1S9S63P000P018P036P004(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='1' AND A(27)='0' )then
          cVar1S10S63P000P018P036P004(0) <='1';
          else
          cVar1S10S63P000P018P036P004(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='1' AND A(27)='0' )then
          cVar1S11S63P000P018P036P004(0) <='1';
          else
          cVar1S11S63P000P018P036P004(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='1' AND A(27)='1' )then
          cVar1S12S63P000P018P036P004(0) <='1';
          else
          cVar1S12S63P000P018P036P004(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='0' AND E(19)='0' )then
          cVar1S13S63P000P018N036P057(0) <='1';
          else
          cVar1S13S63P000P018N036P057(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='0' AND E(19)='0' )then
          cVar1S14S63P000P018N036P057(0) <='1';
          else
          cVar1S14S63P000P018N036P057(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='0' AND E(19)='1' )then
          cVar1S15S63P000P018N036P057(0) <='1';
          else
          cVar1S15S63P000P018N036P057(0) <='0';
          end if;
        if(A(29)='0' AND A(20)='1' AND B(20)='0' AND E(19)='1' )then
          cVar1S16S63P000P018N036P057(0) <='1';
          else
          cVar1S16S63P000P018N036P057(0) <='0';
          end if;
        if(A(29)='1' AND B(23)='0' AND B(15)='0' AND B(28)='0' )then
          cVar1S17S63P000P030P027P020(0) <='1';
          else
          cVar1S17S63P000P030P027P020(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='1' )then
          cVar1S0S64P018P061P059P028(0) <='1';
          else
          cVar1S0S64P018P061P059P028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='1' )then
          cVar1S1S64P018P061P059P028(0) <='1';
          else
          cVar1S1S64P018P061P059P028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='0' )then
          cVar1S2S64P018P061P059N028(0) <='1';
          else
          cVar1S2S64P018P061P059N028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='0' )then
          cVar1S3S64P018P061P059N028(0) <='1';
          else
          cVar1S3S64P018P061P059N028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='0' )then
          cVar1S4S64P018P061P059N028(0) <='1';
          else
          cVar1S4S64P018P061P059N028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='0' AND B(24)='0' )then
          cVar1S5S64P018P061P059N028(0) <='1';
          else
          cVar1S5S64P018P061P059N028(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='0' AND D(18)='1' AND A(23)='1' )then
          cVar1S6S64P018P061P059P012(0) <='1';
          else
          cVar1S6S64P018P061P059P012(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S7S64P018P061P059P000(0) <='1';
          else
          cVar1S7S64P018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S8S64P018P061P059P000(0) <='1';
          else
          cVar1S8S64P018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='1' AND A(29)='0' )then
          cVar1S9S64P018P061P059P000(0) <='1';
          else
          cVar1S9S64P018P061P059P000(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='1' )then
          cVar1S10S64P018P061N059P063(0) <='1';
          else
          cVar1S10S64P018P061N059P063(0) <='0';
          end if;
        if(A(20)='0' AND E(18)='1' AND D(18)='0' AND D(17)='0' )then
          cVar1S11S64P018P061N059N063(0) <='1';
          else
          cVar1S11S64P018P061N059N063(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='0' )then
          cVar1S12S64P018P034P039P050(0) <='1';
          else
          cVar1S12S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='0' )then
          cVar1S13S64P018P034P039P050(0) <='1';
          else
          cVar1S13S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='0' )then
          cVar1S14S64P018P034P039P050(0) <='1';
          else
          cVar1S14S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='0' )then
          cVar1S15S64P018P034P039P050(0) <='1';
          else
          cVar1S15S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='1' )then
          cVar1S16S64P018P034P039P050(0) <='1';
          else
          cVar1S16S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='1' )then
          cVar1S17S64P018P034P039P050(0) <='1';
          else
          cVar1S17S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='0' AND D(12)='1' )then
          cVar1S18S64P018P034P039P050(0) <='1';
          else
          cVar1S18S64P018P034P039P050(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(23)='1' AND E( 8)='1' )then
          cVar1S19S64P018P034P039P068nsss(0) <='1';
          else
          cVar1S19S64P018P034P039P068nsss(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='1' AND D(21)='0' AND E(16)='0' )then
          cVar1S20S64P018P034P047P069(0) <='1';
          else
          cVar1S20S64P018P034P047P069(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='1' AND D(21)='0' AND E(16)='0' )then
          cVar1S21S64P018P034P047P069(0) <='1';
          else
          cVar1S21S64P018P034P047P069(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='1' AND D(21)='0' AND E(16)='1' )then
          cVar1S22S64P018P034P047P069(0) <='1';
          else
          cVar1S22S64P018P034P047P069(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='0' AND D(23)='0' )then
          cVar1S0S65P018P034P050P039(0) <='1';
          else
          cVar1S0S65P018P034P050P039(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='0' AND D(23)='0' )then
          cVar1S1S65P018P034P050P039(0) <='1';
          else
          cVar1S1S65P018P034P050P039(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='0' AND D(23)='0' )then
          cVar1S2S65P018P034P050P039(0) <='1';
          else
          cVar1S2S65P018P034P050P039(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='0' AND D(23)='1' )then
          cVar1S3S65P018P034P050P039(0) <='1';
          else
          cVar1S3S65P018P034P050P039(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='0' AND D(23)='1' )then
          cVar1S4S65P018P034P050P039(0) <='1';
          else
          cVar1S4S65P018P034P050P039(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='1' AND E(13)='1' )then
          cVar1S5S65P018P034P050P048(0) <='1';
          else
          cVar1S5S65P018P034P050P048(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='1' AND E(13)='0' )then
          cVar1S6S65P018P034P050N048(0) <='1';
          else
          cVar1S6S65P018P034P050N048(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='0' AND D(12)='1' AND E(13)='0' )then
          cVar1S7S65P018P034P050N048(0) <='1';
          else
          cVar1S7S65P018P034P050N048(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='1' AND D(21)='0' AND E(16)='0' )then
          cVar1S8S65P018P034P047P069(0) <='1';
          else
          cVar1S8S65P018P034P047P069(0) <='0';
          end if;
        if(A(20)='1' AND B(21)='1' AND D(21)='0' AND E(16)='1' )then
          cVar1S9S65P018P034P047P069(0) <='1';
          else
          cVar1S9S65P018P034P047P069(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='1' AND B(23)='0' AND A(24)='1' )then
          cVar1S10S65N018P028P030P010(0) <='1';
          else
          cVar1S10S65N018P028P030P010(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='1' AND B(23)='0' AND A(24)='1' )then
          cVar1S11S65N018P028P030P010(0) <='1';
          else
          cVar1S11S65N018P028P030P010(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='1' AND B(23)='0' AND A(24)='1' )then
          cVar1S12S65N018P028P030P010(0) <='1';
          else
          cVar1S12S65N018P028P030P010(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='1' AND B(23)='0' AND A(24)='0' )then
          cVar1S13S65N018P028P030N010(0) <='1';
          else
          cVar1S13S65N018P028P030N010(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S14S65N018N028P041P039(0) <='1';
          else
          cVar1S14S65N018N028P041P039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='1' AND D(23)='1' )then
          cVar1S15S65N018N028P041P039(0) <='1';
          else
          cVar1S15S65N018N028P041P039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='1' AND D(23)='0' )then
          cVar1S16S65N018N028P041N039(0) <='1';
          else
          cVar1S16S65N018N028P041N039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S17S65N018N028N041P039(0) <='1';
          else
          cVar1S17S65N018N028N041P039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S18S65N018N028N041P039(0) <='1';
          else
          cVar1S18S65N018N028N041P039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='0' AND D(23)='0' )then
          cVar1S19S65N018N028N041P039(0) <='1';
          else
          cVar1S19S65N018N028N041P039(0) <='0';
          end if;
        if(A(20)='0' AND B(24)='0' AND E(23)='0' AND D(23)='1' )then
          cVar1S20S65N018N028N041P039(0) <='1';
          else
          cVar1S20S65N018N028N041P039(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='1' AND E(15)='1' )then
          cVar1S0S66P016P000P002P040nsss(0) <='1';
          else
          cVar1S0S66P016P000P002P040nsss(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='1' AND E(15)='0' )then
          cVar1S1S66P016P000P002N040(0) <='1';
          else
          cVar1S1S66P016P000P002N040(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='1' AND E(15)='0' )then
          cVar1S2S66P016P000P002N040(0) <='1';
          else
          cVar1S2S66P016P000P002N040(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='0' AND B(21)='0' )then
          cVar1S3S66P016P000N002P034(0) <='1';
          else
          cVar1S3S66P016P000N002P034(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='0' AND B(21)='0' )then
          cVar1S4S66P016P000N002P034(0) <='1';
          else
          cVar1S4S66P016P000N002P034(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='0' AND B(21)='0' )then
          cVar1S5S66P016P000N002P034(0) <='1';
          else
          cVar1S5S66P016P000N002P034(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='0' AND A(28)='0' AND B(21)='1' )then
          cVar1S6S66P016P000N002P034(0) <='1';
          else
          cVar1S6S66P016P000N002P034(0) <='0';
          end if;
        if(A(21)='0' AND A(29)='1' AND E(20)='0' AND B(13)='0' )then
          cVar1S7S66P016P000P053P031(0) <='1';
          else
          cVar1S7S66P016P000P053P031(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='0' )then
          cVar1S8S66P016P039P022P041(0) <='1';
          else
          cVar1S8S66P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='1' )then
          cVar1S9S66P016P039P022P041(0) <='1';
          else
          cVar1S9S66P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='1' AND A(10)='1' )then
          cVar1S10S66P016P039P022P019(0) <='1';
          else
          cVar1S10S66P016P039P022P019(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(16)='0' AND A(17)='1' )then
          cVar1S11S66P016P039P007P005nsss(0) <='1';
          else
          cVar1S11S66P016P039P007P005nsss(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(16)='0' AND A(17)='0' )then
          cVar1S12S66P016P039P007N005(0) <='1';
          else
          cVar1S12S66P016P039P007N005(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND B(15)='0' AND E(14)='0' )then
          cVar1S0S67P014P024P027P044(0) <='1';
          else
          cVar1S0S67P014P024P027P044(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND B(15)='0' AND E(14)='0' )then
          cVar1S1S67P014P024P027P044(0) <='1';
          else
          cVar1S1S67P014P024P027P044(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND B(15)='0' AND E(14)='0' )then
          cVar1S2S67P014P024P027P044(0) <='1';
          else
          cVar1S2S67P014P024P027P044(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND B(15)='0' AND E(14)='1' )then
          cVar1S3S67P014P024P027P044(0) <='1';
          else
          cVar1S3S67P014P024P027P044(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S4S67P014P024P027P009nsss(0) <='1';
          else
          cVar1S4S67P014P024P027P009nsss(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND D(22)='1' )then
          cVar1S5S67P014P024P031P043nsss(0) <='1';
          else
          cVar1S5S67P014P024P031P043nsss(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(15)='1' AND D(12)='1' )then
          cVar1S6S67N014P027P009P050nsss(0) <='1';
          else
          cVar1S6S67N014P027P009P050nsss(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(15)='1' AND D(12)='0' )then
          cVar1S7S67N014P027P009N050(0) <='1';
          else
          cVar1S7S67N014P027P009N050(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(15)='0' AND A(29)='0' )then
          cVar1S8S67N014P027N009P000(0) <='1';
          else
          cVar1S8S67N014P027N009P000(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='0' AND B(26)='1' )then
          cVar1S9S67N014N027P050P024(0) <='1';
          else
          cVar1S9S67N014N027P050P024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='0' AND B(26)='1' )then
          cVar1S10S67N014N027P050P024(0) <='1';
          else
          cVar1S10S67N014N027P050P024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='0' AND B(26)='0' )then
          cVar1S11S67N014N027P050N024(0) <='1';
          else
          cVar1S11S67N014N027P050N024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='0' AND B(26)='0' )then
          cVar1S12S67N014N027P050N024(0) <='1';
          else
          cVar1S12S67N014N027P050N024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='1' AND B(22)='0' )then
          cVar1S13S67N014N027P050P032(0) <='1';
          else
          cVar1S13S67N014N027P050P032(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='1' AND B(22)='0' )then
          cVar1S14S67N014N027P050P032(0) <='1';
          else
          cVar1S14S67N014N027P050P032(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND D(12)='1' AND B(22)='0' )then
          cVar1S15S67N014N027P050P032(0) <='1';
          else
          cVar1S15S67N014N027P050P032(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='0' AND B(25)='0' )then
          cVar1S0S68P006P024P049P026(0) <='1';
          else
          cVar1S0S68P006P024P049P026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='0' AND B(25)='0' )then
          cVar1S1S68P006P024P049P026(0) <='1';
          else
          cVar1S1S68P006P024P049P026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='0' AND B(25)='0' )then
          cVar1S2S68P006P024P049P026(0) <='1';
          else
          cVar1S2S68P006P024P049P026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='0' AND B(25)='1' )then
          cVar1S3S68P006P024P049P026(0) <='1';
          else
          cVar1S3S68P006P024P049P026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='1' AND B(25)='1' )then
          cVar1S4S68P006P024P049P026nsss(0) <='1';
          else
          cVar1S4S68P006P024P049P026nsss(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='1' AND B(25)='0' )then
          cVar1S5S68P006P024P049N026(0) <='1';
          else
          cVar1S5S68P006P024P049N026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='0' AND E(21)='1' AND B(25)='0' )then
          cVar1S6S68P006P024P049N026(0) <='1';
          else
          cVar1S6S68P006P024P049N026(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(24)='0' AND D(21)='1' )then
          cVar1S7S68P006P024P010P047nsss(0) <='1';
          else
          cVar1S7S68P006P024P010P047nsss(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(24)='0' AND D(21)='0' )then
          cVar1S8S68P006P024P010N047(0) <='1';
          else
          cVar1S8S68P006P024P010N047(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(24)='0' AND D(21)='0' )then
          cVar1S9S68P006P024P010N047(0) <='1';
          else
          cVar1S9S68P006P024P010N047(0) <='0';
          end if;
        if(A(26)='0' AND B(26)='1' AND A(24)='1' AND A(10)='0' )then
          cVar1S10S68P006P024P010P019(0) <='1';
          else
          cVar1S10S68P006P024P010P019(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='1' AND A(28)='0' AND A(14)='0' )then
          cVar1S11S68P006P024P002P011(0) <='1';
          else
          cVar1S11S68P006P024P002P011(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='1' AND A(28)='0' AND A(14)='0' )then
          cVar1S12S68P006P024P002P011(0) <='1';
          else
          cVar1S12S68P006P024P002P011(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='0' AND E(17)='0' AND B(21)='0' )then
          cVar1S13S68P006N024P065P034(0) <='1';
          else
          cVar1S13S68P006N024P065P034(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='0' AND E(17)='0' AND B(21)='0' )then
          cVar1S14S68P006N024P065P034(0) <='1';
          else
          cVar1S14S68P006N024P065P034(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='0' AND E(17)='0' AND B(21)='1' )then
          cVar1S15S68P006N024P065P034(0) <='1';
          else
          cVar1S15S68P006N024P065P034(0) <='0';
          end if;
        if(A(26)='1' AND B(26)='0' AND E(17)='1' AND A(13)='0' )then
          cVar1S16S68P006N024P065P013(0) <='1';
          else
          cVar1S16S68P006N024P065P013(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='1' AND E(19)='1' )then
          cVar1S0S69P055P026P010P057(0) <='1';
          else
          cVar1S0S69P055P026P010P057(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='1' AND E(19)='1' )then
          cVar1S1S69P055P026P010P057(0) <='1';
          else
          cVar1S1S69P055P026P010P057(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='1' AND E(19)='0' )then
          cVar1S2S69P055P026P010N057(0) <='1';
          else
          cVar1S2S69P055P026P010N057(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='0' AND E(17)='1' )then
          cVar1S3S69P055P026N010P065nsss(0) <='1';
          else
          cVar1S3S69P055P026N010P065nsss(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='0' AND E(17)='0' )then
          cVar1S4S69P055P026N010N065(0) <='1';
          else
          cVar1S4S69P055P026N010N065(0) <='0';
          end if;
        if(D(19)='1' AND B(25)='0' AND A(24)='0' AND E(17)='0' )then
          cVar1S5S69P055P026N010N065(0) <='1';
          else
          cVar1S5S69P055P026N010N065(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='0' AND B(25)='1' AND A(27)='0' )then
          cVar1S6S69N055P030P026P004(0) <='1';
          else
          cVar1S6S69N055P030P026P004(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='0' AND B(25)='1' AND A(27)='0' )then
          cVar1S7S69N055P030P026P004(0) <='1';
          else
          cVar1S7S69N055P030P026P004(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='0' AND B(25)='0' AND E(19)='0' )then
          cVar1S8S69N055P030N026P057(0) <='1';
          else
          cVar1S8S69N055P030N026P057(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='0' AND B(25)='0' AND E(19)='0' )then
          cVar1S9S69N055P030N026P057(0) <='1';
          else
          cVar1S9S69N055P030N026P057(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='1' AND D(17)='0' AND A(28)='1' )then
          cVar1S10S69N055P030P063P002nsss(0) <='1';
          else
          cVar1S10S69N055P030P063P002nsss(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='1' AND D(17)='0' AND A(28)='0' )then
          cVar1S11S69N055P030P063N002(0) <='1';
          else
          cVar1S11S69N055P030P063N002(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='1' AND D(17)='0' AND A(28)='0' )then
          cVar1S12S69N055P030P063N002(0) <='1';
          else
          cVar1S12S69N055P030P063N002(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='1' AND D(17)='0' AND A(28)='0' )then
          cVar1S13S69N055P030P063N002(0) <='1';
          else
          cVar1S13S69N055P030P063N002(0) <='0';
          end if;
        if(D(19)='0' AND B(23)='1' AND D(17)='1' AND A(22)='0' )then
          cVar1S14S69N055P030P063P014(0) <='1';
          else
          cVar1S14S69N055P030P063P014(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='0' )then
          cVar1S0S70P050P027P048P025(0) <='1';
          else
          cVar1S0S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='0' )then
          cVar1S1S70P050P027P048P025(0) <='1';
          else
          cVar1S1S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='0' )then
          cVar1S2S70P050P027P048P025(0) <='1';
          else
          cVar1S2S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='1' )then
          cVar1S3S70P050P027P048P025(0) <='1';
          else
          cVar1S3S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='1' )then
          cVar1S4S70P050P027P048P025(0) <='1';
          else
          cVar1S4S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='0' AND B(16)='1' )then
          cVar1S5S70P050P027P048P025(0) <='1';
          else
          cVar1S5S70P050P027P048P025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='1' AND B(16)='1' )then
          cVar1S6S70P050P027P048P025nsss(0) <='1';
          else
          cVar1S6S70P050P027P048P025nsss(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='1' AND B(16)='0' )then
          cVar1S7S70P050P027P048N025(0) <='1';
          else
          cVar1S7S70P050P027P048N025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='1' AND B(16)='0' )then
          cVar1S8S70P050P027P048N025(0) <='1';
          else
          cVar1S8S70P050P027P048N025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='0' AND E(13)='1' AND B(16)='0' )then
          cVar1S9S70P050P027P048N025(0) <='1';
          else
          cVar1S9S70P050P027P048N025(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='1' AND A(29)='0' AND B(11)='0' )then
          cVar1S10S70P050P027P000P035(0) <='1';
          else
          cVar1S10S70P050P027P000P035(0) <='0';
          end if;
        if(D(12)='0' AND B(15)='1' AND A(29)='0' AND B(11)='0' )then
          cVar1S11S70P050P027P000P035(0) <='1';
          else
          cVar1S11S70P050P027P000P035(0) <='0';
          end if;
        if(D(12)='1' AND D(22)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S12S70P050P043P027P009nsss(0) <='1';
          else
          cVar1S12S70P050P043P027P009nsss(0) <='0';
          end if;
        if(D(12)='1' AND D(22)='0' AND B(15)='1' AND A(15)='0' )then
          cVar1S13S70P050P043P027N009(0) <='1';
          else
          cVar1S13S70P050P043P027N009(0) <='0';
          end if;
        if(D(12)='1' AND D(22)='0' AND B(15)='0' AND B(28)='0' )then
          cVar1S14S70P050P043N027P020(0) <='1';
          else
          cVar1S14S70P050P043N027P020(0) <='0';
          end if;
        if(D(12)='1' AND D(22)='0' AND B(15)='0' AND B(28)='0' )then
          cVar1S15S70P050P043N027P020(0) <='1';
          else
          cVar1S15S70P050P043N027P020(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' )then
          cVar1S0S71P021P040nsss(0) <='1';
          else
          cVar1S0S71P021P040nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(13)='0' AND D(23)='1' )then
          cVar1S1S71P021N040P048P039nsss(0) <='1';
          else
          cVar1S1S71P021N040P048P039nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(13)='0' AND D(23)='0' )then
          cVar1S2S71P021N040P048N039(0) <='1';
          else
          cVar1S2S71P021N040P048N039(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='1' )then
          cVar1S3S71N021P038P040P057(0) <='1';
          else
          cVar1S3S71N021P038P040P057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='1' )then
          cVar1S4S71N021P038P040P057(0) <='1';
          else
          cVar1S4S71N021P038P040P057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='0' )then
          cVar1S5S71N021P038P040N057(0) <='1';
          else
          cVar1S5S71N021P038P040N057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='0' )then
          cVar1S6S71N021P038P040N057(0) <='1';
          else
          cVar1S6S71N021P038P040N057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='0' )then
          cVar1S7S71N021P038P040N057(0) <='1';
          else
          cVar1S7S71N021P038P040N057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S8S71N021P038P040P059(0) <='1';
          else
          cVar1S8S71N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S9S71N021P038P040P059(0) <='1';
          else
          cVar1S9S71N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S10S71N021P038P040P059(0) <='1';
          else
          cVar1S10S71N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(15)='1' AND A(12)='1' )then
          cVar1S11S71N021P038P040P015nsss(0) <='1';
          else
          cVar1S11S71N021P038P040P015nsss(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(15)='1' AND A(12)='0' )then
          cVar1S12S71N021P038P040N015(0) <='1';
          else
          cVar1S12S71N021P038P040N015(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(15)='0' AND A(24)='1' )then
          cVar1S13S71N021P038N040P010nsss(0) <='1';
          else
          cVar1S13S71N021P038N040P010nsss(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='1' AND D(15)='1' )then
          cVar1S0S72P016P021P038nsss(0) <='1';
          else
          cVar1S0S72P016P021P038nsss(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='1' AND D(15)='0' AND A(14)='0' )then
          cVar1S1S72P016P021N038P011(0) <='1';
          else
          cVar1S1S72P016P021N038P011(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='1' AND D(15)='0' AND A(14)='0' )then
          cVar1S2S72P016P021N038P011(0) <='1';
          else
          cVar1S2S72P016P021N038P011(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S3S72P016N021P040P038(0) <='1';
          else
          cVar1S3S72P016N021P040P038(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S4S72P016N021P040P038(0) <='1';
          else
          cVar1S4S72P016N021P040P038(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S5S72P016N021P040P038(0) <='1';
          else
          cVar1S5S72P016N021P040P038(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='0' AND D(15)='1' )then
          cVar1S6S72P016N021P040P038(0) <='1';
          else
          cVar1S6S72P016N021P040P038(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='1' AND A(28)='1' )then
          cVar1S7S72P016N021P040P002nsss(0) <='1';
          else
          cVar1S7S72P016N021P040P002nsss(0) <='0';
          end if;
        if(A(21)='0' AND B(18)='0' AND E(15)='1' AND A(28)='0' )then
          cVar1S8S72P016N021P040N002(0) <='1';
          else
          cVar1S8S72P016N021P040N002(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='0' )then
          cVar1S9S72P016P039P041P022(0) <='1';
          else
          cVar1S9S72P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='0' )then
          cVar1S10S72P016P039P041P022(0) <='1';
          else
          cVar1S10S72P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='1' )then
          cVar1S11S72P016P039P041P022(0) <='1';
          else
          cVar1S11S72P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='1' AND E(16)='0' )then
          cVar1S12S72P016P039P041P069(0) <='1';
          else
          cVar1S12S72P016P039P041P069(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND D(11)='0' AND A(17)='1' )then
          cVar1S13S72P016P039P054P005nsss(0) <='1';
          else
          cVar1S13S72P016P039P054P005nsss(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND D(11)='0' AND A(17)='0' )then
          cVar1S14S72P016P039P054N005(0) <='1';
          else
          cVar1S14S72P016P039P054N005(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' )then
          cVar1S0S73P021P040nsss(0) <='1';
          else
          cVar1S0S73P021P040nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(13)='0' AND E(11)='0' )then
          cVar1S1S73P021N040P048P056(0) <='1';
          else
          cVar1S1S73P021N040P048P056(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(13)='0' AND E(11)='0' )then
          cVar1S2S73P021N040P048P056(0) <='1';
          else
          cVar1S2S73P021N040P048P056(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='1' )then
          cVar1S3S73N021P038P040P057(0) <='1';
          else
          cVar1S3S73N021P038P040P057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='1' )then
          cVar1S4S73N021P038P040P057(0) <='1';
          else
          cVar1S4S73N021P038P040P057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='0' )then
          cVar1S5S73N021P038P040N057(0) <='1';
          else
          cVar1S5S73N021P038P040N057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND E(19)='0' )then
          cVar1S6S73N021P038P040N057(0) <='1';
          else
          cVar1S6S73N021P038P040N057(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S7S73N021P038P040P059(0) <='1';
          else
          cVar1S7S73N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S8S73N021P038P040P059(0) <='1';
          else
          cVar1S8S73N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S9S73N021P038P040P059(0) <='1';
          else
          cVar1S9S73N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND B(28)='1' )then
          cVar1S10S73N021P038P020nsss(0) <='1';
          else
          cVar1S10S73N021P038P020nsss(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND B(28)='0' AND D(17)='0' )then
          cVar1S11S73N021P038N020P063(0) <='1';
          else
          cVar1S11S73N021P038N020P063(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND B(28)='0' AND D(17)='0' )then
          cVar1S12S73N021P038N020P063(0) <='1';
          else
          cVar1S12S73N021P038N020P063(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(28)='0' AND A(15)='1' )then
          cVar1S0S74P014P027P002P009nsss(0) <='1';
          else
          cVar1S0S74P014P027P002P009nsss(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(28)='0' AND A(15)='0' )then
          cVar1S1S74P014P027P002N009(0) <='1';
          else
          cVar1S1S74P014P027P002N009(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='1' AND A(28)='0' AND A(15)='0' )then
          cVar1S2S74P014P027P002N009(0) <='1';
          else
          cVar1S2S74P014P027P002N009(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='1' AND B(24)='1' )then
          cVar1S3S74P014N027P010P028(0) <='1';
          else
          cVar1S3S74P014N027P010P028(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='1' AND B(24)='1' )then
          cVar1S4S74P014N027P010P028(0) <='1';
          else
          cVar1S4S74P014N027P010P028(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='1' AND B(24)='0' )then
          cVar1S5S74P014N027P010N028(0) <='1';
          else
          cVar1S5S74P014N027P010N028(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='1' AND B(24)='0' )then
          cVar1S6S74P014N027P010N028(0) <='1';
          else
          cVar1S6S74P014N027P010N028(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='1' )then
          cVar1S7S74P014N027N010P024(0) <='1';
          else
          cVar1S7S74P014N027N010P024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='1' )then
          cVar1S8S74P014N027N010P024(0) <='1';
          else
          cVar1S8S74P014N027N010P024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='0' )then
          cVar1S9S74P014N027N010N024(0) <='1';
          else
          cVar1S9S74P014N027N010N024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='0' )then
          cVar1S10S74P014N027N010N024(0) <='1';
          else
          cVar1S10S74P014N027N010N024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='0' )then
          cVar1S11S74P014N027N010N024(0) <='1';
          else
          cVar1S11S74P014N027N010N024(0) <='0';
          end if;
        if(A(22)='0' AND B(15)='0' AND A(24)='0' AND B(26)='0' )then
          cVar1S12S74P014N027N010N024(0) <='1';
          else
          cVar1S12S74P014N027N010N024(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(10)='1' )then
          cVar1S13S74P014P024P044P037(0) <='1';
          else
          cVar1S13S74P014P024P044P037(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(10)='0' )then
          cVar1S14S74P014P024P044N037(0) <='1';
          else
          cVar1S14S74P014P024P044N037(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(10)='0' )then
          cVar1S15S74P014P024P044N037(0) <='1';
          else
          cVar1S15S74P014P024P044N037(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(10)='0' )then
          cVar1S16S74P014P024P044N037(0) <='1';
          else
          cVar1S16S74P014P024P044N037(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='1' AND E(17)='0' )then
          cVar1S17S74P014P024P044P065(0) <='1';
          else
          cVar1S17S74P014P024P044P065(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='1' )then
          cVar1S18S74P014P024P031P045nsss(0) <='1';
          else
          cVar1S18S74P014P024P031P045nsss(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='0' )then
          cVar1S19S74P014P024P031N045(0) <='1';
          else
          cVar1S19S74P014P024P031N045(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='0' )then
          cVar1S20S74P014P024P031N045(0) <='1';
          else
          cVar1S20S74P014P024P031N045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='1' AND A(18)='0' )then
          cVar1S0S75P010P024P028P003(0) <='1';
          else
          cVar1S0S75P010P024P028P003(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='0' )then
          cVar1S1S75P010P024N028P045(0) <='1';
          else
          cVar1S1S75P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='0' )then
          cVar1S2S75P010P024N028P045(0) <='1';
          else
          cVar1S2S75P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='0' )then
          cVar1S3S75P010P024N028P045(0) <='1';
          else
          cVar1S3S75P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='1' )then
          cVar1S4S75P010P024N028P045(0) <='1';
          else
          cVar1S4S75P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S5S75P010P024P064P019(0) <='1';
          else
          cVar1S5S75P010P024P064P019(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S6S75P010P024P064P019(0) <='1';
          else
          cVar1S6S75P010P024P064P019(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='0' )then
          cVar1S7S75N010P014P024P056(0) <='1';
          else
          cVar1S7S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='0' )then
          cVar1S8S75N010P014P024P056(0) <='1';
          else
          cVar1S8S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='0' )then
          cVar1S9S75N010P014P024P056(0) <='1';
          else
          cVar1S9S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='0' )then
          cVar1S10S75N010P014P024P056(0) <='1';
          else
          cVar1S10S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='1' )then
          cVar1S11S75N010P014P024P056(0) <='1';
          else
          cVar1S11S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='0' AND E(11)='1' )then
          cVar1S12S75N010P014P024P056(0) <='1';
          else
          cVar1S12S75N010P014P024P056(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='1' AND B(26)='1' AND D(20)='0' )then
          cVar1S13S75N010P014P024P051(0) <='1';
          else
          cVar1S13S75N010P014P024P051(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='1' AND D(12)='1' )then
          cVar1S14S75N010N014P027P050nsss(0) <='1';
          else
          cVar1S14S75N010N014P027P050nsss(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S15S75N010N014P027N050(0) <='1';
          else
          cVar1S15S75N010N014P027N050(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S16S75N010N014P027N050(0) <='1';
          else
          cVar1S16S75N010N014P027N050(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S17S75N010N014P027N050(0) <='1';
          else
          cVar1S17S75N010N014P027N050(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='0' AND B(26)='1' )then
          cVar1S18S75N010N014N027P024(0) <='1';
          else
          cVar1S18S75N010N014N027P024(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='0' AND B(26)='1' )then
          cVar1S19S75N010N014N027P024(0) <='1';
          else
          cVar1S19S75N010N014N027P024(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S20S75N010N014N027N024(0) <='1';
          else
          cVar1S20S75N010N014N027N024(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S21S75N010N014N027N024(0) <='1';
          else
          cVar1S21S75N010N014N027N024(0) <='0';
          end if;
        if(A(24)='0' AND A(22)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S22S75N010N014N027N024(0) <='1';
          else
          cVar1S22S75N010N014N027N024(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='1' AND B(22)='0' AND B(18)='0' )then
          cVar1S0S76P014P010P032P021(0) <='1';
          else
          cVar1S0S76P014P010P032P021(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='1' AND B(22)='0' AND B(18)='0' )then
          cVar1S1S76P014P010P032P021(0) <='1';
          else
          cVar1S1S76P014P010P032P021(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='1' AND B(22)='1' AND A(11)='1' )then
          cVar1S2S76P014P010P032P017(0) <='1';
          else
          cVar1S2S76P014P010P032P017(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='1' AND D(12)='1' )then
          cVar1S3S76P014N010P027P050nsss(0) <='1';
          else
          cVar1S3S76P014N010P027P050nsss(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S4S76P014N010P027N050(0) <='1';
          else
          cVar1S4S76P014N010P027N050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='1' AND D(12)='0' )then
          cVar1S5S76P014N010P027N050(0) <='1';
          else
          cVar1S5S76P014N010P027N050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S6S76P014N010N027P050(0) <='1';
          else
          cVar1S6S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S7S76P014N010N027P050(0) <='1';
          else
          cVar1S7S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S8S76P014N010N027P050(0) <='1';
          else
          cVar1S8S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='0' )then
          cVar1S9S76P014N010N027P050(0) <='1';
          else
          cVar1S9S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='1' )then
          cVar1S10S76P014N010N027P050(0) <='1';
          else
          cVar1S10S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='0' AND A(24)='0' AND B(15)='0' AND D(12)='1' )then
          cVar1S11S76P014N010N027P050(0) <='1';
          else
          cVar1S11S76P014N010N027P050(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(15)='0' )then
          cVar1S12S76P014P024P044P027(0) <='1';
          else
          cVar1S12S76P014P024P044P027(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(15)='0' )then
          cVar1S13S76P014P024P044P027(0) <='1';
          else
          cVar1S13S76P014P024P044P027(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(15)='1' )then
          cVar1S14S76P014P024P044P027(0) <='1';
          else
          cVar1S14S76P014P024P044P027(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='0' AND B(15)='1' )then
          cVar1S15S76P014P024P044P027(0) <='1';
          else
          cVar1S15S76P014P024P044P027(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='0' AND E(14)='1' AND D( 9)='0' )then
          cVar1S16S76P014P024P044P062(0) <='1';
          else
          cVar1S16S76P014P024P044P062(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='1' )then
          cVar1S17S76P014P024P031P045nsss(0) <='1';
          else
          cVar1S17S76P014P024P031P045nsss(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='0' )then
          cVar1S18S76P014P024P031N045(0) <='1';
          else
          cVar1S18S76P014P024P031N045(0) <='0';
          end if;
        if(A(22)='1' AND B(26)='1' AND B(13)='0' AND E(22)='0' )then
          cVar1S19S76P014P024P031N045(0) <='1';
          else
          cVar1S19S76P014P024P031N045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='1' AND A(18)='0' )then
          cVar1S0S77P010P024P028P003(0) <='1';
          else
          cVar1S0S77P010P024P028P003(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='1' AND A(18)='0' )then
          cVar1S1S77P010P024P028P003(0) <='1';
          else
          cVar1S1S77P010P024P028P003(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='1' AND A(18)='0' )then
          cVar1S2S77P010P024P028P003(0) <='1';
          else
          cVar1S2S77P010P024P028P003(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='0' )then
          cVar1S3S77P010P024N028P045(0) <='1';
          else
          cVar1S3S77P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='0' )then
          cVar1S4S77P010P024N028P045(0) <='1';
          else
          cVar1S4S77P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='0' AND B(24)='0' AND E(22)='1' )then
          cVar1S5S77P010P024N028P045(0) <='1';
          else
          cVar1S5S77P010P024N028P045(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S6S77P010P024P064P019(0) <='1';
          else
          cVar1S6S77P010P024P064P019(0) <='0';
          end if;
        if(A(24)='1' AND B(26)='1' AND E( 9)='0' AND A(10)='0' )then
          cVar1S7S77P010P024P064P019(0) <='1';
          else
          cVar1S7S77P010P024P064P019(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='1' AND D(13)='1' )then
          cVar1S8S77N010P025P046nsss(0) <='1';
          else
          cVar1S8S77N010P025P046nsss(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='1' AND D(13)='0' AND A(16)='1' )then
          cVar1S9S77N010P025N046P007nsss(0) <='1';
          else
          cVar1S9S77N010P025N046P007nsss(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='1' AND D(13)='0' AND A(16)='0' )then
          cVar1S10S77N010P025N046N007(0) <='1';
          else
          cVar1S10S77N010P025N046N007(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='1' AND D(13)='0' AND A(16)='0' )then
          cVar1S11S77N010P025N046N007(0) <='1';
          else
          cVar1S11S77N010P025N046N007(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='0' AND A(28)='1' )then
          cVar1S12S77N010N025P046P002(0) <='1';
          else
          cVar1S12S77N010N025P046P002(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='0' AND A(28)='1' )then
          cVar1S13S77N010N025P046P002(0) <='1';
          else
          cVar1S13S77N010N025P046P002(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='0' AND A(28)='1' )then
          cVar1S14S77N010N025P046P002(0) <='1';
          else
          cVar1S14S77N010N025P046P002(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='0' AND A(28)='0' )then
          cVar1S15S77N010N025P046N002(0) <='1';
          else
          cVar1S15S77N010N025P046N002(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='1' AND D(21)='1' )then
          cVar1S16S77N010N025P046P047nsss(0) <='1';
          else
          cVar1S16S77N010N025P046P047nsss(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='1' AND D(21)='0' )then
          cVar1S17S77N010N025P046N047(0) <='1';
          else
          cVar1S17S77N010N025P046N047(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='1' AND D(21)='0' )then
          cVar1S18S77N010N025P046N047(0) <='1';
          else
          cVar1S18S77N010N025P046N047(0) <='0';
          end if;
        if(A(24)='0' AND B(16)='0' AND D(13)='1' AND D(21)='0' )then
          cVar1S19S77N010N025P046N047(0) <='1';
          else
          cVar1S19S77N010N025P046N047(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='0' AND D(12)='1' )then
          cVar1S0S78P039P041P020P050(0) <='1';
          else
          cVar1S0S78P039P041P020P050(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='0' AND D(12)='0' )then
          cVar1S1S78P039P041P020N050(0) <='1';
          else
          cVar1S1S78P039P041P020N050(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='0' AND D(12)='0' )then
          cVar1S2S78P039P041P020N050(0) <='1';
          else
          cVar1S2S78P039P041P020N050(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='0' AND D(12)='0' )then
          cVar1S3S78P039P041P020N050(0) <='1';
          else
          cVar1S3S78P039P041P020N050(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='1' AND E(15)='1' )then
          cVar1S4S78P039P041P020P040nsss(0) <='1';
          else
          cVar1S4S78P039P041P020P040nsss(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='1' AND E(15)='0' )then
          cVar1S5S78P039P041P020N040(0) <='1';
          else
          cVar1S5S78P039P041P020N040(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='0' AND B(28)='1' AND E(15)='0' )then
          cVar1S6S78P039P041P020N040(0) <='1';
          else
          cVar1S6S78P039P041P020N040(0) <='0';
          end if;
        if(D(23)='0' AND E(23)='1' AND B(12)='1' )then
          cVar1S7S78P039P041P033nsss(0) <='1';
          else
          cVar1S7S78P039P041P033nsss(0) <='0';
          end if;
        if(D(23)='1' AND B(28)='1' AND E(23)='1' )then
          cVar1S8S78P039P020P041nsss(0) <='1';
          else
          cVar1S8S78P039P020P041nsss(0) <='0';
          end if;
        if(D(23)='1' AND B(28)='0' AND A(23)='0' AND E(10)='0' )then
          cVar1S9S78P039N020P012P060(0) <='1';
          else
          cVar1S9S78P039N020P012P060(0) <='0';
          end if;
        if(D(23)='1' AND B(28)='0' AND A(23)='0' AND E(10)='0' )then
          cVar1S10S78P039N020P012P060(0) <='1';
          else
          cVar1S10S78P039N020P012P060(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='1' )then
          cVar1S0S79P021P040nsss(0) <='1';
          else
          cVar1S0S79P021P040nsss(0) <='0';
          end if;
        if(B(18)='1' AND E(15)='0' AND E(13)='0' AND E(10)='0' )then
          cVar1S1S79P021N040P048P060(0) <='1';
          else
          cVar1S1S79P021N040P048P060(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='1' )then
          cVar1S2S79N021P038P040P050(0) <='1';
          else
          cVar1S2S79N021P038P040P050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='1' )then
          cVar1S3S79N021P038P040P050(0) <='1';
          else
          cVar1S3S79N021P038P040P050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='0' )then
          cVar1S4S79N021P038P040N050(0) <='1';
          else
          cVar1S4S79N021P038P040N050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='0' )then
          cVar1S5S79N021P038P040N050(0) <='1';
          else
          cVar1S5S79N021P038P040N050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='0' )then
          cVar1S6S79N021P038P040N050(0) <='1';
          else
          cVar1S6S79N021P038P040N050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='0' AND D(12)='0' )then
          cVar1S7S79N021P038P040N050(0) <='1';
          else
          cVar1S7S79N021P038P040N050(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S8S79N021P038P040P059(0) <='1';
          else
          cVar1S8S79N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S9S79N021P038P040P059(0) <='1';
          else
          cVar1S9S79N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='0' AND E(15)='1' AND D(18)='0' )then
          cVar1S10S79N021P038P040P059(0) <='1';
          else
          cVar1S10S79N021P038P040P059(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(17)='0' AND B(28)='1' )then
          cVar1S11S79N021P038P065P020nsss(0) <='1';
          else
          cVar1S11S79N021P038P065P020nsss(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(17)='0' AND B(28)='0' )then
          cVar1S12S79N021P038P065N020(0) <='1';
          else
          cVar1S12S79N021P038P065N020(0) <='0';
          end if;
        if(B(18)='0' AND D(15)='1' AND E(17)='0' AND B(28)='0' )then
          cVar1S13S79N021P038P065N020(0) <='1';
          else
          cVar1S13S79N021P038P065N020(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='1' )then
          cVar1S0S80P037P048P025nsss(0) <='1';
          else
          cVar1S0S80P037P048P025nsss(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND B(15)='1' )then
          cVar1S1S80P037P048N025P027nsss(0) <='1';
          else
          cVar1S1S80P037P048N025P027nsss(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND B(15)='0' )then
          cVar1S2S80P037P048N025N027(0) <='1';
          else
          cVar1S2S80P037P048N025N027(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND B(15)='0' )then
          cVar1S3S80P037P048N025N027(0) <='1';
          else
          cVar1S3S80P037P048N025N027(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND B(15)='0' )then
          cVar1S4S80P037P048N025N027(0) <='1';
          else
          cVar1S4S80P037P048N025N027(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='0' )then
          cVar1S5S80P037N048P046P064(0) <='1';
          else
          cVar1S5S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='0' )then
          cVar1S6S80P037N048P046P064(0) <='1';
          else
          cVar1S6S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='0' )then
          cVar1S7S80P037N048P046P064(0) <='1';
          else
          cVar1S7S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='1' )then
          cVar1S8S80P037N048P046P064(0) <='1';
          else
          cVar1S8S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='1' )then
          cVar1S9S80P037N048P046P064(0) <='1';
          else
          cVar1S9S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND E( 9)='1' )then
          cVar1S10S80P037N048P046P064(0) <='1';
          else
          cVar1S10S80P037N048P046P064(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='1' AND A(18)='0' )then
          cVar1S11S80P037N048P046P003(0) <='1';
          else
          cVar1S11S80P037N048P046P003(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='1' AND A(18)='0' )then
          cVar1S12S80P037N048P046P003(0) <='1';
          else
          cVar1S12S80P037N048P046P003(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND E( 9)='1' )then
          cVar1S13S80P037P013P048P064(0) <='1';
          else
          cVar1S13S80P037P013P048P064(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND E( 9)='1' )then
          cVar1S14S80P037P013P048P064(0) <='1';
          else
          cVar1S14S80P037P013P048P064(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND E( 9)='0' )then
          cVar1S15S80P037P013P048N064(0) <='1';
          else
          cVar1S15S80P037P013P048N064(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND E( 9)='0' )then
          cVar1S16S80P037P013P048N064(0) <='1';
          else
          cVar1S16S80P037P013P048N064(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='1' AND B(11)='0' )then
          cVar1S17S80P037P013P048P035(0) <='1';
          else
          cVar1S17S80P037P013P048P035(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND A(12)='0' )then
          cVar1S18S80P037P013P018P015(0) <='1';
          else
          cVar1S18S80P037P013P018P015(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND A(12)='0' )then
          cVar1S19S80P037P013P018P015(0) <='1';
          else
          cVar1S19S80P037P013P018P015(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND A(12)='1' )then
          cVar1S20S80P037P013P018P015(0) <='1';
          else
          cVar1S20S80P037P013P018P015(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND A(12)='1' )then
          cVar1S21S80P037P013P018P015(0) <='1';
          else
          cVar1S21S80P037P013P018P015(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='0' AND B(13)='1' )then
          cVar1S22S80P037P013N018P031nsss(0) <='1';
          else
          cVar1S22S80P037P013N018P031nsss(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='0' AND B(13)='0' )then
          cVar1S23S80P037P013N018N031(0) <='1';
          else
          cVar1S23S80P037P013N018N031(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='0' AND B(13)='0' )then
          cVar1S24S80P037P013N018N031(0) <='1';
          else
          cVar1S24S80P037P013N018N031(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='1' AND E(20)='0' )then
          cVar1S0S81P019P017P055P053(0) <='1';
          else
          cVar1S0S81P019P017P055P053(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S1S81P019P017N055P057(0) <='1';
          else
          cVar1S1S81P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S2S81P019P017N055P057(0) <='1';
          else
          cVar1S2S81P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S3S81P019P017N055P057(0) <='1';
          else
          cVar1S3S81P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S4S81P019P017N055P057(0) <='1';
          else
          cVar1S4S81P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='1' )then
          cVar1S5S81P019P017N055P057(0) <='1';
          else
          cVar1S5S81P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='0' AND B(14)='0' )then
          cVar1S6S81P019P017P064P029(0) <='1';
          else
          cVar1S6S81P019P017P064P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='0' AND B(14)='0' )then
          cVar1S7S81P019P017P064P029(0) <='1';
          else
          cVar1S7S81P019P017P064P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='0' AND B(14)='0' )then
          cVar1S8S81P019P017P064P029(0) <='1';
          else
          cVar1S8S81P019P017P064P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='0' AND B(14)='1' )then
          cVar1S9S81P019P017P064P029(0) <='1';
          else
          cVar1S9S81P019P017P064P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='1' AND A(14)='1' )then
          cVar1S10S81P019P017P064P011(0) <='1';
          else
          cVar1S10S81P019P017P064P011(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='1' AND A(14)='1' )then
          cVar1S11S81P019P017P064P011(0) <='1';
          else
          cVar1S11S81P019P017P064P011(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E( 9)='1' AND A(14)='0' )then
          cVar1S12S81P019P017P064N011(0) <='1';
          else
          cVar1S12S81P019P017P064N011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='0' AND B(11)='0' )then
          cVar1S13S81N019P037P003P035(0) <='1';
          else
          cVar1S13S81N019P037P003P035(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='0' AND B(11)='0' )then
          cVar1S14S81N019P037P003P035(0) <='1';
          else
          cVar1S14S81N019P037P003P035(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='0' AND B(11)='0' )then
          cVar1S15S81N019P037P003P035(0) <='1';
          else
          cVar1S15S81N019P037P003P035(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='0' AND B(11)='1' )then
          cVar1S16S81N019P037P003P035(0) <='1';
          else
          cVar1S16S81N019P037P003P035(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='0' AND B(11)='1' )then
          cVar1S17S81N019P037P003P035(0) <='1';
          else
          cVar1S17S81N019P037P003P035(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='1' AND B(21)='1' )then
          cVar1S18S81N019P037P003P034nsss(0) <='1';
          else
          cVar1S18S81N019P037P003P034nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND A(18)='1' AND B(21)='0' )then
          cVar1S19S81N019P037P003N034(0) <='1';
          else
          cVar1S19S81N019P037P003N034(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='1' AND D( 9)='1' )then
          cVar1S20S81N019N037P048P062nsss(0) <='1';
          else
          cVar1S20S81N019N037P048P062nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='1' AND D( 9)='0' )then
          cVar1S21S81N019N037P048N062(0) <='1';
          else
          cVar1S21S81N019N037P048N062(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='1' AND D( 9)='0' )then
          cVar1S22S81N019N037P048N062(0) <='1';
          else
          cVar1S22S81N019N037P048N062(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='1' AND D( 9)='0' )then
          cVar1S23S81N019N037P048N062(0) <='1';
          else
          cVar1S23S81N019N037P048N062(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='1' )then
          cVar1S24S81N019N037N048P057(0) <='1';
          else
          cVar1S24S81N019N037N048P057(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='1' )then
          cVar1S25S81N019N037N048P057(0) <='1';
          else
          cVar1S25S81N019N037N048P057(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='1' )then
          cVar1S26S81N019N037N048P057(0) <='1';
          else
          cVar1S26S81N019N037N048P057(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='0' )then
          cVar1S27S81N019N037N048N057(0) <='1';
          else
          cVar1S27S81N019N037N048N057(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='0' )then
          cVar1S28S81N019N037N048N057(0) <='1';
          else
          cVar1S28S81N019N037N048N057(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(13)='0' AND E(19)='0' )then
          cVar1S29S81N019N037N048N057(0) <='1';
          else
          cVar1S29S81N019N037N048N057(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='1' AND B(18)='1' )then
          cVar1S0S82P019P030P040P021nsss(0) <='1';
          else
          cVar1S0S82P019P030P040P021nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='1' AND B(18)='0' )then
          cVar1S1S82P019P030P040N021(0) <='1';
          else
          cVar1S1S82P019P030P040N021(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='1' AND B(18)='0' )then
          cVar1S2S82P019P030P040N021(0) <='1';
          else
          cVar1S2S82P019P030P040N021(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S3S82P019P030N040P038(0) <='1';
          else
          cVar1S3S82P019P030N040P038(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S4S82P019P030N040P038(0) <='1';
          else
          cVar1S4S82P019P030N040P038(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S5S82P019P030N040P038(0) <='1';
          else
          cVar1S5S82P019P030N040P038(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='1' AND E(22)='0' AND E(11)='1' )then
          cVar1S6S82P019P030P045P056nsss(0) <='1';
          else
          cVar1S6S82P019P030P045P056nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='1' AND E(22)='0' AND E(11)='0' )then
          cVar1S7S82P019P030P045N056(0) <='1';
          else
          cVar1S7S82P019P030P045N056(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='1' AND E(22)='0' AND E(11)='0' )then
          cVar1S8S82P019P030P045N056(0) <='1';
          else
          cVar1S8S82P019P030P045N056(0) <='0';
          end if;
        if(A(10)='0' AND B(23)='1' AND E(22)='0' AND E(11)='0' )then
          cVar1S9S82P019P030P045N056(0) <='1';
          else
          cVar1S9S82P019P030P045N056(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='1' AND E(17)='1' )then
          cVar1S10S82P019P017P055P065nsss(0) <='1';
          else
          cVar1S10S82P019P017P055P065nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='1' AND E(17)='0' )then
          cVar1S11S82P019P017P055N065(0) <='1';
          else
          cVar1S11S82P019P017P055N065(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S12S82P019P017N055P057(0) <='1';
          else
          cVar1S12S82P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S13S82P019P017N055P057(0) <='1';
          else
          cVar1S13S82P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='0' )then
          cVar1S14S82P019P017N055P057(0) <='1';
          else
          cVar1S14S82P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND D(19)='0' AND E(19)='1' )then
          cVar1S15S82P019P017N055P057(0) <='1';
          else
          cVar1S15S82P019P017N055P057(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='0' AND B(14)='0' )then
          cVar1S16S82P019P017P053P029(0) <='1';
          else
          cVar1S16S82P019P017P053P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='0' AND B(14)='0' )then
          cVar1S17S82P019P017P053P029(0) <='1';
          else
          cVar1S17S82P019P017P053P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='1' AND B(10)='1' )then
          cVar1S18S82P019P017P053P037(0) <='1';
          else
          cVar1S18S82P019P017P053P037(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='1' AND B(10)='0' )then
          cVar1S19S82P019P017P053N037(0) <='1';
          else
          cVar1S19S82P019P017P053N037(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='1' )then
          cVar1S0S83P015P051P017P012(0) <='1';
          else
          cVar1S0S83P015P051P017P012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='1' )then
          cVar1S1S83P015P051P017P012(0) <='1';
          else
          cVar1S1S83P015P051P017P012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='0' )then
          cVar1S2S83P015P051P017N012(0) <='1';
          else
          cVar1S2S83P015P051P017N012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='0' )then
          cVar1S3S83P015P051P017N012(0) <='1';
          else
          cVar1S3S83P015P051P017N012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='0' )then
          cVar1S4S83P015P051P017N012(0) <='1';
          else
          cVar1S4S83P015P051P017N012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='0' AND A(23)='0' )then
          cVar1S5S83P015P051P017N012(0) <='1';
          else
          cVar1S5S83P015P051P017N012(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='1' AND E(18)='0' )then
          cVar1S6S83P015P051P017P061(0) <='1';
          else
          cVar1S6S83P015P051P017P061(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='1' AND E(18)='0' )then
          cVar1S7S83P015P051P017P061(0) <='1';
          else
          cVar1S7S83P015P051P017P061(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='0' AND A(11)='1' AND E(18)='1' )then
          cVar1S8S83P015P051P017P061(0) <='1';
          else
          cVar1S8S83P015P051P017P061(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='1' AND A(29)='0' )then
          cVar1S9S83P015P051P053P000(0) <='1';
          else
          cVar1S9S83P015P051P053P000(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='1' AND A(29)='0' )then
          cVar1S10S83P015P051P053P000(0) <='1';
          else
          cVar1S10S83P015P051P053P000(0) <='0';
          end if;
        if(A(12)='1' AND D(20)='1' AND E(20)='0' AND A(22)='0' )then
          cVar1S11S83P015P051N053P014(0) <='1';
          else
          cVar1S11S83P015P051N053P014(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='1' AND D(15)='1' )then
          cVar1S12S83N015P021P038nsss(0) <='1';
          else
          cVar1S12S83N015P021P038nsss(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='1' AND D(15)='0' AND E(16)='0' )then
          cVar1S13S83N015P021N038P069(0) <='1';
          else
          cVar1S13S83N015P021N038P069(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='1' AND D(15)='0' AND E(16)='0' )then
          cVar1S14S83N015P021N038P069(0) <='1';
          else
          cVar1S14S83N015P021N038P069(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='1' )then
          cVar1S15S83N015N021P038P067(0) <='1';
          else
          cVar1S15S83N015N021P038P067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='1' )then
          cVar1S16S83N015N021P038P067(0) <='1';
          else
          cVar1S16S83N015N021P038P067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='1' )then
          cVar1S17S83N015N021P038P067(0) <='1';
          else
          cVar1S17S83N015N021P038P067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='0' )then
          cVar1S18S83N015N021P038N067(0) <='1';
          else
          cVar1S18S83N015N021P038N067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='0' )then
          cVar1S19S83N015N021P038N067(0) <='1';
          else
          cVar1S19S83N015N021P038N067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='0' AND D(16)='0' )then
          cVar1S20S83N015N021P038N067(0) <='1';
          else
          cVar1S20S83N015N021P038N067(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='1' AND E(16)='0' )then
          cVar1S21S83N015N021P038P069(0) <='1';
          else
          cVar1S21S83N015N021P038P069(0) <='0';
          end if;
        if(A(12)='0' AND B(18)='0' AND D(15)='1' AND E(16)='0' )then
          cVar1S22S83N015N021P038P069(0) <='1';
          else
          cVar1S22S83N015N021P038P069(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='1' AND E(15)='1' )then
          cVar1S0S84P067P037P021P040nsss(0) <='1';
          else
          cVar1S0S84P067P037P021P040nsss(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S1S84P067P037P021N040(0) <='1';
          else
          cVar1S1S84P067P037P021N040(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S2S84P067P037P021N040(0) <='1';
          else
          cVar1S2S84P067P037P021N040(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='1' )then
          cVar1S3S84P067P037N021P013(0) <='1';
          else
          cVar1S3S84P067P037N021P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='1' )then
          cVar1S4S84P067P037N021P013(0) <='1';
          else
          cVar1S4S84P067P037N021P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='1' )then
          cVar1S5S84P067P037N021P013(0) <='1';
          else
          cVar1S5S84P067P037N021P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='0' )then
          cVar1S6S84P067P037N021N013(0) <='1';
          else
          cVar1S6S84P067P037N021N013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='0' )then
          cVar1S7S84P067P037N021N013(0) <='1';
          else
          cVar1S7S84P067P037N021N013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='0' AND B(18)='0' AND A(13)='0' )then
          cVar1S8S84P067P037N021N013(0) <='1';
          else
          cVar1S8S84P067P037N021N013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='1' )then
          cVar1S9S84P067P037P028nsss(0) <='1';
          else
          cVar1S9S84P067P037P028nsss(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='0' AND A(13)='0' )then
          cVar1S10S84P067P037N028P013(0) <='1';
          else
          cVar1S10S84P067P037N028P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='0' AND A(13)='0' )then
          cVar1S11S84P067P037N028P013(0) <='1';
          else
          cVar1S11S84P067P037N028P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='0' AND A(13)='0' )then
          cVar1S12S84P067P037N028P013(0) <='1';
          else
          cVar1S12S84P067P037N028P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='0' AND A(13)='1' )then
          cVar1S13S84P067P037N028P013(0) <='1';
          else
          cVar1S13S84P067P037N028P013(0) <='0';
          end if;
        if(D(16)='0' AND B(10)='1' AND B(24)='0' AND A(13)='1' )then
          cVar1S14S84P067P037N028P013(0) <='1';
          else
          cVar1S14S84P067P037N028P013(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='1' AND A(24)='0' )then
          cVar1S15S84P067P051P065P010(0) <='1';
          else
          cVar1S15S84P067P051P065P010(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='1' AND A(24)='0' )then
          cVar1S16S84P067P051P065P010(0) <='1';
          else
          cVar1S16S84P067P051P065P010(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='1' AND A(24)='1' )then
          cVar1S17S84P067P051P065P010(0) <='1';
          else
          cVar1S17S84P067P051P065P010(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='0' AND E( 9)='1' )then
          cVar1S18S84P067P051N065P064(0) <='1';
          else
          cVar1S18S84P067P051N065P064(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='0' AND E( 9)='0' )then
          cVar1S19S84P067P051N065N064(0) <='1';
          else
          cVar1S19S84P067P051N065N064(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='0' AND E( 9)='0' )then
          cVar1S20S84P067P051N065N064(0) <='1';
          else
          cVar1S20S84P067P051N065N064(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='0' AND E(17)='0' AND E( 9)='0' )then
          cVar1S21S84P067P051N065N064(0) <='1';
          else
          cVar1S21S84P067P051N065N064(0) <='0';
          end if;
        if(D(16)='1' AND D(20)='1' AND A(26)='0' AND B(21)='0' )then
          cVar1S22S84P067P051P006P034(0) <='1';
          else
          cVar1S22S84P067P051P006P034(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND D(19)='1' )then
          cVar1S0S85P037P013P048P055(0) <='1';
          else
          cVar1S0S85P037P013P048P055(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND D(19)='1' )then
          cVar1S1S85P037P013P048P055(0) <='1';
          else
          cVar1S1S85P037P013P048P055(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND D(19)='0' )then
          cVar1S2S85P037P013P048N055(0) <='1';
          else
          cVar1S2S85P037P013P048N055(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND D(19)='0' )then
          cVar1S3S85P037P013P048N055(0) <='1';
          else
          cVar1S3S85P037P013P048N055(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='0' AND D(19)='0' )then
          cVar1S4S85P037P013P048N055(0) <='1';
          else
          cVar1S4S85P037P013P048N055(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='0' AND E(13)='1' AND B(11)='0' )then
          cVar1S5S85P037P013P048P035(0) <='1';
          else
          cVar1S5S85P037P013P048P035(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND D(12)='0' )then
          cVar1S6S85P037P013P018P050(0) <='1';
          else
          cVar1S6S85P037P013P018P050(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND D(12)='0' )then
          cVar1S7S85P037P013P018P050(0) <='1';
          else
          cVar1S7S85P037P013P018P050(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND D(12)='0' )then
          cVar1S8S85P037P013P018P050(0) <='1';
          else
          cVar1S8S85P037P013P018P050(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='1' AND D(12)='0' )then
          cVar1S9S85P037P013P018P050(0) <='1';
          else
          cVar1S9S85P037P013P018P050(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='0' AND E(23)='0' )then
          cVar1S10S85P037P013N018P041(0) <='1';
          else
          cVar1S10S85P037P013N018P041(0) <='0';
          end if;
        if(B(10)='1' AND A(13)='1' AND A(20)='0' AND E(23)='0' )then
          cVar1S11S85P037P013N018P041(0) <='1';
          else
          cVar1S11S85P037P013N018P041(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='0' AND B(13)='1' )then
          cVar1S12S85N037P058P011P031nsss(0) <='1';
          else
          cVar1S12S85N037P058P011P031nsss(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='0' AND B(13)='0' )then
          cVar1S13S85N037P058P011N031(0) <='1';
          else
          cVar1S13S85N037P058P011N031(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='0' AND B(13)='0' )then
          cVar1S14S85N037P058P011N031(0) <='1';
          else
          cVar1S14S85N037P058P011N031(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='0' AND B(13)='0' )then
          cVar1S15S85N037P058P011N031(0) <='1';
          else
          cVar1S15S85N037P058P011N031(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='0' AND B(13)='0' )then
          cVar1S16S85N037P058P011N031(0) <='1';
          else
          cVar1S16S85N037P058P011N031(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='1' AND A(15)='0' )then
          cVar1S17S85N037P058P011P009(0) <='1';
          else
          cVar1S17S85N037P058P011P009(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='1' AND A(14)='1' AND A(15)='0' )then
          cVar1S18S85N037P058P011P009(0) <='1';
          else
          cVar1S18S85N037P058P011P009(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='1' AND E(15)='1' )then
          cVar1S19S85N037N058P021P040nsss(0) <='1';
          else
          cVar1S19S85N037N058P021P040nsss(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S20S85N037N058P021N040(0) <='1';
          else
          cVar1S20S85N037N058P021N040(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='1' AND E(15)='0' )then
          cVar1S21S85N037N058P021N040(0) <='1';
          else
          cVar1S21S85N037N058P021N040(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='0' AND E(13)='1' )then
          cVar1S22S85N037N058N021P048(0) <='1';
          else
          cVar1S22S85N037N058N021P048(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='0' AND E(13)='1' )then
          cVar1S23S85N037N058N021P048(0) <='1';
          else
          cVar1S23S85N037N058N021P048(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='0' AND E(13)='1' )then
          cVar1S24S85N037N058N021P048(0) <='1';
          else
          cVar1S24S85N037N058N021P048(0) <='0';
          end if;
        if(B(10)='0' AND D(10)='0' AND B(18)='0' AND E(13)='0' )then
          cVar1S25S85N037N058N021N048(0) <='1';
          else
          cVar1S25S85N037N058N021N048(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='1' )then
          cVar1S0S86P037P048P025nsss(0) <='1';
          else
          cVar1S0S86P037P048P025nsss(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND D(12)='1' )then
          cVar1S1S86P037P048N025P050(0) <='1';
          else
          cVar1S1S86P037P048N025P050(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND D(12)='1' )then
          cVar1S2S86P037P048N025P050(0) <='1';
          else
          cVar1S2S86P037P048N025P050(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND D(12)='0' )then
          cVar1S3S86P037P048N025N050(0) <='1';
          else
          cVar1S3S86P037P048N025N050(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='1' AND B(16)='0' AND D(12)='0' )then
          cVar1S4S86P037P048N025N050(0) <='1';
          else
          cVar1S4S86P037P048N025N050(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='1' )then
          cVar1S5S86P037N048P046P036(0) <='1';
          else
          cVar1S5S86P037N048P046P036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='1' )then
          cVar1S6S86P037N048P046P036(0) <='1';
          else
          cVar1S6S86P037N048P046P036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='1' )then
          cVar1S7S86P037N048P046P036(0) <='1';
          else
          cVar1S7S86P037N048P046P036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='0' )then
          cVar1S8S86P037N048P046N036(0) <='1';
          else
          cVar1S8S86P037N048P046N036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='0' )then
          cVar1S9S86P037N048P046N036(0) <='1';
          else
          cVar1S9S86P037N048P046N036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='0' AND B(20)='0' )then
          cVar1S10S86P037N048P046N036(0) <='1';
          else
          cVar1S10S86P037N048P046N036(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='1' AND D( 9)='0' )then
          cVar1S11S86P037N048P046P062(0) <='1';
          else
          cVar1S11S86P037N048P046P062(0) <='0';
          end if;
        if(B(10)='0' AND E(13)='0' AND D(13)='1' AND D( 9)='0' )then
          cVar1S12S86P037N048P046P062(0) <='1';
          else
          cVar1S12S86P037N048P046P062(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='0' AND B(13)='1' AND B(11)='0' )then
          cVar1S13S86P037P004P031P035(0) <='1';
          else
          cVar1S13S86P037P004P031P035(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='0' AND B(13)='0' AND D(19)='1' )then
          cVar1S14S86P037P004N031P055(0) <='1';
          else
          cVar1S14S86P037P004N031P055(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='0' AND B(13)='0' AND D(19)='1' )then
          cVar1S15S86P037P004N031P055(0) <='1';
          else
          cVar1S15S86P037P004N031P055(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='0' AND B(13)='0' AND D(19)='0' )then
          cVar1S16S86P037P004N031N055(0) <='1';
          else
          cVar1S16S86P037P004N031N055(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='0' AND B(13)='0' AND D(19)='0' )then
          cVar1S17S86P037P004N031N055(0) <='1';
          else
          cVar1S17S86P037P004N031N055(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='1' AND D(20)='0' AND B(20)='0' )then
          cVar1S18S86P037P004P051P036(0) <='1';
          else
          cVar1S18S86P037P004P051P036(0) <='0';
          end if;
        if(B(10)='1' AND A(27)='1' AND D(20)='0' AND B(20)='0' )then
          cVar1S19S86P037P004P051P036(0) <='1';
          else
          cVar1S19S86P037P004P051P036(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='1' AND B(25)='0' )then
          cVar1S0S87P019P017P035P026(0) <='1';
          else
          cVar1S0S87P019P017P035P026(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='1' AND B(25)='0' )then
          cVar1S1S87P019P017P035P026(0) <='1';
          else
          cVar1S1S87P019P017P035P026(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='1' AND B(25)='0' )then
          cVar1S2S87P019P017P035P026(0) <='1';
          else
          cVar1S2S87P019P017P035P026(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='1' AND B(25)='0' )then
          cVar1S3S87P019P017P035P026(0) <='1';
          else
          cVar1S3S87P019P017P035P026(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='1' )then
          cVar1S4S87P019P017N035P066(0) <='1';
          else
          cVar1S4S87P019P017N035P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='1' )then
          cVar1S5S87P019P017N035P066(0) <='1';
          else
          cVar1S5S87P019P017N035P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='1' )then
          cVar1S6S87P019P017N035P066(0) <='1';
          else
          cVar1S6S87P019P017N035P066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='0' )then
          cVar1S7S87P019P017N035N066(0) <='1';
          else
          cVar1S7S87P019P017N035N066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='0' )then
          cVar1S8S87P019P017N035N066(0) <='1';
          else
          cVar1S8S87P019P017N035N066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='0' AND B(11)='0' AND D( 8)='0' )then
          cVar1S9S87P019P017N035N066(0) <='1';
          else
          cVar1S9S87P019P017N035N066(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='0' AND B(14)='0' )then
          cVar1S10S87P019P017P053P029(0) <='1';
          else
          cVar1S10S87P019P017P053P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='0' AND B(14)='0' )then
          cVar1S11S87P019P017P053P029(0) <='1';
          else
          cVar1S11S87P019P017P053P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='0' AND B(14)='1' )then
          cVar1S12S87P019P017P053P029(0) <='1';
          else
          cVar1S12S87P019P017P053P029(0) <='0';
          end if;
        if(A(10)='1' AND A(11)='1' AND E(20)='1' AND B(10)='1' )then
          cVar1S13S87P019P017P053P037(0) <='1';
          else
          cVar1S13S87P019P017P053P037(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='1' AND E( 8)='0' AND D(23)='0' )then
          cVar1S14S87N019P009P068P039(0) <='1';
          else
          cVar1S14S87N019P009P068P039(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='1' AND E( 8)='0' AND D(23)='0' )then
          cVar1S15S87N019P009P068P039(0) <='1';
          else
          cVar1S15S87N019P009P068P039(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='1' AND E( 8)='0' AND D(23)='0' )then
          cVar1S16S87N019P009P068P039(0) <='1';
          else
          cVar1S16S87N019P009P068P039(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='1' AND E( 8)='1' AND E(20)='1' )then
          cVar1S17S87N019P009P068P053nsss(0) <='1';
          else
          cVar1S17S87N019P009P068P053nsss(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='1' AND B(18)='1' )then
          cVar1S18S87N019N009P040P021nsss(0) <='1';
          else
          cVar1S18S87N019N009P040P021nsss(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='1' AND B(18)='0' )then
          cVar1S19S87N019N009P040N021(0) <='1';
          else
          cVar1S19S87N019N009P040N021(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='1' AND B(18)='0' )then
          cVar1S20S87N019N009P040N021(0) <='1';
          else
          cVar1S20S87N019N009P040N021(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='1' AND B(18)='0' )then
          cVar1S21S87N019N009P040N021(0) <='1';
          else
          cVar1S21S87N019N009P040N021(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S22S87N019N009N040P038(0) <='1';
          else
          cVar1S22S87N019N009N040P038(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S23S87N019N009N040P038(0) <='1';
          else
          cVar1S23S87N019N009N040P038(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='0' AND D(15)='0' )then
          cVar1S24S87N019N009N040P038(0) <='1';
          else
          cVar1S24S87N019N009N040P038(0) <='0';
          end if;
        if(A(10)='0' AND A(15)='0' AND E(15)='0' AND D(15)='1' )then
          cVar1S25S87N019N009N040P038(0) <='1';
          else
          cVar1S25S87N019N009N040P038(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='0' AND D(17)='0' )then
          cVar1S0S88P060P009P068P063(0) <='1';
          else
          cVar1S0S88P060P009P068P063(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='0' AND D(17)='0' )then
          cVar1S1S88P060P009P068P063(0) <='1';
          else
          cVar1S1S88P060P009P068P063(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='0' AND D(17)='0' )then
          cVar1S2S88P060P009P068P063(0) <='1';
          else
          cVar1S2S88P060P009P068P063(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='0' AND D(17)='1' )then
          cVar1S3S88P060P009P068P063(0) <='1';
          else
          cVar1S3S88P060P009P068P063(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='0' AND D(17)='1' )then
          cVar1S4S88P060P009P068P063(0) <='1';
          else
          cVar1S4S88P060P009P068P063(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='1' AND A(28)='0' )then
          cVar1S5S88P060P009P068P002(0) <='1';
          else
          cVar1S5S88P060P009P068P002(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='1' AND E( 8)='1' AND A(28)='0' )then
          cVar1S6S88P060P009P068P002(0) <='1';
          else
          cVar1S6S88P060P009P068P002(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='0' AND D(19)='1' )then
          cVar1S7S88P060N009P053P055(0) <='1';
          else
          cVar1S7S88P060N009P053P055(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='0' AND D(19)='0' )then
          cVar1S8S88P060N009P053N055(0) <='1';
          else
          cVar1S8S88P060N009P053N055(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='0' AND D(19)='0' )then
          cVar1S9S88P060N009P053N055(0) <='1';
          else
          cVar1S9S88P060N009P053N055(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='0' AND D(19)='0' )then
          cVar1S10S88P060N009P053N055(0) <='1';
          else
          cVar1S10S88P060N009P053N055(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='1' AND B(24)='1' )then
          cVar1S11S88P060N009P053P028nsss(0) <='1';
          else
          cVar1S11S88P060N009P053P028nsss(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='1' AND B(24)='0' )then
          cVar1S12S88P060N009P053N028(0) <='1';
          else
          cVar1S12S88P060N009P053N028(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='1' AND B(24)='0' )then
          cVar1S13S88P060N009P053N028(0) <='1';
          else
          cVar1S13S88P060N009P053N028(0) <='0';
          end if;
        if(E(10)='0' AND A(15)='0' AND E(20)='1' AND B(24)='0' )then
          cVar1S14S88P060N009P053N028(0) <='1';
          else
          cVar1S14S88P060N009P053N028(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='1' AND D(20)='0' )then
          cVar1S15S88P060P039P062P051(0) <='1';
          else
          cVar1S15S88P060P039P062P051(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='1' AND D(20)='0' )then
          cVar1S16S88P060P039P062P051(0) <='1';
          else
          cVar1S16S88P060P039P062P051(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='0' AND B(13)='1' )then
          cVar1S17S88P060P039N062P031(0) <='1';
          else
          cVar1S17S88P060P039N062P031(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='0' AND B(13)='1' )then
          cVar1S18S88P060P039N062P031(0) <='1';
          else
          cVar1S18S88P060P039N062P031(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='0' AND B(13)='0' )then
          cVar1S19S88P060P039N062N031(0) <='1';
          else
          cVar1S19S88P060P039N062N031(0) <='0';
          end if;
        if(E(10)='1' AND D(23)='0' AND D( 9)='0' AND B(13)='0' )then
          cVar1S20S88P060P039N062N031(0) <='1';
          else
          cVar1S20S88P060P039N062N031(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='0' AND D(17)='0' AND A(16)='1' )then
          cVar1S0S89P009P068P063P007(0) <='1';
          else
          cVar1S0S89P009P068P063P007(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='0' AND D(17)='0' AND A(16)='1' )then
          cVar1S1S89P009P068P063P007(0) <='1';
          else
          cVar1S1S89P009P068P063P007(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='0' AND D(17)='0' AND A(16)='0' )then
          cVar1S2S89P009P068P063N007(0) <='1';
          else
          cVar1S2S89P009P068P063N007(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='0' AND D(17)='1' AND A(25)='0' )then
          cVar1S3S89P009P068P063P008(0) <='1';
          else
          cVar1S3S89P009P068P063P008(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='1' AND A(28)='0' AND D(21)='1' )then
          cVar1S4S89P009P068P002P047nsss(0) <='1';
          else
          cVar1S4S89P009P068P002P047nsss(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='1' AND A(28)='0' AND D(21)='0' )then
          cVar1S5S89P009P068P002N047(0) <='1';
          else
          cVar1S5S89P009P068P002N047(0) <='0';
          end if;
        if(A(15)='1' AND E( 8)='1' AND A(28)='0' AND D(21)='0' )then
          cVar1S6S89P009P068P002N047(0) <='1';
          else
          cVar1S6S89P009P068P002N047(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='1' AND A(17)='1' )then
          cVar1S7S89N009P049P023P005nsss(0) <='1';
          else
          cVar1S7S89N009P049P023P005nsss(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S8S89N009P049P023N005(0) <='1';
          else
          cVar1S8S89N009P049P023N005(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S9S89N009P049P023N005(0) <='1';
          else
          cVar1S9S89N009P049P023N005(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='1' AND A(17)='0' )then
          cVar1S10S89N009P049P023N005(0) <='1';
          else
          cVar1S10S89N009P049P023N005(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='0' AND D(22)='0' )then
          cVar1S11S89N009P049N023P043(0) <='1';
          else
          cVar1S11S89N009P049N023P043(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='0' AND D(22)='0' )then
          cVar1S12S89N009P049N023P043(0) <='1';
          else
          cVar1S12S89N009P049N023P043(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='0' AND D(22)='1' )then
          cVar1S13S89N009P049N023P043(0) <='1';
          else
          cVar1S13S89N009P049N023P043(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='0' AND D(22)='1' )then
          cVar1S14S89N009P049N023P043(0) <='1';
          else
          cVar1S14S89N009P049N023P043(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='0' AND B(17)='0' AND D(22)='1' )then
          cVar1S15S89N009P049N023P043(0) <='1';
          else
          cVar1S15S89N009P049N023P043(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='1' AND B(25)='1' AND A(22)='0' )then
          cVar1S16S89N009P049P026P014nsss(0) <='1';
          else
          cVar1S16S89N009P049P026P014nsss(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='1' AND B(25)='0' AND B(26)='1' )then
          cVar1S17S89N009P049N026P024(0) <='1';
          else
          cVar1S17S89N009P049N026P024(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='1' AND B(25)='0' AND B(26)='0' )then
          cVar1S18S89N009P049N026N024(0) <='1';
          else
          cVar1S18S89N009P049N026N024(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='1' AND B(25)='0' AND B(26)='0' )then
          cVar1S19S89N009P049N026N024(0) <='1';
          else
          cVar1S19S89N009P049N026N024(0) <='0';
          end if;
        if(A(15)='0' AND E(21)='1' AND B(25)='0' AND B(26)='0' )then
          cVar1S20S89N009P049N026N024(0) <='1';
          else
          cVar1S20S89N009P049N026N024(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='1' AND E(16)='0' )then
          cVar1S0S90P049P052P065P069nsss(0) <='1';
          else
          cVar1S0S90P049P052P065P069nsss(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='1' )then
          cVar1S1S90P049P052N065P062(0) <='1';
          else
          cVar1S1S90P049P052N065P062(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S2S90P049P052N065N062(0) <='1';
          else
          cVar1S2S90P049P052N065N062(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S3S90P049P052N065N062(0) <='1';
          else
          cVar1S3S90P049P052N065N062(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S4S90P049P052N065N062(0) <='1';
          else
          cVar1S4S90P049P052N065N062(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S5S90P049P052N065N062(0) <='1';
          else
          cVar1S5S90P049P052N065N062(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='1' )then
          cVar1S6S90P049N052P029P055(0) <='1';
          else
          cVar1S6S90P049N052P029P055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='1' )then
          cVar1S7S90P049N052P029P055(0) <='1';
          else
          cVar1S7S90P049N052P029P055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='0' )then
          cVar1S8S90P049N052P029N055(0) <='1';
          else
          cVar1S8S90P049N052P029N055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='0' )then
          cVar1S9S90P049N052P029N055(0) <='1';
          else
          cVar1S9S90P049N052P029N055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='0' )then
          cVar1S10S90P049N052P029N055(0) <='1';
          else
          cVar1S10S90P049N052P029N055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='0' AND D(19)='0' )then
          cVar1S11S90P049N052P029N055(0) <='1';
          else
          cVar1S11S90P049N052P029N055(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='1' AND E(11)='1' )then
          cVar1S12S90P049N052P029P056(0) <='1';
          else
          cVar1S12S90P049N052P029P056(0) <='0';
          end if;
        if(E(21)='0' AND E(12)='0' AND B(14)='1' AND E(11)='0' )then
          cVar1S13S90P049N052P029N056(0) <='1';
          else
          cVar1S13S90P049N052P029N056(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='1' AND D(17)='0' )then
          cVar1S14S90P049P026P063nsss(0) <='1';
          else
          cVar1S14S90P049P026P063nsss(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='0' AND B(15)='1' AND A(15)='1' )then
          cVar1S15S90P049N026P027P009nsss(0) <='1';
          else
          cVar1S15S90P049N026P027P009nsss(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='0' AND B(15)='0' AND B(26)='1' )then
          cVar1S16S90P049N026N027P024(0) <='1';
          else
          cVar1S16S90P049N026N027P024(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S17S90P049N026N027N024(0) <='1';
          else
          cVar1S17S90P049N026N027N024(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S18S90P049N026N027N024(0) <='1';
          else
          cVar1S18S90P049N026N027N024(0) <='0';
          end if;
        if(E(21)='1' AND B(25)='0' AND B(15)='0' AND B(26)='0' )then
          cVar1S19S90P049N026N027N024(0) <='1';
          else
          cVar1S19S90P049N026N027N024(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='1' AND E(16)='0' )then
          cVar1S0S91P052P065P069nsss(0) <='1';
          else
          cVar1S0S91P052P065P069nsss(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='1' AND B(11)='0' )then
          cVar1S1S91P052N065P062P035nsss(0) <='1';
          else
          cVar1S1S91P052N065P062P035nsss(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='0' AND D(12)='1' )then
          cVar1S2S91P052N065N062P050(0) <='1';
          else
          cVar1S2S91P052N065N062P050(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='0' AND D(12)='1' )then
          cVar1S3S91P052N065N062P050(0) <='1';
          else
          cVar1S3S91P052N065N062P050(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='0' AND D(12)='0' )then
          cVar1S4S91P052N065N062N050(0) <='1';
          else
          cVar1S4S91P052N065N062N050(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='0' AND D(12)='0' )then
          cVar1S5S91P052N065N062N050(0) <='1';
          else
          cVar1S5S91P052N065N062N050(0) <='0';
          end if;
        if(E(12)='1' AND E(17)='0' AND D( 9)='0' AND D(12)='0' )then
          cVar1S6S91P052N065N062N050(0) <='1';
          else
          cVar1S6S91P052N065N062N050(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='0' AND A(16)='1' )then
          cVar1S7S91N052P048P061P007(0) <='1';
          else
          cVar1S7S91N052P048P061P007(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='0' AND A(16)='1' )then
          cVar1S8S91N052P048P061P007(0) <='1';
          else
          cVar1S8S91N052P048P061P007(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='0' AND A(16)='0' )then
          cVar1S9S91N052P048P061N007(0) <='1';
          else
          cVar1S9S91N052P048P061N007(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='0' AND A(16)='0' )then
          cVar1S10S91N052P048P061N007(0) <='1';
          else
          cVar1S10S91N052P048P061N007(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='0' AND A(16)='0' )then
          cVar1S11S91N052P048P061N007(0) <='1';
          else
          cVar1S11S91N052P048P061N007(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='1' AND E(18)='1' AND A(22)='1' )then
          cVar1S12S91N052P048P061P014nsss(0) <='1';
          else
          cVar1S12S91N052P048P061P014nsss(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='0' AND D(12)='0' AND D(19)='1' )then
          cVar1S13S91N052N048P050P055(0) <='1';
          else
          cVar1S13S91N052N048P050P055(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='0' AND D(12)='0' AND D(19)='0' )then
          cVar1S14S91N052N048P050N055(0) <='1';
          else
          cVar1S14S91N052N048P050N055(0) <='0';
          end if;
        if(E(12)='0' AND E(13)='0' AND D(12)='1' AND A(27)='0' )then
          cVar1S15S91N052N048P050P004(0) <='1';
          else
          cVar1S15S91N052N048P050P004(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='1' AND D(11)='1' )then
          cVar1S0S92P019P068P029P054nsss(0) <='1';
          else
          cVar1S0S92P019P068P029P054nsss(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='1' AND D(11)='0' )then
          cVar1S1S92P019P068P029N054(0) <='1';
          else
          cVar1S1S92P019P068P029N054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='1' AND D(11)='0' )then
          cVar1S2S92P019P068P029N054(0) <='1';
          else
          cVar1S2S92P019P068P029N054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='1' AND D(11)='0' )then
          cVar1S3S92P019P068P029N054(0) <='1';
          else
          cVar1S3S92P019P068P029N054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S4S92P019P068N029P054(0) <='1';
          else
          cVar1S4S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S5S92P019P068N029P054(0) <='1';
          else
          cVar1S5S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S6S92P019P068N029P054(0) <='1';
          else
          cVar1S6S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S7S92P019P068N029P054(0) <='1';
          else
          cVar1S7S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S8S92P019P068N029P054(0) <='1';
          else
          cVar1S8S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S9S92P019P068N029P054(0) <='1';
          else
          cVar1S9S92P019P068N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND D(19)='0' AND D(12)='1' )then
          cVar1S10S92P019P068P055P050(0) <='1';
          else
          cVar1S10S92P019P068P055P050(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND D(19)='0' AND D(12)='0' )then
          cVar1S11S92P019P068P055N050(0) <='1';
          else
          cVar1S11S92P019P068P055N050(0) <='0';
          end if;
        if(A(10)='0' AND E( 8)='1' AND D(19)='1' AND A(24)='1' )then
          cVar1S12S92P019P068P055P010nsss(0) <='1';
          else
          cVar1S12S92P019P068P055P010nsss(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='0' AND D(13)='1' )then
          cVar1S13S92P019P066P009P046nsss(0) <='1';
          else
          cVar1S13S92P019P066P009P046nsss(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='0' AND D(13)='0' )then
          cVar1S14S92P019P066P009N046(0) <='1';
          else
          cVar1S14S92P019P066P009N046(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='0' AND D(13)='0' )then
          cVar1S15S92P019P066P009N046(0) <='1';
          else
          cVar1S15S92P019P066P009N046(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='0' AND D(13)='0' )then
          cVar1S16S92P019P066P009N046(0) <='1';
          else
          cVar1S16S92P019P066P009N046(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='1' AND E( 8)='1' )then
          cVar1S17S92P019P066P009P068(0) <='1';
          else
          cVar1S17S92P019P066P009P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='1' AND A(15)='1' AND E( 8)='1' )then
          cVar1S18S92P019P066P009P068(0) <='1';
          else
          cVar1S18S92P019P066P009P068(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='0' AND E(18)='0' )then
          cVar1S19S92P019N066P051P061(0) <='1';
          else
          cVar1S19S92P019N066P051P061(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='0' AND E(18)='0' )then
          cVar1S20S92P019N066P051P061(0) <='1';
          else
          cVar1S20S92P019N066P051P061(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='0' AND E(18)='0' )then
          cVar1S21S92P019N066P051P061(0) <='1';
          else
          cVar1S21S92P019N066P051P061(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='0' AND E(18)='1' )then
          cVar1S22S92P019N066P051P061(0) <='1';
          else
          cVar1S22S92P019N066P051P061(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='0' AND E(18)='1' )then
          cVar1S23S92P019N066P051P061(0) <='1';
          else
          cVar1S23S92P019N066P051P061(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='1' AND A(21)='0' )then
          cVar1S24S92P019N066P051P016(0) <='1';
          else
          cVar1S24S92P019N066P051P016(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='1' AND A(21)='0' )then
          cVar1S25S92P019N066P051P016(0) <='1';
          else
          cVar1S25S92P019N066P051P016(0) <='0';
          end if;
        if(A(10)='1' AND D( 8)='0' AND D(20)='1' AND A(21)='1' )then
          cVar1S26S92P019N066P051P016(0) <='1';
          else
          cVar1S26S92P019N066P051P016(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='1' )then
          cVar1S0S93P019P051P002P000(0) <='1';
          else
          cVar1S0S93P019P051P002P000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='1' )then
          cVar1S1S93P019P051P002P000(0) <='1';
          else
          cVar1S1S93P019P051P002P000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='1' )then
          cVar1S2S93P019P051P002P000(0) <='1';
          else
          cVar1S2S93P019P051P002P000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='0' )then
          cVar1S3S93P019P051P002N000(0) <='1';
          else
          cVar1S3S93P019P051P002N000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='0' )then
          cVar1S4S93P019P051P002N000(0) <='1';
          else
          cVar1S4S93P019P051P002N000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='0' )then
          cVar1S5S93P019P051P002N000(0) <='1';
          else
          cVar1S5S93P019P051P002N000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='0' AND A(29)='0' )then
          cVar1S6S93P019P051P002N000(0) <='1';
          else
          cVar1S6S93P019P051P002N000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(28)='1' AND D(11)='0' )then
          cVar1S7S93P019P051P002P054(0) <='1';
          else
          cVar1S7S93P019P051P002P054(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(26)='0' AND B(10)='1' )then
          cVar1S8S93P019P051P024P037(0) <='1';
          else
          cVar1S8S93P019P051P024P037(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(26)='0' AND B(10)='0' )then
          cVar1S9S93P019P051P024N037(0) <='1';
          else
          cVar1S9S93P019P051P024N037(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(26)='0' AND B(10)='0' )then
          cVar1S10S93P019P051P024N037(0) <='1';
          else
          cVar1S10S93P019P051P024N037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='1' AND D(11)='1' AND A(13)='1' )then
          cVar1S11S93N019P056P054P013nsss(0) <='1';
          else
          cVar1S11S93N019P056P054P013nsss(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='1' AND D(11)='1' AND A(13)='0' )then
          cVar1S12S93N019P056P054N013(0) <='1';
          else
          cVar1S12S93N019P056P054N013(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='1' AND D(11)='0' AND D(10)='1' )then
          cVar1S13S93N019P056N054P058(0) <='1';
          else
          cVar1S13S93N019P056N054P058(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='1' AND D(11)='0' AND D(10)='1' )then
          cVar1S14S93N019P056N054P058(0) <='1';
          else
          cVar1S14S93N019P056N054P058(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='1' AND D(11)='0' AND D(10)='0' )then
          cVar1S15S93N019P056N054N058(0) <='1';
          else
          cVar1S15S93N019P056N054N058(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='0' AND B(10)='1' )then
          cVar1S16S93N019N056P054P037(0) <='1';
          else
          cVar1S16S93N019N056P054P037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='0' AND B(10)='1' )then
          cVar1S17S93N019N056P054P037(0) <='1';
          else
          cVar1S17S93N019N056P054P037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='0' AND B(10)='0' )then
          cVar1S18S93N019N056P054N037(0) <='1';
          else
          cVar1S18S93N019N056P054N037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='0' AND B(10)='0' )then
          cVar1S19S93N019N056P054N037(0) <='1';
          else
          cVar1S19S93N019N056P054N037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='0' AND B(10)='0' )then
          cVar1S20S93N019N056P054N037(0) <='1';
          else
          cVar1S20S93N019N056P054N037(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='1' AND A(17)='0' )then
          cVar1S21S93N019N056P054P005(0) <='1';
          else
          cVar1S21S93N019N056P054P005(0) <='0';
          end if;
        if(A(10)='0' AND E(11)='0' AND D(11)='1' AND A(17)='0' )then
          cVar1S22S93N019N056P054P005(0) <='1';
          else
          cVar1S22S93N019N056P054P005(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S0S94P019P037P029P011(0) <='1';
          else
          cVar1S0S94P019P037P029P011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S1S94P019P037P029P011(0) <='1';
          else
          cVar1S1S94P019P037P029P011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S2S94P019P037P029P011(0) <='1';
          else
          cVar1S2S94P019P037P029P011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S3S94P019P037P029N011(0) <='1';
          else
          cVar1S3S94P019P037P029N011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S4S94P019P037P029N011(0) <='1';
          else
          cVar1S4S94P019P037P029N011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S5S94P019P037P029N011(0) <='1';
          else
          cVar1S5S94P019P037P029N011(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='0' AND E(22)='1' )then
          cVar1S6S94P019P037N029P045(0) <='1';
          else
          cVar1S6S94P019P037N029P045(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='0' AND E(22)='1' )then
          cVar1S7S94P019P037N029P045(0) <='1';
          else
          cVar1S7S94P019P037N029P045(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='0' AND E(22)='1' )then
          cVar1S8S94P019P037N029P045(0) <='1';
          else
          cVar1S8S94P019P037N029P045(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='0' AND E(22)='0' )then
          cVar1S9S94P019P037N029N045(0) <='1';
          else
          cVar1S9S94P019P037N029N045(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND B(14)='0' AND E(22)='0' )then
          cVar1S10S94P019P037N029N045(0) <='1';
          else
          cVar1S10S94P019P037N029N045(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='0' AND B(24)='1' )then
          cVar1S11S94P019P037P059P028nsss(0) <='1';
          else
          cVar1S11S94P019P037P059P028nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='0' AND B(24)='0' )then
          cVar1S12S94P019P037P059N028(0) <='1';
          else
          cVar1S12S94P019P037P059N028(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='1' AND E( 9)='0' )then
          cVar1S13S94P019P037P059P064(0) <='1';
          else
          cVar1S13S94P019P037P059P064(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='1' AND E( 9)='0' )then
          cVar1S14S94P019P037P059P064(0) <='1';
          else
          cVar1S14S94P019P037P059P064(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='1' AND D(20)='0' AND B(14)='0' )then
          cVar1S15S94P019P069P051P029(0) <='1';
          else
          cVar1S15S94P019P069P051P029(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='1' AND D(20)='0' AND B(14)='0' )then
          cVar1S16S94P019P069P051P029(0) <='1';
          else
          cVar1S16S94P019P069P051P029(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='1' AND D(20)='1' AND A(13)='0' )then
          cVar1S17S94P019P069P051P013(0) <='1';
          else
          cVar1S17S94P019P069P051P013(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='0' AND B(23)='0' )then
          cVar1S18S94P019N069P057P030(0) <='1';
          else
          cVar1S18S94P019N069P057P030(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='0' AND B(23)='0' )then
          cVar1S19S94P019N069P057P030(0) <='1';
          else
          cVar1S19S94P019N069P057P030(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='0' AND B(23)='0' )then
          cVar1S20S94P019N069P057P030(0) <='1';
          else
          cVar1S20S94P019N069P057P030(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='1' AND E(18)='0' )then
          cVar1S21S94P019N069P057P061(0) <='1';
          else
          cVar1S21S94P019N069P057P061(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='1' AND E(18)='0' )then
          cVar1S22S94P019N069P057P061(0) <='1';
          else
          cVar1S22S94P019N069P057P061(0) <='0';
          end if;
        if(A(10)='1' AND E(16)='0' AND E(19)='1' AND E(18)='0' )then
          cVar1S23S94P019N069P057P061(0) <='1';
          else
          cVar1S23S94P019N069P057P061(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='1' AND A(15)='1' )then
          cVar1S0S95P019P057P036P009(0) <='1';
          else
          cVar1S0S95P019P057P036P009(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='1' AND A(15)='1' )then
          cVar1S1S95P019P057P036P009(0) <='1';
          else
          cVar1S1S95P019P057P036P009(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='1' AND A(15)='1' )then
          cVar1S2S95P019P057P036P009(0) <='1';
          else
          cVar1S2S95P019P057P036P009(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='1' AND A(15)='0' )then
          cVar1S3S95P019P057P036N009(0) <='1';
          else
          cVar1S3S95P019P057P036N009(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='1' AND A(15)='0' )then
          cVar1S4S95P019P057P036N009(0) <='1';
          else
          cVar1S4S95P019P057P036N009(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='0' AND E(11)='0' )then
          cVar1S5S95P019P057N036P056(0) <='1';
          else
          cVar1S5S95P019P057N036P056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='0' AND E(11)='0' )then
          cVar1S6S95P019P057N036P056(0) <='1';
          else
          cVar1S6S95P019P057N036P056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='0' AND E(11)='0' )then
          cVar1S7S95P019P057N036P056(0) <='1';
          else
          cVar1S7S95P019P057N036P056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='0' AND E(11)='1' )then
          cVar1S8S95P019P057N036P056(0) <='1';
          else
          cVar1S8S95P019P057N036P056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='0' AND B(20)='0' AND E(11)='1' )then
          cVar1S9S95P019P057N036P056(0) <='1';
          else
          cVar1S9S95P019P057N036P056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='1' AND B(23)='1' AND E(11)='1' )then
          cVar1S10S95P019P057P030P056nsss(0) <='1';
          else
          cVar1S10S95P019P057P030P056nsss(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='1' AND B(23)='1' AND E(11)='0' )then
          cVar1S11S95P019P057P030N056(0) <='1';
          else
          cVar1S11S95P019P057P030N056(0) <='0';
          end if;
        if(A(10)='1' AND E(19)='1' AND B(23)='0' AND A(27)='0' )then
          cVar1S12S95P019P057N030P004(0) <='1';
          else
          cVar1S12S95P019P057N030P004(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND D( 9)='0' AND A(17)='1' )then
          cVar1S13S95N019P045P062P005nsss(0) <='1';
          else
          cVar1S13S95N019P045P062P005nsss(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND D( 9)='0' AND A(17)='0' )then
          cVar1S14S95N019P045P062N005(0) <='1';
          else
          cVar1S14S95N019P045P062N005(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND D( 9)='0' AND A(17)='0' )then
          cVar1S15S95N019P045P062N005(0) <='1';
          else
          cVar1S15S95N019P045P062N005(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S16S95N019N045P029P011(0) <='1';
          else
          cVar1S16S95N019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S17S95N019N045P029P011(0) <='1';
          else
          cVar1S17S95N019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S18S95N019N045P029P011(0) <='1';
          else
          cVar1S18S95N019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S19S95N019N045P029N011(0) <='1';
          else
          cVar1S19S95N019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S20S95N019N045P029N011(0) <='1';
          else
          cVar1S20S95N019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='1' )then
          cVar1S21S95N019N045N029P031(0) <='1';
          else
          cVar1S21S95N019N045N029P031(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='1' )then
          cVar1S22S95N019N045N029P031(0) <='1';
          else
          cVar1S22S95N019N045N029P031(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='1' )then
          cVar1S23S95N019N045N029P031(0) <='1';
          else
          cVar1S23S95N019N045N029P031(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='0' )then
          cVar1S24S95N019N045N029N031(0) <='1';
          else
          cVar1S24S95N019N045N029N031(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='0' )then
          cVar1S25S95N019N045N029N031(0) <='1';
          else
          cVar1S25S95N019N045N029N031(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND B(13)='0' )then
          cVar1S26S95N019N045N029N031(0) <='1';
          else
          cVar1S26S95N019N045N029N031(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='1' AND A(17)='1' )then
          cVar1S0S96P019P037P045P005nsss(0) <='1';
          else
          cVar1S0S96P019P037P045P005nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='1' AND A(17)='0' )then
          cVar1S1S96P019P037P045N005(0) <='1';
          else
          cVar1S1S96P019P037P045N005(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='1' AND A(17)='0' )then
          cVar1S2S96P019P037P045N005(0) <='1';
          else
          cVar1S2S96P019P037P045N005(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='1' )then
          cVar1S3S96P019P037N045P029(0) <='1';
          else
          cVar1S3S96P019P037N045P029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='1' )then
          cVar1S4S96P019P037N045P029(0) <='1';
          else
          cVar1S4S96P019P037N045P029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='1' )then
          cVar1S5S96P019P037N045P029(0) <='1';
          else
          cVar1S5S96P019P037N045P029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='0' )then
          cVar1S6S96P019P037N045N029(0) <='1';
          else
          cVar1S6S96P019P037N045N029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='0' )then
          cVar1S7S96P019P037N045N029(0) <='1';
          else
          cVar1S7S96P019P037N045N029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='0' AND E(22)='0' AND B(14)='0' )then
          cVar1S8S96P019P037N045N029(0) <='1';
          else
          cVar1S8S96P019P037N045N029(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='0' AND B(24)='1' )then
          cVar1S9S96P019P037P059P028nsss(0) <='1';
          else
          cVar1S9S96P019P037P059P028nsss(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='0' AND B(24)='0' )then
          cVar1S10S96P019P037P059N028(0) <='1';
          else
          cVar1S10S96P019P037P059N028(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='0' AND B(24)='0' )then
          cVar1S11S96P019P037P059N028(0) <='1';
          else
          cVar1S11S96P019P037P059N028(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='1' AND E( 9)='0' )then
          cVar1S12S96P019P037P059P064(0) <='1';
          else
          cVar1S12S96P019P037P059P064(0) <='0';
          end if;
        if(A(10)='0' AND B(10)='1' AND D(18)='1' AND E( 9)='0' )then
          cVar1S13S96P019P037P059P064(0) <='1';
          else
          cVar1S13S96P019P037P059P064(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='0' AND A(15)='1' )then
          cVar1S14S96P019P036P006P009(0) <='1';
          else
          cVar1S14S96P019P036P006P009(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='0' AND A(15)='0' )then
          cVar1S15S96P019P036P006N009(0) <='1';
          else
          cVar1S15S96P019P036P006N009(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='0' AND A(15)='0' )then
          cVar1S16S96P019P036P006N009(0) <='1';
          else
          cVar1S16S96P019P036P006N009(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='0' AND A(15)='0' )then
          cVar1S17S96P019P036P006N009(0) <='1';
          else
          cVar1S17S96P019P036P006N009(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='1' AND A(27)='0' )then
          cVar1S18S96P019P036P006P004(0) <='1';
          else
          cVar1S18S96P019P036P006P004(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='1' AND A(26)='1' AND A(27)='0' )then
          cVar1S19S96P019P036P006P004(0) <='1';
          else
          cVar1S19S96P019P036P006P004(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='1' )then
          cVar1S20S96P019N036P009P063(0) <='1';
          else
          cVar1S20S96P019N036P009P063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='1' )then
          cVar1S21S96P019N036P009P063(0) <='1';
          else
          cVar1S21S96P019N036P009P063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='1' )then
          cVar1S22S96P019N036P009P063(0) <='1';
          else
          cVar1S22S96P019N036P009P063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='0' )then
          cVar1S23S96P019N036P009N063(0) <='1';
          else
          cVar1S23S96P019N036P009N063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='0' )then
          cVar1S24S96P019N036P009N063(0) <='1';
          else
          cVar1S24S96P019N036P009N063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='0' AND D(17)='0' )then
          cVar1S25S96P019N036P009N063(0) <='1';
          else
          cVar1S25S96P019N036P009N063(0) <='0';
          end if;
        if(A(10)='1' AND B(20)='0' AND A(15)='1' AND B(24)='0' )then
          cVar1S26S96P019N036P009P028(0) <='1';
          else
          cVar1S26S96P019N036P009P028(0) <='0';
          end if;
        if(E(22)='1' AND B(11)='0' AND B(16)='1' )then
          cVar1S0S97P045P035P025nsss(0) <='1';
          else
          cVar1S0S97P045P035P025nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(11)='0' AND B(16)='0' AND B(27)='1' )then
          cVar1S1S97P045P035N025P022nsss(0) <='1';
          else
          cVar1S1S97P045P035N025P022nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(11)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S2S97P045P035N025N022(0) <='1';
          else
          cVar1S2S97P045P035N025N022(0) <='0';
          end if;
        if(E(22)='1' AND B(11)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S3S97P045P035N025N022(0) <='1';
          else
          cVar1S3S97P045P035N025N022(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='1' AND B(17)='0' )then
          cVar1S4S97N045P043P019P023(0) <='1';
          else
          cVar1S4S97N045P043P019P023(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='1' AND B(17)='0' )then
          cVar1S5S97N045P043P019P023(0) <='1';
          else
          cVar1S5S97N045P043P019P023(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='1' AND B(17)='1' )then
          cVar1S6S97N045P043P019P023(0) <='1';
          else
          cVar1S6S97N045P043P019P023(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='0' AND B(26)='0' )then
          cVar1S7S97N045P043N019P024(0) <='1';
          else
          cVar1S7S97N045P043N019P024(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='0' AND B(26)='0' )then
          cVar1S8S97N045P043N019P024(0) <='1';
          else
          cVar1S8S97N045P043N019P024(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='0' AND B(26)='0' )then
          cVar1S9S97N045P043N019P024(0) <='1';
          else
          cVar1S9S97N045P043N019P024(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='0' AND B(26)='0' )then
          cVar1S10S97N045P043N019P024(0) <='1';
          else
          cVar1S10S97N045P043N019P024(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='0' AND A(10)='0' AND B(26)='1' )then
          cVar1S11S97N045P043N019P024(0) <='1';
          else
          cVar1S11S97N045P043N019P024(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='1' AND B(27)='1' )then
          cVar1S12S97N045P043P022nsss(0) <='1';
          else
          cVar1S12S97N045P043P022nsss(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='1' AND B(27)='0' AND E(19)='1' )then
          cVar1S13S97N045P043N022P057nsss(0) <='1';
          else
          cVar1S13S97N045P043N022P057nsss(0) <='0';
          end if;
        if(E(22)='0' AND D(22)='1' AND B(27)='0' AND E(19)='0' )then
          cVar1S14S97N045P043N022N057(0) <='1';
          else
          cVar1S14S97N045P043N022N057(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S0S98P019P045P026P062(0) <='1';
          else
          cVar1S0S98P019P045P026P062(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S1S98P019P045P026P062(0) <='1';
          else
          cVar1S1S98P019P045P026P062(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='0' AND B(14)='1' )then
          cVar1S2S98P019N045P024P029(0) <='1';
          else
          cVar1S2S98P019N045P024P029(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='0' AND B(14)='1' )then
          cVar1S3S98P019N045P024P029(0) <='1';
          else
          cVar1S3S98P019N045P024P029(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='0' AND B(14)='0' )then
          cVar1S4S98P019N045P024N029(0) <='1';
          else
          cVar1S4S98P019N045P024N029(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='0' AND B(14)='0' )then
          cVar1S5S98P019N045P024N029(0) <='1';
          else
          cVar1S5S98P019N045P024N029(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='0' AND B(14)='0' )then
          cVar1S6S98P019N045P024N029(0) <='1';
          else
          cVar1S6S98P019N045P024N029(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(26)='1' AND A(19)='0' )then
          cVar1S7S98P019N045P024P001(0) <='1';
          else
          cVar1S7S98P019N045P024P001(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='1' AND A(21)='0' )then
          cVar1S8S98P019P051P025P016(0) <='1';
          else
          cVar1S8S98P019P051P025P016(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='1' AND A(21)='0' )then
          cVar1S9S98P019P051P025P016(0) <='1';
          else
          cVar1S9S98P019P051P025P016(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='1' AND A(21)='1' )then
          cVar1S10S98P019P051P025P016(0) <='1';
          else
          cVar1S10S98P019P051P025P016(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='0' AND B(14)='0' )then
          cVar1S11S98P019P051N025P029(0) <='1';
          else
          cVar1S11S98P019P051N025P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='0' AND B(14)='0' )then
          cVar1S12S98P019P051N025P029(0) <='1';
          else
          cVar1S12S98P019P051N025P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='0' AND B(14)='0' )then
          cVar1S13S98P019P051N025P029(0) <='1';
          else
          cVar1S13S98P019P051N025P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='0' AND B(14)='0' )then
          cVar1S14S98P019P051N025P029(0) <='1';
          else
          cVar1S14S98P019P051N025P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND B(16)='0' AND B(14)='1' )then
          cVar1S15S98P019P051N025P029(0) <='1';
          else
          cVar1S15S98P019P051N025P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='1' AND B(26)='0' )then
          cVar1S16S98P019P051P037P024(0) <='1';
          else
          cVar1S16S98P019P051P037P024(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='0' AND A(25)='1' )then
          cVar1S17S98P019P051N037P008(0) <='1';
          else
          cVar1S17S98P019P051N037P008(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='0' AND A(25)='0' )then
          cVar1S18S98P019P051N037N008(0) <='1';
          else
          cVar1S18S98P019P051N037N008(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='1' )then
          cVar1S0S99P045P030P025nsss(0) <='1';
          else
          cVar1S0S99P045P030P025nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='1' )then
          cVar1S1S99P045P030N025P022nsss(0) <='1';
          else
          cVar1S1S99P045P030N025P022nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S2S99P045P030N025N022(0) <='1';
          else
          cVar1S2S99P045P030N025N022(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S3S99P045P030N025N022(0) <='1';
          else
          cVar1S3S99P045P030N025N022(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND D(20)='0' )then
          cVar1S4S99N045P019P043P051(0) <='1';
          else
          cVar1S4S99N045P019P043P051(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND D(20)='0' )then
          cVar1S5S99N045P019P043P051(0) <='1';
          else
          cVar1S5S99N045P019P043P051(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND D(20)='0' )then
          cVar1S6S99N045P019P043P051(0) <='1';
          else
          cVar1S6S99N045P019P043P051(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND D(20)='1' )then
          cVar1S7S99N045P019P043P051(0) <='1';
          else
          cVar1S7S99N045P019P043P051(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND D(20)='1' )then
          cVar1S8S99N045P019P043P051(0) <='1';
          else
          cVar1S8S99N045P019P043P051(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='1' AND A(22)='0' )then
          cVar1S9S99N045P019P043P014(0) <='1';
          else
          cVar1S9S99N045P019P043P014(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='1' AND A(22)='0' )then
          cVar1S10S99N045P019P043P014(0) <='1';
          else
          cVar1S10S99N045P019P043P014(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S11S99N045N019P029P011(0) <='1';
          else
          cVar1S11S99N045N019P029P011(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S12S99N045N019P029P011(0) <='1';
          else
          cVar1S12S99N045N019P029P011(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S13S99N045N019P029P011(0) <='1';
          else
          cVar1S13S99N045N019P029P011(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S14S99N045N019P029N011(0) <='1';
          else
          cVar1S14S99N045N019P029N011(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S15S99N045N019P029N011(0) <='1';
          else
          cVar1S15S99N045N019P029N011(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND B(22)='1' )then
          cVar1S16S99N045N019N029P032(0) <='1';
          else
          cVar1S16S99N045N019N029P032(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND B(22)='1' )then
          cVar1S17S99N045N019N029P032(0) <='1';
          else
          cVar1S17S99N045N019N029P032(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND B(22)='0' )then
          cVar1S18S99N045N019N029N032(0) <='1';
          else
          cVar1S18S99N045N019N029N032(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND B(22)='0' )then
          cVar1S19S99N045N019N029N032(0) <='1';
          else
          cVar1S19S99N045N019N029N032(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S0S100P019P045P026P062(0) <='1';
          else
          cVar1S0S100P019P045P026P062(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND D( 9)='0' )then
          cVar1S1S100P019P045P026P062(0) <='1';
          else
          cVar1S1S100P019P045P026P062(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S2S100P019N045P029P011(0) <='1';
          else
          cVar1S2S100P019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S3S100P019N045P029P011(0) <='1';
          else
          cVar1S3S100P019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S4S100P019N045P029P011(0) <='1';
          else
          cVar1S4S100P019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S5S100P019N045P029N011(0) <='1';
          else
          cVar1S5S100P019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S6S100P019N045P029N011(0) <='1';
          else
          cVar1S6S100P019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND A(25)='0' )then
          cVar1S7S100P019N045N029P008(0) <='1';
          else
          cVar1S7S100P019N045N029P008(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND A(25)='0' )then
          cVar1S8S100P019N045N029P008(0) <='1';
          else
          cVar1S8S100P019N045N029P008(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND A(25)='0' )then
          cVar1S9S100P019N045N029P008(0) <='1';
          else
          cVar1S9S100P019N045N029P008(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND A(25)='1' )then
          cVar1S10S100P019N045N029P008(0) <='1';
          else
          cVar1S10S100P019N045N029P008(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND A(25)='1' )then
          cVar1S11S100P019N045N029P008(0) <='1';
          else
          cVar1S11S100P019N045N029P008(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='1' AND D(22)='1' )then
          cVar1S12S100P019P013P045P043nsss(0) <='1';
          else
          cVar1S12S100P019P013P045P043nsss(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='1' AND D(22)='0' )then
          cVar1S13S100P019P013P045N043(0) <='1';
          else
          cVar1S13S100P019P013P045N043(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='1' AND D(22)='0' )then
          cVar1S14S100P019P013P045N043(0) <='1';
          else
          cVar1S14S100P019P013P045N043(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='0' AND D(16)='1' )then
          cVar1S15S100P019P013N045P067(0) <='1';
          else
          cVar1S15S100P019P013N045P067(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='0' AND D(16)='1' )then
          cVar1S16S100P019P013N045P067(0) <='1';
          else
          cVar1S16S100P019P013N045P067(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='0' AND D(16)='0' )then
          cVar1S17S100P019P013N045N067(0) <='1';
          else
          cVar1S17S100P019P013N045N067(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='0' AND E(22)='0' AND D(16)='0' )then
          cVar1S18S100P019P013N045N067(0) <='1';
          else
          cVar1S18S100P019P013N045N067(0) <='0';
          end if;
        if(A(10)='1' AND A(13)='1' AND D(23)='0' AND E(23)='0' )then
          cVar1S19S100P019P013P039P041(0) <='1';
          else
          cVar1S19S100P019P013P039P041(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='1' )then
          cVar1S0S101P045P030P035P025nsss(0) <='1';
          else
          cVar1S0S101P045P030P035P025nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='0' )then
          cVar1S1S101P045P030P035N025(0) <='1';
          else
          cVar1S1S101P045P030P035N025(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='0' )then
          cVar1S2S101P045P030P035N025(0) <='1';
          else
          cVar1S2S101P045P030P035N025(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='0' )then
          cVar1S3S101P045P030P035N025(0) <='1';
          else
          cVar1S3S101P045P030P035N025(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND B(17)='0' )then
          cVar1S4S101N045P019P043P023(0) <='1';
          else
          cVar1S4S101N045P019P043P023(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND B(17)='0' )then
          cVar1S5S101N045P019P043P023(0) <='1';
          else
          cVar1S5S101N045P019P043P023(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND B(17)='0' )then
          cVar1S6S101N045P019P043P023(0) <='1';
          else
          cVar1S6S101N045P019P043P023(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='0' AND B(17)='1' )then
          cVar1S7S101N045P019P043P023(0) <='1';
          else
          cVar1S7S101N045P019P043P023(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='1' AND A(22)='0' )then
          cVar1S8S101N045P019P043P014(0) <='1';
          else
          cVar1S8S101N045P019P043P014(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='1' AND D(22)='1' AND A(22)='0' )then
          cVar1S9S101N045P019P043P014(0) <='1';
          else
          cVar1S9S101N045P019P043P014(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND B(26)='0' )then
          cVar1S10S101N045N019P029P024(0) <='1';
          else
          cVar1S10S101N045N019P029P024(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='1' AND B(26)='0' )then
          cVar1S11S101N045N019P029P024(0) <='1';
          else
          cVar1S11S101N045N019P029P024(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND E(15)='1' )then
          cVar1S12S101N045N019N029P040(0) <='1';
          else
          cVar1S12S101N045N019N029P040(0) <='0';
          end if;
        if(E(22)='0' AND A(10)='0' AND B(14)='0' AND E(15)='1' )then
          cVar1S13S101N045N019N029P040(0) <='1';
          else
          cVar1S13S101N045N019N029P040(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND A(17)='1' )then
          cVar1S0S102P019P045P026P005nsss(0) <='1';
          else
          cVar1S0S102P019P045P026P005nsss(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND A(17)='0' )then
          cVar1S1S102P019P045P026N005(0) <='1';
          else
          cVar1S1S102P019P045P026N005(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND E(18)='0' )then
          cVar1S2S102P019N045P029P061(0) <='1';
          else
          cVar1S2S102P019N045P029P061(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND E(18)='0' )then
          cVar1S3S102P019N045P029P061(0) <='1';
          else
          cVar1S3S102P019N045P029P061(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S4S102P019N045N029P054(0) <='1';
          else
          cVar1S4S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S5S102P019N045N029P054(0) <='1';
          else
          cVar1S5S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S6S102P019N045N029P054(0) <='1';
          else
          cVar1S6S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='0' )then
          cVar1S7S102P019N045N029P054(0) <='1';
          else
          cVar1S7S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S8S102P019N045N029P054(0) <='1';
          else
          cVar1S8S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S9S102P019N045N029P054(0) <='1';
          else
          cVar1S9S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND D(11)='1' )then
          cVar1S10S102P019N045N029P054(0) <='1';
          else
          cVar1S10S102P019N045N029P054(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='1' AND E(19)='0' )then
          cVar1S11S102P019P051P018P057(0) <='1';
          else
          cVar1S11S102P019P051P018P057(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='1' AND E(19)='0' )then
          cVar1S12S102P019P051P018P057(0) <='1';
          else
          cVar1S12S102P019P051P018P057(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='1' AND E(19)='0' )then
          cVar1S13S102P019P051P018P057(0) <='1';
          else
          cVar1S13S102P019P051P018P057(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='1' AND E(19)='1' )then
          cVar1S14S102P019P051P018P057(0) <='1';
          else
          cVar1S14S102P019P051P018P057(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='0' AND E(20)='0' )then
          cVar1S15S102P019P051N018P053(0) <='1';
          else
          cVar1S15S102P019P051N018P053(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='0' AND E(20)='0' )then
          cVar1S16S102P019P051N018P053(0) <='1';
          else
          cVar1S16S102P019P051N018P053(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='0' AND E(20)='0' )then
          cVar1S17S102P019P051N018P053(0) <='1';
          else
          cVar1S17S102P019P051N018P053(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND A(20)='0' AND E(20)='1' )then
          cVar1S18S102P019P051N018P053(0) <='1';
          else
          cVar1S18S102P019P051N018P053(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(26)='0' AND B(10)='1' )then
          cVar1S19S102P019P051P024P037(0) <='1';
          else
          cVar1S19S102P019P051P024P037(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(26)='0' AND B(10)='0' )then
          cVar1S20S102P019P051P024N037(0) <='1';
          else
          cVar1S20S102P019P051P024N037(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='1' )then
          cVar1S0S103P045P030P025nsss(0) <='1';
          else
          cVar1S0S103P045P030P025nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='1' )then
          cVar1S1S103P045P030N025P022nsss(0) <='1';
          else
          cVar1S1S103P045P030N025P022nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S2S103P045P030N025N022(0) <='1';
          else
          cVar1S2S103P045P030N025N022(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(16)='0' AND B(27)='0' )then
          cVar1S3S103P045P030N025N022(0) <='1';
          else
          cVar1S3S103P045P030N025N022(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='1' AND E(17)='1' )then
          cVar1S4S103N045P052P065nsss(0) <='1';
          else
          cVar1S4S103N045P052P065nsss(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='1' )then
          cVar1S5S103N045P052N065P062nsss(0) <='1';
          else
          cVar1S5S103N045P052N065P062nsss(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S6S103N045P052N065N062(0) <='1';
          else
          cVar1S6S103N045P052N065N062(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='1' AND E(17)='0' AND D( 9)='0' )then
          cVar1S7S103N045P052N065N062(0) <='1';
          else
          cVar1S7S103N045P052N065N062(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='0' AND A(20)='0' )then
          cVar1S8S103N045N052P043P018(0) <='1';
          else
          cVar1S8S103N045N052P043P018(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='0' AND A(20)='0' )then
          cVar1S9S103N045N052P043P018(0) <='1';
          else
          cVar1S9S103N045N052P043P018(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='0' AND A(20)='1' )then
          cVar1S10S103N045N052P043P018(0) <='1';
          else
          cVar1S10S103N045N052P043P018(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='0' AND A(20)='1' )then
          cVar1S11S103N045N052P043P018(0) <='1';
          else
          cVar1S11S103N045N052P043P018(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='0' AND A(20)='1' )then
          cVar1S12S103N045N052P043P018(0) <='1';
          else
          cVar1S12S103N045N052P043P018(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='1' AND D(17)='0' )then
          cVar1S13S103N045N052P043P063(0) <='1';
          else
          cVar1S13S103N045N052P043P063(0) <='0';
          end if;
        if(E(22)='0' AND E(12)='0' AND D(22)='1' AND D(17)='0' )then
          cVar1S14S103N045N052P043P063(0) <='1';
          else
          cVar1S14S103N045N052P043P063(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND A(17)='1' )then
          cVar1S0S104P019P045P026P005nsss(0) <='1';
          else
          cVar1S0S104P019P045P026P005nsss(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='1' AND B(25)='0' AND A(17)='0' )then
          cVar1S1S104P019P045P026N005(0) <='1';
          else
          cVar1S1S104P019P045P026N005(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S2S104P019N045P029P011(0) <='1';
          else
          cVar1S2S104P019N045P029P011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S3S104P019N045P029N011(0) <='1';
          else
          cVar1S3S104P019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S4S104P019N045P029N011(0) <='1';
          else
          cVar1S4S104P019N045P029N011(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND E(16)='0' )then
          cVar1S5S104P019N045N029P069(0) <='1';
          else
          cVar1S5S104P019N045N029P069(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND E(16)='0' )then
          cVar1S6S104P019N045N029P069(0) <='1';
          else
          cVar1S6S104P019N045N029P069(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND E(16)='0' )then
          cVar1S7S104P019N045N029P069(0) <='1';
          else
          cVar1S7S104P019N045N029P069(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND E(16)='1' )then
          cVar1S8S104P019N045N029P069(0) <='1';
          else
          cVar1S8S104P019N045N029P069(0) <='0';
          end if;
        if(A(10)='0' AND E(22)='0' AND B(14)='0' AND E(16)='1' )then
          cVar1S9S104P019N045N029P069(0) <='1';
          else
          cVar1S9S104P019N045N029P069(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='1' AND A(26)='1' )then
          cVar1S10S104P019P067P047P006nsss(0) <='1';
          else
          cVar1S10S104P019P067P047P006nsss(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='1' AND A(26)='0' )then
          cVar1S11S104P019P067P047N006(0) <='1';
          else
          cVar1S11S104P019P067P047N006(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='1' AND A(26)='0' )then
          cVar1S12S104P019P067P047N006(0) <='1';
          else
          cVar1S12S104P019P067P047N006(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='0' AND E(16)='0' )then
          cVar1S13S104P019P067N047P069(0) <='1';
          else
          cVar1S13S104P019P067N047P069(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='0' AND E(16)='0' )then
          cVar1S14S104P019P067N047P069(0) <='1';
          else
          cVar1S14S104P019P067N047P069(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='0' AND E(16)='1' )then
          cVar1S15S104P019P067N047P069(0) <='1';
          else
          cVar1S15S104P019P067N047P069(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='0' AND D(21)='0' AND E(16)='1' )then
          cVar1S16S104P019P067N047P069(0) <='1';
          else
          cVar1S16S104P019P067N047P069(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='1' AND B(26)='0' AND D(14)='1' )then
          cVar1S17S104P019P067P024P042nsss(0) <='1';
          else
          cVar1S17S104P019P067P024P042nsss(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='1' AND B(26)='0' AND D(14)='0' )then
          cVar1S18S104P019P067P024N042(0) <='1';
          else
          cVar1S18S104P019P067P024N042(0) <='0';
          end if;
        if(A(10)='1' AND D(16)='1' AND B(26)='1' AND E(16)='1' )then
          cVar1S19S104P019P067P024P069(0) <='1';
          else
          cVar1S19S104P019P067P024P069(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='1' )then
          cVar1S0S105P045P030P035P025nsss(0) <='1';
          else
          cVar1S0S105P045P030P035P025nsss(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='0' )then
          cVar1S1S105P045P030P035N025(0) <='1';
          else
          cVar1S1S105P045P030P035N025(0) <='0';
          end if;
        if(E(22)='1' AND B(23)='0' AND B(11)='0' AND B(16)='0' )then
          cVar1S2S105P045P030P035N025(0) <='1';
          else
          cVar1S2S105P045P030P035N025(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='1' AND D(18)='0' AND B(24)='0' )then
          cVar1S3S105N045P029P059P028(0) <='1';
          else
          cVar1S3S105N045P029P059P028(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='1' AND D(18)='0' AND B(24)='0' )then
          cVar1S4S105N045P029P059P028(0) <='1';
          else
          cVar1S4S105N045P029P059P028(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='0' AND D( 9)='1' )then
          cVar1S5S105N045N029P043P062(0) <='1';
          else
          cVar1S5S105N045N029P043P062(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='0' AND D( 9)='1' )then
          cVar1S6S105N045N029P043P062(0) <='1';
          else
          cVar1S6S105N045N029P043P062(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='0' AND D( 9)='0' )then
          cVar1S7S105N045N029P043N062(0) <='1';
          else
          cVar1S7S105N045N029P043N062(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='0' AND D( 9)='0' )then
          cVar1S8S105N045N029P043N062(0) <='1';
          else
          cVar1S8S105N045N029P043N062(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='0' AND D( 9)='0' )then
          cVar1S9S105N045N029P043N062(0) <='1';
          else
          cVar1S9S105N045N029P043N062(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='1' AND B(27)='1' )then
          cVar1S10S105N045N029P043P022nsss(0) <='1';
          else
          cVar1S10S105N045N029P043P022nsss(0) <='0';
          end if;
        if(E(22)='0' AND B(14)='0' AND D(22)='1' AND B(27)='0' )then
          cVar1S11S105N045N029P043N022(0) <='1';
          else
          cVar1S11S105N045N029P043N022(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='0' )then
          cVar1S0S106P020P039P041P002(0) <='1';
          else
          cVar1S0S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='0' )then
          cVar1S1S106P020P039P041P002(0) <='1';
          else
          cVar1S1S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='0' )then
          cVar1S2S106P020P039P041P002(0) <='1';
          else
          cVar1S2S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='0' )then
          cVar1S3S106P020P039P041P002(0) <='1';
          else
          cVar1S3S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='1' )then
          cVar1S4S106P020P039P041P002(0) <='1';
          else
          cVar1S4S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='1' )then
          cVar1S5S106P020P039P041P002(0) <='1';
          else
          cVar1S5S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='0' AND A(28)='1' )then
          cVar1S6S106P020P039P041P002(0) <='1';
          else
          cVar1S6S106P020P039P041P002(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='0' AND E(23)='1' AND B(12)='1' )then
          cVar1S7S106P020P039P041P033nsss(0) <='1';
          else
          cVar1S7S106P020P039P041P033nsss(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='1' AND A(23)='0' AND E(10)='0' )then
          cVar1S8S106P020P039P012P060(0) <='1';
          else
          cVar1S8S106P020P039P012P060(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='1' AND A(23)='0' AND E(10)='0' )then
          cVar1S9S106P020P039P012P060(0) <='1';
          else
          cVar1S9S106P020P039P012P060(0) <='0';
          end if;
        if(B(28)='0' AND D(23)='1' AND A(23)='0' AND E(10)='0' )then
          cVar1S10S106P020P039P012P060(0) <='1';
          else
          cVar1S10S106P020P039P012P060(0) <='0';
          end if;
        if(B(28)='1' AND D(23)='1' AND E(23)='1' )then
          cVar1S11S106P020P039P041nsss(0) <='1';
          else
          cVar1S11S106P020P039P041nsss(0) <='0';
          end if;
        if(B(28)='1' AND D(23)='0' AND A(29)='0' AND A(11)='1' )then
          cVar1S12S106P020N039P000P017(0) <='1';
          else
          cVar1S12S106P020N039P000P017(0) <='0';
          end if;
        if(B(28)='1' AND D(23)='0' AND A(29)='0' AND A(11)='1' )then
          cVar1S13S106P020N039P000P017(0) <='1';
          else
          cVar1S13S106P020N039P000P017(0) <='0';
          end if;
        if(B(28)='1' AND D(23)='0' AND A(29)='0' AND A(11)='0' )then
          cVar1S14S106P020N039P000N017(0) <='1';
          else
          cVar1S14S106P020N039P000N017(0) <='0';
          end if;
        if(D(20)='1' AND E(23)='0' AND B(26)='0' AND E(20)='1' )then
          cVar1S0S107P051P041P024P053(0) <='1';
          else
          cVar1S0S107P051P041P024P053(0) <='0';
          end if;
        if(D(20)='1' AND E(23)='0' AND B(26)='0' AND E(20)='0' )then
          cVar1S1S107P051P041P024N053(0) <='1';
          else
          cVar1S1S107P051P041P024N053(0) <='0';
          end if;
        if(D(20)='1' AND E(23)='0' AND B(26)='0' AND E(20)='0' )then
          cVar1S2S107P051P041P024N053(0) <='1';
          else
          cVar1S2S107P051P041P024N053(0) <='0';
          end if;
        if(D(20)='1' AND E(23)='0' AND B(26)='1' AND D(16)='0' )then
          cVar1S3S107P051P041P024P067(0) <='1';
          else
          cVar1S3S107P051P041P024P067(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='1' AND B(16)='1' )then
          cVar1S4S107N051P053P007P025nsss(0) <='1';
          else
          cVar1S4S107N051P053P007P025nsss(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='1' AND B(16)='0' )then
          cVar1S5S107N051P053P007N025(0) <='1';
          else
          cVar1S5S107N051P053P007N025(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='1' AND B(16)='0' )then
          cVar1S6S107N051P053P007N025(0) <='1';
          else
          cVar1S6S107N051P053P007N025(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='1' AND B(16)='0' )then
          cVar1S7S107N051P053P007N025(0) <='1';
          else
          cVar1S7S107N051P053P007N025(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='0' AND E(13)='0' )then
          cVar1S8S107N051P053N007P048(0) <='1';
          else
          cVar1S8S107N051P053N007P048(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='0' AND E(13)='0' )then
          cVar1S9S107N051P053N007P048(0) <='1';
          else
          cVar1S9S107N051P053N007P048(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='0' AND A(16)='0' AND E(13)='1' )then
          cVar1S10S107N051P053N007P048(0) <='1';
          else
          cVar1S10S107N051P053N007P048(0) <='0';
          end if;
        if(D(20)='0' AND E(20)='1' AND B(15)='0' AND B(23)='0' )then
          cVar1S11S107N051P053P027P030(0) <='1';
          else
          cVar1S11S107N051P053P027P030(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='1' AND D(23)='0' )then
          cVar1S0S108P061P059P051P039(0) <='1';
          else
          cVar1S0S108P061P059P051P039(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='1' AND D(23)='0' )then
          cVar1S1S108P061P059P051P039(0) <='1';
          else
          cVar1S1S108P061P059P051P039(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='1' )then
          cVar1S2S108P061P059N051P045(0) <='1';
          else
          cVar1S2S108P061P059N051P045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='1' )then
          cVar1S3S108P061P059N051P045(0) <='1';
          else
          cVar1S3S108P061P059N051P045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='1' )then
          cVar1S4S108P061P059N051P045(0) <='1';
          else
          cVar1S4S108P061P059N051P045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='0' )then
          cVar1S5S108P061P059N051N045(0) <='1';
          else
          cVar1S5S108P061P059N051N045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='0' )then
          cVar1S6S108P061P059N051N045(0) <='1';
          else
          cVar1S6S108P061P059N051N045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='0' )then
          cVar1S7S108P061P059N051N045(0) <='1';
          else
          cVar1S7S108P061P059N051N045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='0' AND D(20)='0' AND E(22)='0' )then
          cVar1S8S108P061P059N051N045(0) <='1';
          else
          cVar1S8S108P061P059N051N045(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='1' AND E(12)='0' AND D( 9)='0' )then
          cVar1S9S108P061P059P052P062(0) <='1';
          else
          cVar1S9S108P061P059P052P062(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='1' AND E(12)='0' AND D( 9)='0' )then
          cVar1S10S108P061P059P052P062(0) <='1';
          else
          cVar1S10S108P061P059P052P062(0) <='0';
          end if;
        if(E(18)='0' AND D(18)='1' AND E(12)='0' AND D( 9)='0' )then
          cVar1S11S108P061P059P052P062(0) <='1';
          else
          cVar1S11S108P061P059P052P062(0) <='0';
          end if;
        if(E(18)='1' AND E(15)='0' AND B(12)='1' AND A(12)='1' )then
          cVar1S12S108P061P040P033P015(0) <='1';
          else
          cVar1S12S108P061P040P033P015(0) <='0';
          end if;
        if(E(18)='1' AND E(15)='0' AND B(12)='1' AND A(12)='0' )then
          cVar1S13S108P061P040P033N015(0) <='1';
          else
          cVar1S13S108P061P040P033N015(0) <='0';
          end if;
        if(E(18)='1' AND E(15)='0' AND B(12)='0' AND E(23)='0' )then
          cVar1S14S108P061P040N033P041(0) <='1';
          else
          cVar1S14S108P061P040N033P041(0) <='0';
          end if;
        if(E(18)='1' AND E(15)='0' AND B(12)='0' AND E(23)='0' )then
          cVar1S15S108P061P040N033P041(0) <='1';
          else
          cVar1S15S108P061P040N033P041(0) <='0';
          end if;
        if(E(18)='1' AND E(15)='0' AND B(12)='0' AND E(23)='0' )then
          cVar1S16S108P061P040N033P041(0) <='1';
          else
          cVar1S16S108P061P040N033P041(0) <='0';
          end if;
        if(B(27)='1' AND D(22)='1' )then
          cVar1S0S109P022P043nsss(0) <='1';
          else
          cVar1S0S109P022P043nsss(0) <='0';
          end if;
        if(B(27)='1' AND D(22)='0' AND A(28)='1' )then
          cVar1S1S109P022N043P002nsss(0) <='1';
          else
          cVar1S1S109P022N043P002nsss(0) <='0';
          end if;
        if(B(27)='1' AND D(22)='0' AND A(28)='0' AND A(18)='0' )then
          cVar1S2S109P022N043N002P003(0) <='1';
          else
          cVar1S2S109P022N043N002P003(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='0' AND A(29)='0' AND E(11)='1' )then
          cVar1S3S109N022P043P000P056(0) <='1';
          else
          cVar1S3S109N022P043P000P056(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='0' AND A(29)='0' AND E(11)='1' )then
          cVar1S4S109N022P043P000P056(0) <='1';
          else
          cVar1S4S109N022P043P000P056(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='0' AND A(29)='0' AND E(11)='0' )then
          cVar1S5S109N022P043P000N056(0) <='1';
          else
          cVar1S5S109N022P043P000N056(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='0' AND A(29)='0' AND E(11)='0' )then
          cVar1S6S109N022P043P000N056(0) <='1';
          else
          cVar1S6S109N022P043P000N056(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='1' AND B(16)='1' )then
          cVar1S7S109N022P043P025nsss(0) <='1';
          else
          cVar1S7S109N022P043P025nsss(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='1' AND B(16)='0' AND D(12)='0' )then
          cVar1S8S109N022P043N025P050(0) <='1';
          else
          cVar1S8S109N022P043N025P050(0) <='0';
          end if;
        if(B(27)='0' AND D(22)='1' AND B(16)='0' AND D(12)='0' )then
          cVar1S9S109N022P043N025P050(0) <='1';
          else
          cVar1S9S109N022P043N025P050(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='1' AND E(23)='0' AND E(20)='1' )then
          cVar1S0S110P000P051P041P053(0) <='1';
          else
          cVar1S0S110P000P051P041P053(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='1' AND E(23)='0' AND E(20)='1' )then
          cVar1S1S110P000P051P041P053(0) <='1';
          else
          cVar1S1S110P000P051P041P053(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='1' AND E(23)='0' AND E(20)='1' )then
          cVar1S2S110P000P051P041P053(0) <='1';
          else
          cVar1S2S110P000P051P041P053(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='1' AND E(23)='0' AND E(20)='0' )then
          cVar1S3S110P000P051P041N053(0) <='1';
          else
          cVar1S3S110P000P051P041N053(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='1' AND E(23)='0' AND E(20)='0' )then
          cVar1S4S110P000P051P041N053(0) <='1';
          else
          cVar1S4S110P000P051P041N053(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='0' AND E(14)='1' )then
          cVar1S5S110P000N051P053P044(0) <='1';
          else
          cVar1S5S110P000N051P053P044(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='0' AND E(14)='1' )then
          cVar1S6S110P000N051P053P044(0) <='1';
          else
          cVar1S6S110P000N051P053P044(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='0' AND E(14)='0' )then
          cVar1S7S110P000N051P053N044(0) <='1';
          else
          cVar1S7S110P000N051P053N044(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='0' AND E(14)='0' )then
          cVar1S8S110P000N051P053N044(0) <='1';
          else
          cVar1S8S110P000N051P053N044(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='0' AND E(14)='0' )then
          cVar1S9S110P000N051P053N044(0) <='1';
          else
          cVar1S9S110P000N051P053N044(0) <='0';
          end if;
        if(A(29)='0' AND D(20)='0' AND E(20)='1' AND B(23)='0' )then
          cVar1S10S110P000N051P053P030(0) <='1';
          else
          cVar1S10S110P000N051P053P030(0) <='0';
          end if;
        if(A(29)='1' AND B(23)='0' AND B(15)='0' AND E(10)='0' )then
          cVar1S11S110P000P030P027P060(0) <='1';
          else
          cVar1S11S110P000P030P027P060(0) <='0';
          end if;
        if(E(20)='1' AND A(27)='0' AND D(20)='1' AND A(29)='0' )then
          cVar1S0S111P053P004P051P000(0) <='1';
          else
          cVar1S0S111P053P004P051P000(0) <='0';
          end if;
        if(E(20)='1' AND A(27)='0' AND D(20)='1' AND A(29)='0' )then
          cVar1S1S111P053P004P051P000(0) <='1';
          else
          cVar1S1S111P053P004P051P000(0) <='0';
          end if;
        if(E(20)='1' AND A(27)='0' AND D(20)='1' AND A(29)='0' )then
          cVar1S2S111P053P004P051P000(0) <='1';
          else
          cVar1S2S111P053P004P051P000(0) <='0';
          end if;
        if(E(20)='1' AND A(27)='0' AND D(20)='0' AND B(23)='0' )then
          cVar1S3S111P053P004N051P030(0) <='1';
          else
          cVar1S3S111P053P004N051P030(0) <='0';
          end if;
        if(E(20)='1' AND A(27)='0' AND D(20)='0' AND B(23)='0' )then
          cVar1S4S111P053P004N051P030(0) <='1';
          else
          cVar1S4S111P053P004N051P030(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='1' AND B(16)='1' )then
          cVar1S5S111N053P044P025nsss(0) <='1';
          else
          cVar1S5S111N053P044P025nsss(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S6S111N053P044N025P023nsss(0) <='1';
          else
          cVar1S6S111N053P044N025P023nsss(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='1' AND B(16)='0' AND B(17)='0' )then
          cVar1S7S111N053P044N025N023(0) <='1';
          else
          cVar1S7S111N053P044N025N023(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='0' AND B(17)='0' )then
          cVar1S8S111N053N044P042P023(0) <='1';
          else
          cVar1S8S111N053N044P042P023(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='0' AND B(17)='0' )then
          cVar1S9S111N053N044P042P023(0) <='1';
          else
          cVar1S9S111N053N044P042P023(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='0' AND B(17)='1' )then
          cVar1S10S111N053N044P042P023(0) <='1';
          else
          cVar1S10S111N053N044P042P023(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='0' AND B(17)='1' )then
          cVar1S11S111N053N044P042P023(0) <='1';
          else
          cVar1S11S111N053N044P042P023(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='1' AND A(17)='1' )then
          cVar1S12S111N053N044P042P005nsss(0) <='1';
          else
          cVar1S12S111N053N044P042P005nsss(0) <='0';
          end if;
        if(E(20)='0' AND E(14)='0' AND D(14)='1' AND A(17)='0' )then
          cVar1S13S111N053N044P042N005(0) <='1';
          else
          cVar1S13S111N053N044P042N005(0) <='0';
          end if;
        if(E(14)='1' AND B(17)='1' )then
          cVar1S0S112P044P023nsss(0) <='1';
          else
          cVar1S0S112P044P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S112P044N023P025nsss(0) <='1';
          else
          cVar1S1S112P044N023P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(17)='0' AND B(16)='0' AND B(22)='0' )then
          cVar1S2S112P044N023N025P032(0) <='1';
          else
          cVar1S2S112P044N023N025P032(0) <='0';
          end if;
        if(E(14)='1' AND B(17)='0' AND B(16)='0' AND B(22)='0' )then
          cVar1S3S112P044N023N025P032(0) <='1';
          else
          cVar1S3S112P044N023N025P032(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='1' )then
          cVar1S4S112N044P042P023P051(0) <='1';
          else
          cVar1S4S112N044P042P023P051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='1' )then
          cVar1S5S112N044P042P023P051(0) <='1';
          else
          cVar1S5S112N044P042P023P051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='0' )then
          cVar1S6S112N044P042P023N051(0) <='1';
          else
          cVar1S6S112N044P042P023N051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='0' )then
          cVar1S7S112N044P042P023N051(0) <='1';
          else
          cVar1S7S112N044P042P023N051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S8S112N044P042P023P024(0) <='1';
          else
          cVar1S8S112N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S9S112N044P042P023P024(0) <='1';
          else
          cVar1S9S112N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND D( 9)='0' )then
          cVar1S10S112N044P042P024P062(0) <='1';
          else
          cVar1S10S112N044P042P024P062(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND D( 9)='0' )then
          cVar1S11S112N044P042P024P062(0) <='1';
          else
          cVar1S11S112N044P042P024P062(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S113P044P025nsss(0) <='1';
          else
          cVar1S0S113P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S113P044N025P023nsss(0) <='1';
          else
          cVar1S1S113P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND B(22)='0' )then
          cVar1S2S113P044N025N023P032(0) <='1';
          else
          cVar1S2S113P044N025N023P032(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='1' )then
          cVar1S3S113N044P042P023P051(0) <='1';
          else
          cVar1S3S113N044P042P023P051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='1' )then
          cVar1S4S113N044P042P023P051(0) <='1';
          else
          cVar1S4S113N044P042P023P051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='0' )then
          cVar1S5S113N044P042P023N051(0) <='1';
          else
          cVar1S5S113N044P042P023N051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='0' )then
          cVar1S6S113N044P042P023N051(0) <='1';
          else
          cVar1S6S113N044P042P023N051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND D(20)='0' )then
          cVar1S7S113N044P042P023N051(0) <='1';
          else
          cVar1S7S113N044P042P023N051(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S8S113N044P042P023P024(0) <='1';
          else
          cVar1S8S113N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S9S113N044P042P023P024(0) <='1';
          else
          cVar1S9S113N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND D( 9)='0' )then
          cVar1S10S113N044P042P024P062(0) <='1';
          else
          cVar1S10S113N044P042P024P062(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND D( 9)='0' )then
          cVar1S11S113N044P042P024P062(0) <='1';
          else
          cVar1S11S113N044P042P024P062(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='1' )then
          cVar1S0S114P016P044P023nsss(0) <='1';
          else
          cVar1S0S114P016P044P023nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S114P016P044N023P025nsss(0) <='1';
          else
          cVar1S1S114P016P044N023P025nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S2S114P016P044N023N025(0) <='1';
          else
          cVar1S2S114P016P044N023N025(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='1' AND B(28)='1' )then
          cVar1S3S114P016N044P041P020nsss(0) <='1';
          else
          cVar1S3S114P016N044P041P020nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='1' AND B(28)='0' )then
          cVar1S4S114P016N044P041N020(0) <='1';
          else
          cVar1S4S114P016N044P041N020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND B(28)='0' )then
          cVar1S5S114P016N044N041P020(0) <='1';
          else
          cVar1S5S114P016N044N041P020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND B(28)='0' )then
          cVar1S6S114P016N044N041P020(0) <='1';
          else
          cVar1S6S114P016N044N041P020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND B(28)='0' )then
          cVar1S7S114P016N044N041P020(0) <='1';
          else
          cVar1S7S114P016N044N041P020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND B(28)='1' )then
          cVar1S8S114P016N044N041P020(0) <='1';
          else
          cVar1S8S114P016N044N041P020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND B(28)='1' )then
          cVar1S9S114P016N044N041P020(0) <='1';
          else
          cVar1S9S114P016N044N041P020(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='0' )then
          cVar1S10S114P016P039P022P041(0) <='1';
          else
          cVar1S10S114P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='0' )then
          cVar1S11S114P016P039P022P041(0) <='1';
          else
          cVar1S11S114P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='0' )then
          cVar1S12S114P016P039P022P041(0) <='1';
          else
          cVar1S12S114P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='0' AND E(23)='1' )then
          cVar1S13S114P016P039P022P041(0) <='1';
          else
          cVar1S13S114P016P039P022P041(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND B(27)='1' AND A(10)='1' )then
          cVar1S14S114P016P039P022P019(0) <='1';
          else
          cVar1S14S114P016P039P022P019(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(17)='1' )then
          cVar1S15S114P016P039P005nsss(0) <='1';
          else
          cVar1S15S114P016P039P005nsss(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(17)='0' AND E(16)='0' )then
          cVar1S16S114P016P039N005P069(0) <='1';
          else
          cVar1S16S114P016P039N005P069(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S115P044P025nsss(0) <='1';
          else
          cVar1S0S115P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S115P044N025P023nsss(0) <='1';
          else
          cVar1S1S115P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND B(22)='0' )then
          cVar1S2S115P044N025N023P032(0) <='1';
          else
          cVar1S2S115P044N025N023P032(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='1' )then
          cVar1S3S115N044P042P023P008(0) <='1';
          else
          cVar1S3S115N044P042P023P008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='1' )then
          cVar1S4S115N044P042P023P008(0) <='1';
          else
          cVar1S4S115N044P042P023P008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='1' )then
          cVar1S5S115N044P042P023P008(0) <='1';
          else
          cVar1S5S115N044P042P023P008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='0' )then
          cVar1S6S115N044P042P023N008(0) <='1';
          else
          cVar1S6S115N044P042P023N008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='0' )then
          cVar1S7S115N044P042P023N008(0) <='1';
          else
          cVar1S7S115N044P042P023N008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='0' AND A(25)='0' )then
          cVar1S8S115N044P042P023N008(0) <='1';
          else
          cVar1S8S115N044P042P023N008(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S9S115N044P042P023P024(0) <='1';
          else
          cVar1S9S115N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S10S115N044P042P023P024(0) <='1';
          else
          cVar1S10S115N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='0' AND B(17)='1' AND B(26)='0' )then
          cVar1S11S115N044P042P023P024(0) <='1';
          else
          cVar1S11S115N044P042P023P024(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND A(17)='1' )then
          cVar1S12S115N044P042P024P005nsss(0) <='1';
          else
          cVar1S12S115N044P042P024P005nsss(0) <='0';
          end if;
        if(E(14)='0' AND D(14)='1' AND B(26)='0' AND A(17)='0' )then
          cVar1S13S115N044P042P024N005(0) <='1';
          else
          cVar1S13S115N044P042P024N005(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='1' )then
          cVar1S0S116P016P044P023nsss(0) <='1';
          else
          cVar1S0S116P016P044P023nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='0' AND B(16)='1' )then
          cVar1S1S116P016P044N023P025nsss(0) <='1';
          else
          cVar1S1S116P016P044N023P025nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='1' AND B(17)='0' AND B(16)='0' )then
          cVar1S2S116P016P044N023N025(0) <='1';
          else
          cVar1S2S116P016P044N023N025(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='1' AND B(28)='1' )then
          cVar1S3S116P016N044P041P020nsss(0) <='1';
          else
          cVar1S3S116P016N044P041P020nsss(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='1' AND B(28)='0' )then
          cVar1S4S116P016N044P041N020(0) <='1';
          else
          cVar1S4S116P016N044P041N020(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND A(27)='0' )then
          cVar1S5S116P016N044N041P004(0) <='1';
          else
          cVar1S5S116P016N044N041P004(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND A(27)='0' )then
          cVar1S6S116P016N044N041P004(0) <='1';
          else
          cVar1S6S116P016N044N041P004(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND A(27)='0' )then
          cVar1S7S116P016N044N041P004(0) <='1';
          else
          cVar1S7S116P016N044N041P004(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND A(27)='0' )then
          cVar1S8S116P016N044N041P004(0) <='1';
          else
          cVar1S8S116P016N044N041P004(0) <='0';
          end if;
        if(A(21)='0' AND E(14)='0' AND E(23)='0' AND A(27)='1' )then
          cVar1S9S116P016N044N041P004(0) <='1';
          else
          cVar1S9S116P016N044N041P004(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='0' )then
          cVar1S10S116P016P039P041P022(0) <='1';
          else
          cVar1S10S116P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='0' )then
          cVar1S11S116P016P039P041P022(0) <='1';
          else
          cVar1S11S116P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='0' )then
          cVar1S12S116P016P039P041P022(0) <='1';
          else
          cVar1S12S116P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='0' AND B(27)='1' )then
          cVar1S13S116P016P039P041P022(0) <='1';
          else
          cVar1S13S116P016P039P041P022(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='0' AND E(23)='1' AND E(16)='0' )then
          cVar1S14S116P016P039P041P069(0) <='1';
          else
          cVar1S14S116P016P039P041P069(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(17)='1' )then
          cVar1S15S116P016P039P005nsss(0) <='1';
          else
          cVar1S15S116P016P039P005nsss(0) <='0';
          end if;
        if(A(21)='1' AND D(23)='1' AND A(17)='0' AND E(16)='0' )then
          cVar1S16S116P016P039N005P069(0) <='1';
          else
          cVar1S16S116P016P039N005P069(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S117P044P025nsss(0) <='1';
          else
          cVar1S0S117P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S117P044N025P023nsss(0) <='1';
          else
          cVar1S1S117P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND B(22)='0' )then
          cVar1S2S117P044N025N023P032(0) <='1';
          else
          cVar1S2S117P044N025N023P032(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S3S117N044P023P042P002(0) <='1';
          else
          cVar1S3S117N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S4S117N044P023P042P002(0) <='1';
          else
          cVar1S4S117N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S5S117N044P023P042P002(0) <='1';
          else
          cVar1S5S117N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='1' )then
          cVar1S6S117N044P023P042P002(0) <='1';
          else
          cVar1S6S117N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='1' )then
          cVar1S7S117N044P023P042P002(0) <='1';
          else
          cVar1S7S117N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S8S117N044P023P042P024(0) <='1';
          else
          cVar1S8S117N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S9S117N044P023P042P024(0) <='1';
          else
          cVar1S9S117N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S10S117N044P023P042P024(0) <='1';
          else
          cVar1S10S117N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='1' )then
          cVar1S11S117N044P023P024P005nsss(0) <='1';
          else
          cVar1S11S117N044P023P024P005nsss(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='0' )then
          cVar1S12S117N044P023P024N005(0) <='1';
          else
          cVar1S12S117N044P023P024N005(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S118P044P025nsss(0) <='1';
          else
          cVar1S0S118P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S118P044N025P023nsss(0) <='1';
          else
          cVar1S1S118P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND B(22)='0' )then
          cVar1S2S118P044N025N023P032(0) <='1';
          else
          cVar1S2S118P044N025N023P032(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S3S118N044P023P042P002(0) <='1';
          else
          cVar1S3S118N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S4S118N044P023P042P002(0) <='1';
          else
          cVar1S4S118N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='0' )then
          cVar1S5S118N044P023P042P002(0) <='1';
          else
          cVar1S5S118N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND A(28)='1' )then
          cVar1S6S118N044P023P042P002(0) <='1';
          else
          cVar1S6S118N044P023P042P002(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S7S118N044P023P042P024(0) <='1';
          else
          cVar1S7S118N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S8S118N044P023P042P024(0) <='1';
          else
          cVar1S8S118N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S9S118N044P023P042P024(0) <='1';
          else
          cVar1S9S118N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='1' )then
          cVar1S10S118N044P023P024P005nsss(0) <='1';
          else
          cVar1S10S118N044P023P024P005nsss(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='0' )then
          cVar1S11S118N044P023P024N005(0) <='1';
          else
          cVar1S11S118N044P023P024N005(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S119P044P025nsss(0) <='1';
          else
          cVar1S0S119P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S119P044N025P023nsss(0) <='1';
          else
          cVar1S1S119P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND A(29)='0' )then
          cVar1S2S119P044N025N023P000(0) <='1';
          else
          cVar1S2S119P044N025N023P000(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND E(20)='1' )then
          cVar1S3S119N044P023P042P053(0) <='1';
          else
          cVar1S3S119N044P023P042P053(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND E(20)='0' )then
          cVar1S4S119N044P023P042N053(0) <='1';
          else
          cVar1S4S119N044P023P042N053(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S5S119N044P023P042P024(0) <='1';
          else
          cVar1S5S119N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S6S119N044P023P042P024(0) <='1';
          else
          cVar1S6S119N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S7S119N044P023P042P024(0) <='1';
          else
          cVar1S7S119N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='1' )then
          cVar1S8S119N044P023P024P008nsss(0) <='1';
          else
          cVar1S8S119N044P023P024P008nsss(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='0' )then
          cVar1S9S119N044P023P024N008(0) <='1';
          else
          cVar1S9S119N044P023P024N008(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='0' )then
          cVar1S10S119N044P023P024N008(0) <='1';
          else
          cVar1S10S119N044P023P024N008(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='1' )then
          cVar1S0S120P044P025nsss(0) <='1';
          else
          cVar1S0S120P044P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='1' )then
          cVar1S1S120P044N025P023nsss(0) <='1';
          else
          cVar1S1S120P044N025P023nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(16)='0' AND B(17)='0' AND A(29)='0' )then
          cVar1S2S120P044N025N023P000(0) <='1';
          else
          cVar1S2S120P044N025N023P000(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND D(11)='0' )then
          cVar1S3S120N044P023P042P054(0) <='1';
          else
          cVar1S3S120N044P023P042P054(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND D(11)='0' )then
          cVar1S4S120N044P023P042P054(0) <='1';
          else
          cVar1S4S120N044P023P042P054(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND D(11)='1' )then
          cVar1S5S120N044P023P042P054(0) <='1';
          else
          cVar1S5S120N044P023P042P054(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S6S120N044P023P042P024(0) <='1';
          else
          cVar1S6S120N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S7S120N044P023P042P024(0) <='1';
          else
          cVar1S7S120N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='1' )then
          cVar1S8S120N044P023P024P005nsss(0) <='1';
          else
          cVar1S8S120N044P023P024P005nsss(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(17)='0' )then
          cVar1S9S120N044P023P024N005(0) <='1';
          else
          cVar1S9S120N044P023P024N005(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='1' )then
          cVar1S0S121P042P023nsss(0) <='1';
          else
          cVar1S0S121P042P023nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='1' )then
          cVar1S1S121P042N023P002nsss(0) <='1';
          else
          cVar1S1S121P042N023P002nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='1' )then
          cVar1S2S121P042N023N002P055nsss(0) <='1';
          else
          cVar1S2S121P042N023N002P055nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='0' )then
          cVar1S3S121P042N023N002N055(0) <='1';
          else
          cVar1S3S121P042N023N002N055(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='0' )then
          cVar1S4S121P042N023N002N055(0) <='1';
          else
          cVar1S4S121P042N023N002N055(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='1' AND E(17)='1' )then
          cVar1S5S121N042P023P052P065(0) <='1';
          else
          cVar1S5S121N042P023P052P065(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='1' AND E(17)='0' )then
          cVar1S6S121N042P023P052N065(0) <='1';
          else
          cVar1S6S121N042P023P052N065(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='1' AND E(17)='0' )then
          cVar1S7S121N042P023P052N065(0) <='1';
          else
          cVar1S7S121N042P023P052N065(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='1' AND E(17)='0' )then
          cVar1S8S121N042P023P052N065(0) <='1';
          else
          cVar1S8S121N042P023P052N065(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='0' AND D(12)='0' )then
          cVar1S9S121N042P023N052P050(0) <='1';
          else
          cVar1S9S121N042P023N052P050(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='0' AND D(12)='0' )then
          cVar1S10S121N042P023N052P050(0) <='1';
          else
          cVar1S10S121N042P023N052P050(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND E(12)='0' AND D(12)='1' )then
          cVar1S11S121N042P023N052P050(0) <='1';
          else
          cVar1S11S121N042P023N052P050(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='1' )then
          cVar1S12S121N042P023P024P008nsss(0) <='1';
          else
          cVar1S12S121N042P023P024P008nsss(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='0' )then
          cVar1S13S121N042P023P024N008(0) <='1';
          else
          cVar1S13S121N042P023P024N008(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='1' AND B(26)='0' AND A(25)='0' )then
          cVar1S14S121N042P023P024N008(0) <='1';
          else
          cVar1S14S121N042P023P024N008(0) <='0';
          end if;
        if(E(14)='1' AND B(25)='0' AND B(16)='1' )then
          cVar1S0S122P044P026P025nsss(0) <='1';
          else
          cVar1S0S122P044P026P025nsss(0) <='0';
          end if;
        if(E(14)='1' AND B(25)='0' AND B(16)='0' AND A(29)='0' )then
          cVar1S1S122P044P026N025P000(0) <='1';
          else
          cVar1S1S122P044P026N025P000(0) <='0';
          end if;
        if(E(14)='1' AND B(25)='0' AND B(16)='0' AND A(29)='0' )then
          cVar1S2S122P044P026N025P000(0) <='1';
          else
          cVar1S2S122P044P026N025P000(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='1' )then
          cVar1S3S122N044P023P042P020(0) <='1';
          else
          cVar1S3S122N044P023P042P020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='1' )then
          cVar1S4S122N044P023P042P020(0) <='1';
          else
          cVar1S4S122N044P023P042P020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='1' )then
          cVar1S5S122N044P023P042P020(0) <='1';
          else
          cVar1S5S122N044P023P042P020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='0' )then
          cVar1S6S122N044P023P042N020(0) <='1';
          else
          cVar1S6S122N044P023P042N020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='0' )then
          cVar1S7S122N044P023P042N020(0) <='1';
          else
          cVar1S7S122N044P023P042N020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='0' AND B(28)='0' )then
          cVar1S8S122N044P023P042N020(0) <='1';
          else
          cVar1S8S122N044P023P042N020(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S9S122N044P023P042P024(0) <='1';
          else
          cVar1S9S122N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='0' AND D(14)='1' AND B(26)='0' )then
          cVar1S10S122N044P023P042P024(0) <='1';
          else
          cVar1S10S122N044P023P042P024(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(26)='1' )then
          cVar1S11S122N044P023P024P006nsss(0) <='1';
          else
          cVar1S11S122N044P023P024P006nsss(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(26)='0' )then
          cVar1S12S122N044P023P024N006(0) <='1';
          else
          cVar1S12S122N044P023P024N006(0) <='0';
          end if;
        if(E(14)='0' AND B(17)='1' AND B(26)='0' AND A(26)='0' )then
          cVar1S13S122N044P023P024N006(0) <='1';
          else
          cVar1S13S122N044P023P024N006(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='1' )then
          cVar1S0S123P042P023nsss(0) <='1';
          else
          cVar1S0S123P042P023nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='1' )then
          cVar1S1S123P042N023P002nsss(0) <='1';
          else
          cVar1S1S123P042N023P002nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='1' )then
          cVar1S2S123P042N023N002P055nsss(0) <='1';
          else
          cVar1S2S123P042N023N002P055nsss(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='0' )then
          cVar1S3S123P042N023N002N055(0) <='1';
          else
          cVar1S3S123P042N023N002N055(0) <='0';
          end if;
        if(D(14)='1' AND B(17)='0' AND A(28)='0' AND D(19)='0' )then
          cVar1S4S123P042N023N002N055(0) <='1';
          else
          cVar1S4S123P042N023N002N055(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='1' AND A(26)='0' )then
          cVar1S5S123N042P023P019P006(0) <='1';
          else
          cVar1S5S123N042P023P019P006(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='1' AND A(26)='0' )then
          cVar1S6S123N042P023P019P006(0) <='1';
          else
          cVar1S6S123N042P023P019P006(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='1' AND A(26)='0' )then
          cVar1S7S123N042P023P019P006(0) <='1';
          else
          cVar1S7S123N042P023P019P006(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='1' AND A(26)='1' )then
          cVar1S8S123N042P023P019P006(0) <='1';
          else
          cVar1S8S123N042P023P019P006(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='0' AND E(16)='1' )then
          cVar1S9S123N042P023N019P069(0) <='1';
          else
          cVar1S9S123N042P023N019P069(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='0' AND E(16)='1' )then
          cVar1S10S123N042P023N019P069(0) <='1';
          else
          cVar1S10S123N042P023N019P069(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='0' AND E(16)='0' )then
          cVar1S11S123N042P023N019N069(0) <='1';
          else
          cVar1S11S123N042P023N019N069(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='0' AND E(16)='0' )then
          cVar1S12S123N042P023N019N069(0) <='1';
          else
          cVar1S12S123N042P023N019N069(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='0' AND A(10)='0' AND E(16)='0' )then
          cVar1S13S123N042P023N019N069(0) <='1';
          else
          cVar1S13S123N042P023N019N069(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='1' AND B(26)='0' AND A(16)='1' )then
          cVar1S14S123N042P023P024P007nsss(0) <='1';
          else
          cVar1S14S123N042P023P024P007nsss(0) <='0';
          end if;
        if(D(14)='0' AND B(17)='1' AND B(26)='0' AND A(16)='0' )then
          cVar1S15S123N042P023P024N007(0) <='1';
          else
          cVar1S15S123N042P023P024N007(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='1' )then
          cVar1S0S124P019P018P067P039(0) <='1';
          else
          cVar1S0S124P019P018P067P039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='1' )then
          cVar1S1S124P019P018P067P039(0) <='1';
          else
          cVar1S1S124P019P018P067P039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='1' )then
          cVar1S2S124P019P018P067P039(0) <='1';
          else
          cVar1S2S124P019P018P067P039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='0' )then
          cVar1S3S124P019P018P067N039(0) <='1';
          else
          cVar1S3S124P019P018P067N039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='0' )then
          cVar1S4S124P019P018P067N039(0) <='1';
          else
          cVar1S4S124P019P018P067N039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='0' AND D(23)='0' )then
          cVar1S5S124P019P018P067N039(0) <='1';
          else
          cVar1S5S124P019P018P067N039(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='1' AND B(24)='0' )then
          cVar1S6S124P019P018P067P028(0) <='1';
          else
          cVar1S6S124P019P018P067P028(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='0' AND D(16)='1' AND B(24)='0' )then
          cVar1S7S124P019P018P067P028(0) <='1';
          else
          cVar1S7S124P019P018P067P028(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='1' AND D(23)='0' AND B(12)='1' )then
          cVar1S8S124P019P018P039P033(0) <='1';
          else
          cVar1S8S124P019P018P039P033(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='1' AND D(23)='0' AND B(12)='1' )then
          cVar1S9S124P019P018P039P033(0) <='1';
          else
          cVar1S9S124P019P018P039P033(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='1' AND D(23)='0' AND B(12)='0' )then
          cVar1S10S124P019P018P039N033(0) <='1';
          else
          cVar1S10S124P019P018P039N033(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='1' AND D(23)='0' AND B(12)='0' )then
          cVar1S11S124P019P018P039N033(0) <='1';
          else
          cVar1S11S124P019P018P039N033(0) <='0';
          end if;
        if(A(10)='0' AND A(20)='1' AND D(23)='1' AND A(11)='0' )then
          cVar1S12S124P019P018P039P017(0) <='1';
          else
          cVar1S12S124P019P018P039P017(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='1' AND D(16)='1' )then
          cVar1S13S124P019P051P042P067nsss(0) <='1';
          else
          cVar1S13S124P019P051P042P067nsss(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='1' AND D(16)='0' )then
          cVar1S14S124P019P051P042N067(0) <='1';
          else
          cVar1S14S124P019P051P042N067(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='1' AND D(16)='0' )then
          cVar1S15S124P019P051P042N067(0) <='1';
          else
          cVar1S15S124P019P051P042N067(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='0' AND B(14)='0' )then
          cVar1S16S124P019P051N042P029(0) <='1';
          else
          cVar1S16S124P019P051N042P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='0' AND B(14)='0' )then
          cVar1S17S124P019P051N042P029(0) <='1';
          else
          cVar1S17S124P019P051N042P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='0' AND B(14)='1' )then
          cVar1S18S124P019P051N042P029(0) <='1';
          else
          cVar1S18S124P019P051N042P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='0' AND D(14)='0' AND B(14)='1' )then
          cVar1S19S124P019P051N042P029(0) <='1';
          else
          cVar1S19S124P019P051N042P029(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='1' AND B(26)='0' )then
          cVar1S20S124P019P051P037P024(0) <='1';
          else
          cVar1S20S124P019P051P037P024(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='1' AND B(26)='0' )then
          cVar1S21S124P019P051P037P024(0) <='1';
          else
          cVar1S21S124P019P051P037P024(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='0' AND A(29)='0' )then
          cVar1S22S124P019P051N037P000(0) <='1';
          else
          cVar1S22S124P019P051N037P000(0) <='0';
          end if;
        if(A(10)='1' AND D(20)='1' AND B(10)='0' AND A(29)='0' )then
          cVar1S23S124P019P051N037P000(0) <='1';
          else
          cVar1S23S124P019P051N037P000(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='0' AND B(22)='0' )then
          cVar1S0S125P018P050P029P032(0) <='1';
          else
          cVar1S0S125P018P050P029P032(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='0' AND B(22)='0' )then
          cVar1S1S125P018P050P029P032(0) <='1';
          else
          cVar1S1S125P018P050P029P032(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='0' AND B(22)='0' )then
          cVar1S2S125P018P050P029P032(0) <='1';
          else
          cVar1S2S125P018P050P029P032(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='0' AND B(22)='1' )then
          cVar1S3S125P018P050P029P032(0) <='1';
          else
          cVar1S3S125P018P050P029P032(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='0' AND B(22)='1' )then
          cVar1S4S125P018P050P029P032(0) <='1';
          else
          cVar1S4S125P018P050P029P032(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='1' AND A(14)='1' )then
          cVar1S5S125P018P050P029P011(0) <='1';
          else
          cVar1S5S125P018P050P029P011(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='0' AND B(14)='1' AND A(14)='0' )then
          cVar1S6S125P018P050P029N011(0) <='1';
          else
          cVar1S6S125P018P050P029N011(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='1' AND A(27)='0' AND A(23)='0' )then
          cVar1S7S125P018P050P004P012(0) <='1';
          else
          cVar1S7S125P018P050P004P012(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='1' AND A(27)='0' AND A(23)='0' )then
          cVar1S8S125P018P050P004P012(0) <='1';
          else
          cVar1S8S125P018P050P004P012(0) <='0';
          end if;
        if(A(20)='1' AND D(12)='1' AND A(27)='0' AND A(23)='1' )then
          cVar1S9S125P018P050P004P012(0) <='1';
          else
          cVar1S9S125P018P050P004P012(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='1' AND D(11)='0' AND B(21)='0' )then
          cVar1S10S125N018P039P054P034(0) <='1';
          else
          cVar1S10S125N018P039P054P034(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='1' AND D(11)='0' AND B(21)='0' )then
          cVar1S11S125N018P039P054P034(0) <='1';
          else
          cVar1S11S125N018P039P054P034(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='1' AND E(10)='1' )then
          cVar1S12S125N018N039P014P060(0) <='1';
          else
          cVar1S12S125N018N039P014P060(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='1' AND E(10)='1' )then
          cVar1S13S125N018N039P014P060(0) <='1';
          else
          cVar1S13S125N018N039P014P060(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='1' AND E(10)='1' )then
          cVar1S14S125N018N039P014P060(0) <='1';
          else
          cVar1S14S125N018N039P014P060(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='1' AND E(10)='0' )then
          cVar1S15S125N018N039P014N060(0) <='1';
          else
          cVar1S15S125N018N039P014N060(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='1' AND E(10)='0' )then
          cVar1S16S125N018N039P014N060(0) <='1';
          else
          cVar1S16S125N018N039P014N060(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='0' AND E(14)='1' )then
          cVar1S17S125N018N039N014P044(0) <='1';
          else
          cVar1S17S125N018N039N014P044(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='0' AND E(14)='0' )then
          cVar1S18S125N018N039N014N044(0) <='1';
          else
          cVar1S18S125N018N039N014N044(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='0' AND E(14)='0' )then
          cVar1S19S125N018N039N014N044(0) <='1';
          else
          cVar1S19S125N018N039N014N044(0) <='0';
          end if;
        if(A(20)='0' AND D(23)='0' AND A(22)='0' AND E(14)='0' )then
          cVar1S20S125N018N039N014N044(0) <='1';
          else
          cVar1S20S125N018N039N014N044(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='1' )then
          cVar1S0S126P018P014P037P004(0) <='1';
          else
          cVar1S0S126P018P014P037P004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='1' )then
          cVar1S1S126P018P014P037P004(0) <='1';
          else
          cVar1S1S126P018P014P037P004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='1' )then
          cVar1S2S126P018P014P037P004(0) <='1';
          else
          cVar1S2S126P018P014P037P004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='0' )then
          cVar1S3S126P018P014P037N004(0) <='1';
          else
          cVar1S3S126P018P014P037N004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='0' )then
          cVar1S4S126P018P014P037N004(0) <='1';
          else
          cVar1S4S126P018P014P037N004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='0' )then
          cVar1S5S126P018P014P037N004(0) <='1';
          else
          cVar1S5S126P018P014P037N004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='0' AND A(27)='0' )then
          cVar1S6S126P018P014P037N004(0) <='1';
          else
          cVar1S6S126P018P014P037N004(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='1' AND A(21)='1' )then
          cVar1S7S126P018P014P037P016(0) <='1';
          else
          cVar1S7S126P018P014P037P016(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='1' AND A(21)='1' )then
          cVar1S8S126P018P014P037P016(0) <='1';
          else
          cVar1S8S126P018P014P037P016(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='1' AND A(21)='0' )then
          cVar1S9S126P018P014P037N016(0) <='1';
          else
          cVar1S9S126P018P014P037N016(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='0' AND B(10)='1' AND A(21)='0' )then
          cVar1S10S126P018P014P037N016(0) <='1';
          else
          cVar1S10S126P018P014P037N016(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='1' AND E(10)='1' AND B(22)='1' )then
          cVar1S11S126P018P014P060P032nsss(0) <='1';
          else
          cVar1S11S126P018P014P060P032nsss(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='1' AND E(10)='1' AND B(22)='0' )then
          cVar1S12S126P018P014P060N032(0) <='1';
          else
          cVar1S12S126P018P014P060N032(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='1' AND E(10)='1' AND B(22)='0' )then
          cVar1S13S126P018P014P060N032(0) <='1';
          else
          cVar1S13S126P018P014P060N032(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='1' AND E(10)='1' AND B(22)='0' )then
          cVar1S14S126P018P014P060N032(0) <='1';
          else
          cVar1S14S126P018P014P060N032(0) <='0';
          end if;
        if(A(20)='0' AND A(22)='1' AND E(10)='0' AND E(14)='0' )then
          cVar1S15S126P018P014N060P044(0) <='1';
          else
          cVar1S15S126P018P014N060P044(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='1' AND B(12)='1' )then
          cVar1S16S126P018P061P033nsss(0) <='1';
          else
          cVar1S16S126P018P061P033nsss(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='1' AND B(12)='0' AND E(13)='0' )then
          cVar1S17S126P018P061N033P048(0) <='1';
          else
          cVar1S17S126P018P061N033P048(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='1' AND B(12)='0' AND E(13)='0' )then
          cVar1S18S126P018P061N033P048(0) <='1';
          else
          cVar1S18S126P018P061N033P048(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='1' AND B(12)='0' AND E(13)='0' )then
          cVar1S19S126P018P061N033P048(0) <='1';
          else
          cVar1S19S126P018P061N033P048(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='1' AND D(17)='1' )then
          cVar1S20S126P018N061P042P063nsss(0) <='1';
          else
          cVar1S20S126P018N061P042P063nsss(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='1' AND D(17)='0' )then
          cVar1S21S126P018N061P042N063(0) <='1';
          else
          cVar1S21S126P018N061P042N063(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='1' AND D(17)='0' )then
          cVar1S22S126P018N061P042N063(0) <='1';
          else
          cVar1S22S126P018N061P042N063(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='0' AND D(12)='0' )then
          cVar1S23S126P018N061N042P050(0) <='1';
          else
          cVar1S23S126P018N061N042P050(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='0' AND D(12)='0' )then
          cVar1S24S126P018N061N042P050(0) <='1';
          else
          cVar1S24S126P018N061N042P050(0) <='0';
          end if;
        if(A(20)='1' AND E(18)='0' AND D(14)='0' AND D(12)='1' )then
          cVar1S25S126P018N061N042P050(0) <='1';
          else
          cVar1S25S126P018N061N042P050(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='1' )then
          cVar1S0S127P017P015P014P010(0) <='1';
          else
          cVar1S0S127P017P015P014P010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='1' )then
          cVar1S1S127P017P015P014P010(0) <='1';
          else
          cVar1S1S127P017P015P014P010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='1' )then
          cVar1S2S127P017P015P014P010(0) <='1';
          else
          cVar1S2S127P017P015P014P010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='0' )then
          cVar1S3S127P017P015P014N010(0) <='1';
          else
          cVar1S3S127P017P015P014N010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='0' )then
          cVar1S4S127P017P015P014N010(0) <='1';
          else
          cVar1S4S127P017P015P014N010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='0' AND A(24)='0' )then
          cVar1S5S127P017P015P014N010(0) <='1';
          else
          cVar1S5S127P017P015P014N010(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='1' AND D( 8)='0' )then
          cVar1S6S127P017P015P014P066(0) <='1';
          else
          cVar1S6S127P017P015P014P066(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='1' AND D( 8)='0' )then
          cVar1S7S127P017P015P014P066(0) <='1';
          else
          cVar1S7S127P017P015P014P066(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='1' AND D( 8)='0' )then
          cVar1S8S127P017P015P014P066(0) <='1';
          else
          cVar1S8S127P017P015P014P066(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='1' AND D( 8)='1' )then
          cVar1S9S127P017P015P014P066(0) <='1';
          else
          cVar1S9S127P017P015P014P066(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='0' AND A(22)='1' AND D( 8)='1' )then
          cVar1S10S127P017P015P014P066(0) <='1';
          else
          cVar1S10S127P017P015P014P066(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='0' AND A(10)='1' )then
          cVar1S11S127P017P015P000P019(0) <='1';
          else
          cVar1S11S127P017P015P000P019(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='0' AND A(10)='1' )then
          cVar1S12S127P017P015P000P019(0) <='1';
          else
          cVar1S12S127P017P015P000P019(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='0' AND A(10)='0' )then
          cVar1S13S127P017P015P000N019(0) <='1';
          else
          cVar1S13S127P017P015P000N019(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='0' AND A(10)='0' )then
          cVar1S14S127P017P015P000N019(0) <='1';
          else
          cVar1S14S127P017P015P000N019(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='1' AND A(25)='0' )then
          cVar1S15S127P017P015P000P008(0) <='1';
          else
          cVar1S15S127P017P015P000P008(0) <='0';
          end if;
        if(A(11)='1' AND A(12)='1' AND A(29)='1' AND A(25)='0' )then
          cVar1S16S127P017P015P000P008(0) <='1';
          else
          cVar1S16S127P017P015P000P008(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='1' AND A(22)='0' )then
          cVar1S17S127N017P018P027P014nsss(0) <='1';
          else
          cVar1S17S127N017P018P027P014nsss(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='0' AND A(28)='1' )then
          cVar1S18S127N017P018N027P002(0) <='1';
          else
          cVar1S18S127N017P018N027P002(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='0' AND A(28)='1' )then
          cVar1S19S127N017P018N027P002(0) <='1';
          else
          cVar1S19S127N017P018N027P002(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='0' AND A(28)='0' )then
          cVar1S20S127N017P018N027N002(0) <='1';
          else
          cVar1S20S127N017P018N027N002(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='0' AND A(28)='0' )then
          cVar1S21S127N017P018N027N002(0) <='1';
          else
          cVar1S21S127N017P018N027N002(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='1' AND B(15)='0' AND A(28)='0' )then
          cVar1S22S127N017P018N027N002(0) <='1';
          else
          cVar1S22S127N017P018N027N002(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='1' AND E(22)='0' )then
          cVar1S23S127N017N018P067P045(0) <='1';
          else
          cVar1S23S127N017N018P067P045(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='1' AND E(22)='0' )then
          cVar1S24S127N017N018P067P045(0) <='1';
          else
          cVar1S24S127N017N018P067P045(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='1' AND E(22)='0' )then
          cVar1S25S127N017N018P067P045(0) <='1';
          else
          cVar1S25S127N017N018P067P045(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='0' )then
          cVar1S26S127N017N018N067P009(0) <='1';
          else
          cVar1S26S127N017N018N067P009(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='0' )then
          cVar1S27S127N017N018N067P009(0) <='1';
          else
          cVar1S27S127N017N018N067P009(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='0' )then
          cVar1S28S127N017N018N067P009(0) <='1';
          else
          cVar1S28S127N017N018N067P009(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='1' )then
          cVar1S29S127N017N018N067P009(0) <='1';
          else
          cVar1S29S127N017N018N067P009(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='1' )then
          cVar1S30S127N017N018N067P009(0) <='1';
          else
          cVar1S30S127N017N018N067P009(0) <='0';
          end if;
        if(A(11)='0' AND A(20)='0' AND D(16)='0' AND A(15)='1' )then
          cVar1S31S127N017N018N067P009(0) <='1';
          else
          cVar1S31S127N017N018N067P009(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV2 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar1S0S0P068P069P012P008(0)='1' AND  A(22)='0' AND D(16)='1' )then
          cVar2S0S0P014P067nsss(0) <='1';
          else
          cVar2S0S0P014P067nsss(0) <='0';
          end if;
        if(cVar1S1S0P068P069P012P008(0)='1' AND  A(22)='1' AND A(13)='0' AND A(12)='0' )then
          cVar2S1S0P014P013P015nsss(0) <='1';
          else
          cVar2S1S0P014P013P015nsss(0) <='0';
          end if;
        if(cVar1S2S0P068N069P065P012(0)='1' AND  D(17)='1' AND A(25)='0' )then
          cVar2S2S0P063P008nsss(0) <='1';
          else
          cVar2S2S0P063P008nsss(0) <='0';
          end if;
        if(cVar1S3S0P068N069N065P055(0)='1' AND  B(23)='1' )then
          cVar2S3S0P030nsss(0) <='1';
          else
          cVar2S3S0P030nsss(0) <='0';
          end if;
        if(cVar1S4S0P068N069N065P055(0)='1' AND  B(23)='0' AND E(19)='1' AND A(20)='1' )then
          cVar2S4S0N030P057P018nsss(0) <='1';
          else
          cVar2S4S0N030P057P018nsss(0) <='0';
          end if;
        if(cVar1S5S0P068N069N065N055(0)='1' AND  E(18)='1' AND B(22)='1' )then
          cVar2S5S0P061P032nsss(0) <='1';
          else
          cVar2S5S0P061P032nsss(0) <='0';
          end if;
        if(cVar1S6S0N068P064P063P065(0)='1' AND  A(23)='0' )then
          cVar2S6S0P012nsss(0) <='1';
          else
          cVar2S6S0P012nsss(0) <='0';
          end if;
        if(cVar1S7S0N068P064N063P035(0)='1' AND  D(16)='1' AND A(22)='0' AND A(11)='1' )then
          cVar2S7S0P067P014P017nsss(0) <='1';
          else
          cVar2S7S0P067P014P017nsss(0) <='0';
          end if;
        if(cVar1S8S0N068P064N063P035(0)='1' AND  D(16)='0' AND E(18)='1' )then
          cVar2S8S0N067P061nsss(0) <='1';
          else
          cVar2S8S0N067P061nsss(0) <='0';
          end if;
        if(cVar1S9S0N068P064N063P035(0)='1' AND  D(16)='0' AND E(18)='0' AND D(20)='1' )then
          cVar2S9S0N067N061P051nsss(0) <='1';
          else
          cVar2S9S0N067N061P051nsss(0) <='0';
          end if;
        if(cVar1S10S0N068P064N063N035(0)='1' AND  B(10)='1' AND D(18)='1' )then
          cVar2S10S0P037P059nsss(0) <='1';
          else
          cVar2S10S0P037P059nsss(0) <='0';
          end if;
        if(cVar1S11S0N068P064N063N035(0)='1' AND  B(10)='0' AND B(21)='1' AND A(21)='1' )then
          cVar2S11S0N037P034P016nsss(0) <='1';
          else
          cVar2S11S0N037P034P016nsss(0) <='0';
          end if;
        if(cVar1S12S0N068N064P067P014(0)='1' AND  E(16)='1' AND E(11)='1' AND B(13)='1' )then
          cVar2S12S0P069P056P031nsss(0) <='1';
          else
          cVar2S12S0P069P056P031nsss(0) <='0';
          end if;
        if(cVar1S13S0N068N064P067P014(0)='1' AND  E(10)='1' AND B(12)='1' )then
          cVar2S13S0P060P033nsss(0) <='1';
          else
          cVar2S13S0P060P033nsss(0) <='0';
          end if;
        if(cVar1S14S0N068N064N067P059(0)='1' AND  B(22)='1' AND E(18)='1' )then
          cVar2S14S0P032P061nsss(0) <='1';
          else
          cVar2S14S0P032P061nsss(0) <='0';
          end if;
        if(cVar1S15S0N068N064N067P059(0)='1' AND  B(22)='0' AND B(12)='1' AND E(10)='1' )then
          cVar2S15S0N032P033P060nsss(0) <='1';
          else
          cVar2S15S0N032P033P060nsss(0) <='0';
          end if;
        if(cVar1S16S0N068N064N067N059(0)='1' AND  E(17)='1' AND D(17)='1' AND E(10)='1' )then
          cVar2S16S0P065P063P060nsss(0) <='1';
          else
          cVar2S16S0P065P063P060nsss(0) <='0';
          end if;
        if(cVar1S17S0N068N064N067N059(0)='1' AND  E(17)='0' AND E(11)='1' AND B(13)='1' )then
          cVar2S17S0N065P056P031nsss(0) <='1';
          else
          cVar2S17S0N065P056P031nsss(0) <='0';
          end if;
        if(cVar1S0S1P067P010P068P069(0)='1' AND  A(22)='0' )then
          cVar2S0S1P014nsss(0) <='1';
          else
          cVar2S0S1P014nsss(0) <='0';
          end if;
        if(cVar1S1S1P067P010P068P069(0)='1' AND  A(22)='1' AND B(26)='0' AND A(23)='0' )then
          cVar2S1S1P014P024P012nsss(0) <='1';
          else
          cVar2S1S1P014P024P012nsss(0) <='0';
          end if;
        if(cVar1S2S1P067P010P068N069(0)='1' AND  A(22)='0' AND A(11)='0' AND B(20)='0' )then
          cVar2S2S1P014P017P036nsss(0) <='1';
          else
          cVar2S2S1P014P017P036nsss(0) <='0';
          end if;
        if(cVar1S3S1P067P010P068N069(0)='1' AND  A(22)='0' AND A(11)='1' AND A(25)='0' )then
          cVar2S3S1P014P017P008nsss(0) <='1';
          else
          cVar2S3S1P014P017P008nsss(0) <='0';
          end if;
        if(cVar1S4S1P067P010P068P012(0)='1' AND  A(15)='0' )then
          cVar2S4S1P009nsss(0) <='1';
          else
          cVar2S4S1P009nsss(0) <='0';
          end if;
        if(cVar1S5S1P067P010P068N012(0)='1' AND  A(25)='1' AND A(21)='0' )then
          cVar2S5S1P008P016nsss(0) <='1';
          else
          cVar2S5S1P008P016nsss(0) <='0';
          end if;
        if(cVar1S6S1P067P010P068N012(0)='1' AND  A(25)='0' AND E(16)='0' )then
          cVar2S6S1N008P069nsss(0) <='1';
          else
          cVar2S6S1N008P069nsss(0) <='0';
          end if;
        if(cVar1S8S1P067P010P024N028(0)='1' AND  A(28)='0' AND A(29)='0' AND A(14)='0' )then
          cVar2S8S1P002P000P011nsss(0) <='1';
          else
          cVar2S8S1P002P000P011nsss(0) <='0';
          end if;
        if(cVar1S9S1N067P068P014P063(0)='1' AND  B(22)='0' )then
          cVar2S9S1P032nsss(0) <='1';
          else
          cVar2S9S1P032nsss(0) <='0';
          end if;
        if(cVar1S10S1N067P068P014P063(0)='1' AND  E(16)='1' )then
          cVar2S10S1P069nsss(0) <='1';
          else
          cVar2S10S1P069nsss(0) <='0';
          end if;
        if(cVar1S11S1N067P068P014P063(0)='1' AND  E(16)='0' AND A(23)='1' )then
          cVar2S11S1N069P012nsss(0) <='1';
          else
          cVar2S11S1N069P012nsss(0) <='0';
          end if;
        if(cVar1S12S1N067P068P014P063(0)='1' AND  E(16)='0' AND A(23)='0' AND E(17)='0' )then
          cVar2S12S1N069N012P065nsss(0) <='1';
          else
          cVar2S12S1N069N012P065nsss(0) <='0';
          end if;
        if(cVar1S13S1N067P068P014P066(0)='1' AND  E(10)='1' )then
          cVar2S13S1P060nsss(0) <='1';
          else
          cVar2S13S1P060nsss(0) <='0';
          end if;
        if(cVar1S14S1N067P068P014P066(0)='1' AND  E(10)='0' AND B(10)='1' )then
          cVar2S14S1N060P037nsss(0) <='1';
          else
          cVar2S14S1N060P037nsss(0) <='0';
          end if;
        if(cVar1S15S1N067P068P014P066(0)='1' AND  E(10)='0' AND B(10)='0' AND A(12)='0' )then
          cVar2S15S1N060N037P015nsss(0) <='1';
          else
          cVar2S15S1N060N037P015nsss(0) <='0';
          end if;
        if(cVar1S16S1N067P068P014N066(0)='1' AND  B(20)='0' AND A(11)='0' AND A(23)='1' )then
          cVar2S16S1P036P017P012nsss(0) <='1';
          else
          cVar2S16S1P036P017P012nsss(0) <='0';
          end if;
        if(cVar1S18S1N067N068P055N030(0)='1' AND  B(24)='1' )then
          cVar2S18S1P028nsss(0) <='1';
          else
          cVar2S18S1P028nsss(0) <='0';
          end if;
        if(cVar1S19S1N067N068P055N030(0)='1' AND  B(24)='0' AND B(13)='1' )then
          cVar2S19S1N028P031nsss(0) <='1';
          else
          cVar2S19S1N028P031nsss(0) <='0';
          end if;
        if(cVar1S20S1N067N068P055N030(0)='1' AND  B(24)='0' AND B(13)='0' AND B(14)='1' )then
          cVar2S20S1N028N031P029nsss(0) <='1';
          else
          cVar2S20S1N028N031P029nsss(0) <='0';
          end if;
        if(cVar1S21S1N067N068N055P052(0)='1' AND  B(14)='1' )then
          cVar2S21S1P029nsss(0) <='1';
          else
          cVar2S21S1P029nsss(0) <='0';
          end if;
        if(cVar1S22S1N067N068N055P052(0)='1' AND  B(14)='0' AND B(15)='1' )then
          cVar2S22S1N029P027nsss(0) <='1';
          else
          cVar2S22S1N029P027nsss(0) <='0';
          end if;
        if(cVar1S23S1N067N068N055P052(0)='1' AND  B(14)='0' AND B(15)='0' AND B(25)='1' )then
          cVar2S23S1N029N027P026nsss(0) <='1';
          else
          cVar2S23S1N029N027P026nsss(0) <='0';
          end if;
        if(cVar1S24S1N067N068N055N052(0)='1' AND  D(14)='1' )then
          cVar2S24S1P042nsss(0) <='1';
          else
          cVar2S24S1P042nsss(0) <='0';
          end if;
        if(cVar1S25S1N067N068N055N052(0)='1' AND  D(14)='0' AND E( 9)='1' )then
          cVar2S25S1N042P064nsss(0) <='1';
          else
          cVar2S25S1N042P064nsss(0) <='0';
          end if;
        if(cVar1S26S1N067N068N055N052(0)='1' AND  D(14)='0' AND E( 9)='0' AND E(17)='1' )then
          cVar2S26S1N042N064P065nsss(0) <='1';
          else
          cVar2S26S1N042N064P065nsss(0) <='0';
          end if;
        if(cVar1S1S2P016P047P000N049(0)='1' AND  B(20)='0' AND E(22)='1' )then
          cVar2S1S2P036P045nsss(0) <='1';
          else
          cVar2S1S2P036P045nsss(0) <='0';
          end if;
        if(cVar1S2S2P016P047P000N049(0)='1' AND  B(20)='0' AND E(22)='0' AND A(12)='0' )then
          cVar2S2S2P036N045P015nsss(0) <='1';
          else
          cVar2S2S2P036N045P015nsss(0) <='0';
          end if;
        if(cVar1S4S2P016N047P052N029(0)='1' AND  E(10)='0' )then
          cVar2S4S2P060nsss(0) <='1';
          else
          cVar2S4S2P060nsss(0) <='0';
          end if;
        if(cVar1S5S2P016N047N052P060(0)='1' AND  E(17)='0' AND B(12)='1' AND D(10)='1' )then
          cVar2S5S2P065P033P058nsss(0) <='1';
          else
          cVar2S5S2P065P033P058nsss(0) <='0';
          end if;
        if(cVar1S6S2P016N047N052P060(0)='1' AND  E(17)='0' AND B(12)='0' )then
          cVar2S6S2P065N033psss(0) <='1';
          else
          cVar2S6S2P065N033psss(0) <='0';
          end if;
        if(cVar1S7S2P016N047N052P060(0)='1' AND  E(17)='1' AND E( 9)='1' )then
          cVar2S7S2P065P064nsss(0) <='1';
          else
          cVar2S7S2P065P064nsss(0) <='0';
          end if;
        if(cVar1S8S2P016N047N052N060(0)='1' AND  D(13)='1' )then
          cVar2S8S2P046nsss(0) <='1';
          else
          cVar2S8S2P046nsss(0) <='0';
          end if;
        if(cVar1S9S2P016N047N052N060(0)='1' AND  D(13)='0' AND E(15)='1' )then
          cVar2S9S2N046P040nsss(0) <='1';
          else
          cVar2S9S2N046P040nsss(0) <='0';
          end if;
        if(cVar1S10S2P016N047N052N060(0)='1' AND  D(13)='0' AND E(15)='0' AND A(12)='0' )then
          cVar2S10S2N046N040P015nsss(0) <='1';
          else
          cVar2S10S2N046N040P015nsss(0) <='0';
          end if;
        if(cVar1S11S2P016P014P063P018(0)='1' AND  B(21)='1' AND A(25)='0' )then
          cVar2S11S2P034P008nsss(0) <='1';
          else
          cVar2S11S2P034P008nsss(0) <='0';
          end if;
        if(cVar1S12S2P016P014P063P018(0)='1' AND  B(21)='0' AND B(20)='1' )then
          cVar2S12S2N034P036nsss(0) <='1';
          else
          cVar2S12S2N034P036nsss(0) <='0';
          end if;
        if(cVar1S13S2P016P014P063P018(0)='1' AND  A(10)='0' AND D(16)='1' )then
          cVar2S13S2P019P067nsss(0) <='1';
          else
          cVar2S13S2P019P067nsss(0) <='0';
          end if;
        if(cVar1S14S2P016P014P063P018(0)='1' AND  A(10)='0' AND D(16)='0' AND D( 9)='1' )then
          cVar2S14S2P019N067P062nsss(0) <='1';
          else
          cVar2S14S2P019N067P062nsss(0) <='0';
          end if;
        if(cVar1S15S2P016P014P063P018(0)='1' AND  A(10)='1' AND A(12)='0' AND D( 8)='1' )then
          cVar2S15S2P019P015P066nsss(0) <='1';
          else
          cVar2S15S2P019P015P066nsss(0) <='0';
          end if;
        if(cVar1S16S2P016P014N063P060(0)='1' AND  A(14)='0' AND D(10)='1' )then
          cVar2S16S2P011P058nsss(0) <='1';
          else
          cVar2S16S2P011P058nsss(0) <='0';
          end if;
        if(cVar1S17S2P016P014N063P060(0)='1' AND  A(14)='0' AND D(10)='0' AND D( 9)='1' )then
          cVar2S17S2P011N058P062nsss(0) <='1';
          else
          cVar2S17S2P011N058P062nsss(0) <='0';
          end if;
        if(cVar1S18S2P016P014N063N060(0)='1' AND  E(17)='0' AND D( 9)='1' AND A(23)='0' )then
          cVar2S18S2P065P062P012nsss(0) <='1';
          else
          cVar2S18S2P065P062P012nsss(0) <='0';
          end if;
        if(cVar1S19S2P016P014N063N060(0)='1' AND  E(17)='0' AND D( 9)='0' AND B(15)='1' )then
          cVar2S19S2P065N062P027nsss(0) <='1';
          else
          cVar2S19S2P065N062P027nsss(0) <='0';
          end if;
        if(cVar1S20S2P016P014P008P010(0)='1' AND  D(16)='1' AND D( 9)='1' )then
          cVar2S20S2P067P062nsss(0) <='1';
          else
          cVar2S20S2P067P062nsss(0) <='0';
          end if;
        if(cVar1S21S2P016P014P008P010(0)='1' AND  D(16)='0' AND E(10)='1' AND A(23)='0' )then
          cVar2S21S2N067P060P012nsss(0) <='1';
          else
          cVar2S21S2N067P060P012nsss(0) <='0';
          end if;
        if(cVar1S22S2P016P014P008P010(0)='1' AND  D(16)='0' AND E(10)='0' AND B(14)='1' )then
          cVar2S22S2N067N060P029nsss(0) <='1';
          else
          cVar2S22S2N067N060P029nsss(0) <='0';
          end if;
        if(cVar1S23S2P016P014P008P010(0)='1' AND  E(14)='0' AND B(24)='1' )then
          cVar2S23S2P044P028nsss(0) <='1';
          else
          cVar2S23S2P044P028nsss(0) <='0';
          end if;
        if(cVar1S24S2P016P014P008P004(0)='1' AND  B(25)='1' )then
          cVar2S24S2P026nsss(0) <='1';
          else
          cVar2S24S2P026nsss(0) <='0';
          end if;
        if(cVar1S1S3P047P049P064P014(0)='1' AND  A(23)='0' )then
          cVar2S1S3P012nsss(0) <='1';
          else
          cVar2S1S3P012nsss(0) <='0';
          end if;
        if(cVar1S6S3N047P052N029N027(0)='1' AND  B(24)='1' )then
          cVar2S6S3P028nsss(0) <='1';
          else
          cVar2S6S3P028nsss(0) <='0';
          end if;
        if(cVar1S7S3N047P052N029N027(0)='1' AND  B(24)='0' AND B(25)='1' AND A(25)='1' )then
          cVar2S7S3N028P026P008nsss(0) <='1';
          else
          cVar2S7S3N028P026P008nsss(0) <='0';
          end if;
        if(cVar1S8S3N047P052N029N027(0)='1' AND  B(24)='0' AND B(25)='0' AND D(12)='0' )then
          cVar2S8S3N028N026P050nsss(0) <='1';
          else
          cVar2S8S3N028N026P050nsss(0) <='0';
          end if;
        if(cVar1S9S3N047N052P060P065(0)='1' AND  B(12)='1' AND A(24)='0' )then
          cVar2S9S3P033P010nsss(0) <='1';
          else
          cVar2S9S3P033P010nsss(0) <='0';
          end if;
        if(cVar1S10S3N047N052P060P065(0)='1' AND  B(12)='0' )then
          cVar2S10S3N033psss(0) <='1';
          else
          cVar2S10S3N033psss(0) <='0';
          end if;
        if(cVar1S11S3N047N052P060P065(0)='1' AND  A(24)='0' AND D(18)='1' )then
          cVar2S11S3P010P059nsss(0) <='1';
          else
          cVar2S11S3P010P059nsss(0) <='0';
          end if;
        if(cVar1S12S3N047N052N060P014(0)='1' AND  D(13)='1' AND B(16)='1' )then
          cVar2S12S3P046P025nsss(0) <='1';
          else
          cVar2S12S3P046P025nsss(0) <='0';
          end if;
        if(cVar1S13S3N047N052N060P014(0)='1' AND  D(13)='1' AND B(16)='0' AND B(15)='1' )then
          cVar2S13S3P046N025P027nsss(0) <='1';
          else
          cVar2S13S3P046N025P027nsss(0) <='0';
          end if;
        if(cVar1S14S3N047N052N060P014(0)='1' AND  D(13)='0' AND B(24)='1' )then
          cVar2S14S3N046P028nsss(0) <='1';
          else
          cVar2S14S3N046P028nsss(0) <='0';
          end if;
        if(cVar1S15S3N047N052N060P014(0)='1' AND  D(13)='0' AND B(24)='0' AND E(15)='1' )then
          cVar2S15S3N046N028P040nsss(0) <='1';
          else
          cVar2S15S3N046N028P040nsss(0) <='0';
          end if;
        if(cVar1S16S3N047N052N060P014(0)='1' AND  B(26)='0' AND D(16)='1' AND A(24)='0' )then
          cVar2S16S3P024P067P010nsss(0) <='1';
          else
          cVar2S16S3P024P067P010nsss(0) <='0';
          end if;
        if(cVar1S17S3N047N052N060P014(0)='1' AND  B(26)='0' AND D(16)='0' AND A(17)='1' )then
          cVar2S17S3P024N067P005nsss(0) <='1';
          else
          cVar2S17S3P024N067P005nsss(0) <='0';
          end if;
        if(cVar1S18S3N047N052N060P014(0)='1' AND  B(26)='1' AND E(22)='1' )then
          cVar2S18S3P024P045nsss(0) <='1';
          else
          cVar2S18S3P024P045nsss(0) <='0';
          end if;
        if(cVar1S0S4P014P069P006P010(0)='1' AND  A(27)='0' )then
          cVar2S0S4P004nsss(0) <='1';
          else
          cVar2S0S4P004nsss(0) <='0';
          end if;
        if(cVar1S1S4P014P069P006P010(0)='1' AND  A(27)='1' AND A(20)='1' )then
          cVar2S1S4P004P018nsss(0) <='1';
          else
          cVar2S1S4P004P018nsss(0) <='0';
          end if;
        if(cVar1S2S4P014P069P006P010(0)='1' AND  D( 9)='0' AND E(12)='1' )then
          cVar2S2S4P062P052nsss(0) <='1';
          else
          cVar2S2S4P062P052nsss(0) <='0';
          end if;
        if(cVar1S3S4P014P069P006P010(0)='1' AND  D( 9)='0' AND E(12)='0' AND A(21)='0' )then
          cVar2S3S4P062N052P016nsss(0) <='1';
          else
          cVar2S3S4P062N052P016nsss(0) <='0';
          end if;
        if(cVar1S4S4P014P069P006P013(0)='1' AND  D( 8)='0' AND A(23)='0' )then
          cVar2S4S4P066P012nsss(0) <='1';
          else
          cVar2S4S4P066P012nsss(0) <='0';
          end if;
        if(cVar1S5S4P014N069P053P051(0)='1' AND  B(24)='1' )then
          cVar2S5S4P028nsss(0) <='1';
          else
          cVar2S5S4P028nsss(0) <='0';
          end if;
        if(cVar1S6S4P014N069P053P051(0)='1' AND  B(24)='0' AND E( 9)='0' )then
          cVar2S6S4N028P064nsss(0) <='1';
          else
          cVar2S6S4N028P064nsss(0) <='0';
          end if;
        if(cVar1S7S4P014N069P053N051(0)='1' AND  D(18)='0' AND E( 8)='1' )then
          cVar2S7S4P059P068nsss(0) <='1';
          else
          cVar2S7S4P059P068nsss(0) <='0';
          end if;
        if(cVar1S8S4P014N069N053P045(0)='1' AND  D(22)='1' )then
          cVar2S8S4P043nsss(0) <='1';
          else
          cVar2S8S4P043nsss(0) <='0';
          end if;
        if(cVar1S9S4P014N069N053P045(0)='1' AND  D(22)='0' AND B(26)='1' )then
          cVar2S9S4N043P024nsss(0) <='1';
          else
          cVar2S9S4N043P024nsss(0) <='0';
          end if;
        if(cVar1S10S4P014N069N053P045(0)='1' AND  D(22)='0' AND B(26)='0' AND E( 8)='0' )then
          cVar2S10S4N043N024P068nsss(0) <='1';
          else
          cVar2S10S4N043N024P068nsss(0) <='0';
          end if;
        if(cVar1S11S4P014N069N053N045(0)='1' AND  B(15)='1' )then
          cVar2S11S4P027nsss(0) <='1';
          else
          cVar2S11S4P027nsss(0) <='0';
          end if;
        if(cVar1S12S4P014N069N053N045(0)='1' AND  B(15)='0' AND E(11)='1' AND A(27)='0' )then
          cVar2S12S4N027P056P004nsss(0) <='1';
          else
          cVar2S12S4N027P056P004nsss(0) <='0';
          end if;
        if(cVar1S13S4P014N069N053N045(0)='1' AND  B(15)='0' AND E(11)='0' )then
          cVar2S13S4N027N056psss(0) <='1';
          else
          cVar2S13S4N027N056psss(0) <='0';
          end if;
        if(cVar1S14S4P014P024P060P010(0)='1' AND  A(20)='0' AND A(15)='0' )then
          cVar2S14S4P018P009nsss(0) <='1';
          else
          cVar2S14S4P018P009nsss(0) <='0';
          end if;
        if(cVar1S15S4P014P024P060P010(0)='1' AND  A(20)='1' AND A(23)='0' )then
          cVar2S15S4P018P012nsss(0) <='1';
          else
          cVar2S15S4P018P012nsss(0) <='0';
          end if;
        if(cVar1S16S4P014P024P060P010(0)='1' AND  A(12)='0' )then
          cVar2S16S4P015nsss(0) <='1';
          else
          cVar2S16S4P015nsss(0) <='0';
          end if;
        if(cVar1S17S4P014P024N060P029(0)='1' AND  E(20)='1' )then
          cVar2S17S4P053nsss(0) <='1';
          else
          cVar2S17S4P053nsss(0) <='0';
          end if;
        if(cVar1S18S4P014P024N060P029(0)='1' AND  E(20)='0' AND B(11)='1' )then
          cVar2S18S4N053P035nsss(0) <='1';
          else
          cVar2S18S4N053P035nsss(0) <='0';
          end if;
        if(cVar1S19S4P014P024N060P029(0)='1' AND  E(20)='0' AND B(11)='0' AND A(11)='0' )then
          cVar2S19S4N053N035P017nsss(0) <='1';
          else
          cVar2S19S4N053N035P017nsss(0) <='0';
          end if;
        if(cVar1S20S4P014P024N060N029(0)='1' AND  A(24)='0' AND B(11)='1' AND A(26)='0' )then
          cVar2S20S4P010P035P006nsss(0) <='1';
          else
          cVar2S20S4P010P035P006nsss(0) <='0';
          end if;
        if(cVar1S21S4P014P024N060N029(0)='1' AND  A(24)='0' AND B(11)='0' AND B(16)='1' )then
          cVar2S21S4P010N035P025nsss(0) <='1';
          else
          cVar2S21S4P010N035P025nsss(0) <='0';
          end if;
        if(cVar1S22S4P014P024N060N029(0)='1' AND  A(24)='1' AND B(20)='0' AND A(18)='1' )then
          cVar2S22S4P010P036P003nsss(0) <='1';
          else
          cVar2S22S4P010P036P003nsss(0) <='0';
          end if;
        if(cVar1S1S5P053P051P024N028(0)='1' AND  B(14)='1' )then
          cVar2S1S5P029nsss(0) <='1';
          else
          cVar2S1S5P029nsss(0) <='0';
          end if;
        if(cVar1S2S5P053P051P024N028(0)='1' AND  B(14)='0' AND B(25)='1' )then
          cVar2S2S5N029P026nsss(0) <='1';
          else
          cVar2S2S5N029P026nsss(0) <='0';
          end if;
        if(cVar1S3S5P053P051P024N028(0)='1' AND  B(14)='0' AND B(25)='0' AND B(15)='1' )then
          cVar2S3S5N029N026P027nsss(0) <='1';
          else
          cVar2S3S5N029N026P027nsss(0) <='0';
          end if;
        if(cVar1S5S5P053N051P010N047(0)='1' AND  E(12)='1' )then
          cVar2S5S5P052nsss(0) <='1';
          else
          cVar2S5S5P052nsss(0) <='0';
          end if;
        if(cVar1S6S5P053N051P010N047(0)='1' AND  E(12)='0' AND A(12)='1' AND A(14)='0' )then
          cVar2S6S5N052P015P011nsss(0) <='1';
          else
          cVar2S6S5N052P015P011nsss(0) <='0';
          end if;
        if(cVar1S7S5P053N051P010N047(0)='1' AND  E(12)='0' AND A(12)='0' AND E( 8)='1' )then
          cVar2S7S5N052N015P068nsss(0) <='1';
          else
          cVar2S7S5N052N015P068nsss(0) <='0';
          end if;
        if(cVar1S9S5N053P051P069P010(0)='1' AND  A(27)='0' AND D(19)='1' AND E(17)='0' )then
          cVar2S9S5P004P055P065nsss(0) <='1';
          else
          cVar2S9S5P004P055P065nsss(0) <='0';
          end if;
        if(cVar1S10S5N053P051P069P010(0)='1' AND  A(27)='0' AND D(19)='0' )then
          cVar2S10S5P004N055psss(0) <='1';
          else
          cVar2S10S5P004N055psss(0) <='0';
          end if;
        if(cVar1S11S5N053P051P069P010(0)='1' AND  A(27)='1' AND D( 8)='0' AND D(16)='1' )then
          cVar2S11S5P004P066P067nsss(0) <='1';
          else
          cVar2S11S5P004P066P067nsss(0) <='0';
          end if;
        if(cVar1S12S5N053P051P069P010(0)='1' AND  E(19)='1' )then
          cVar2S12S5P057nsss(0) <='1';
          else
          cVar2S12S5P057nsss(0) <='0';
          end if;
        if(cVar1S13S5N053P051P069P010(0)='1' AND  E(19)='0' AND E(12)='1' )then
          cVar2S13S5N057P052nsss(0) <='1';
          else
          cVar2S13S5N057P052nsss(0) <='0';
          end if;
        if(cVar1S14S5N053P051N069P045(0)='1' AND  D(22)='1' )then
          cVar2S14S5P043nsss(0) <='1';
          else
          cVar2S14S5P043nsss(0) <='0';
          end if;
        if(cVar1S15S5N053P051N069P045(0)='1' AND  D(22)='0' AND D(21)='1' AND A(21)='0' )then
          cVar2S15S5N043P047P016nsss(0) <='1';
          else
          cVar2S15S5N043P047P016nsss(0) <='0';
          end if;
        if(cVar1S16S5N053P051N069N045(0)='1' AND  E(13)='1' )then
          cVar2S16S5P048nsss(0) <='1';
          else
          cVar2S16S5P048nsss(0) <='0';
          end if;
        if(cVar1S17S5N053P051N069N045(0)='1' AND  E(13)='0' AND E(11)='1' AND D(11)='1' )then
          cVar2S17S5N048P056P054nsss(0) <='1';
          else
          cVar2S17S5N048P056P054nsss(0) <='0';
          end if;
        if(cVar1S18S5N053P051N069N045(0)='1' AND  E(13)='0' AND E(11)='0' AND D(15)='1' )then
          cVar2S18S5N048N056P038nsss(0) <='1';
          else
          cVar2S18S5N048N056P038nsss(0) <='0';
          end if;
        if(cVar1S19S5N053P051P049P061(0)='1' AND  D( 9)='0' AND A(11)='0' )then
          cVar2S19S5P062P017nsss(0) <='1';
          else
          cVar2S19S5P062P017nsss(0) <='0';
          end if;
        if(cVar1S20S5N053P051N049P015(0)='1' AND  E(16)='0' AND E(22)='1' )then
          cVar2S20S5P069P045nsss(0) <='1';
          else
          cVar2S20S5P069P045nsss(0) <='0';
          end if;
        if(cVar1S1S6P047P049P064P012(0)='1' AND  A(21)='0' )then
          cVar2S1S6P016nsss(0) <='1';
          else
          cVar2S1S6P016nsss(0) <='0';
          end if;
        if(cVar1S2S6P047N049P034P035(0)='1' AND  A(15)='1' )then
          cVar2S2S6P009nsss(0) <='1';
          else
          cVar2S2S6P009nsss(0) <='0';
          end if;
        if(cVar1S3S6P047N049P034P035(0)='1' AND  A(15)='0' AND E( 8)='0' )then
          cVar2S3S6N009P068nsss(0) <='1';
          else
          cVar2S3S6N009P068nsss(0) <='0';
          end if;
        if(cVar1S4S6N047P024P055P030(0)='1' AND  E(19)='1' )then
          cVar2S4S6P057nsss(0) <='1';
          else
          cVar2S4S6P057nsss(0) <='0';
          end if;
        if(cVar1S5S6N047P024P055N030(0)='1' AND  B(25)='0' AND B(13)='1' )then
          cVar2S5S6P026P031nsss(0) <='1';
          else
          cVar2S5S6P026P031nsss(0) <='0';
          end if;
        if(cVar1S6S6N047P024P055N030(0)='1' AND  B(25)='0' AND B(13)='0' AND A(27)='0' )then
          cVar2S6S6P026N031P004nsss(0) <='1';
          else
          cVar2S6S6P026N031P004nsss(0) <='0';
          end if;
        if(cVar1S7S6N047P024N055P053(0)='1' AND  D(20)='1' )then
          cVar2S7S6P051nsss(0) <='1';
          else
          cVar2S7S6P051nsss(0) <='0';
          end if;
        if(cVar1S8S6N047P024N055P053(0)='1' AND  D(20)='0' AND A(24)='0' AND E(12)='1' )then
          cVar2S8S6N051P010P052nsss(0) <='1';
          else
          cVar2S8S6N051P010P052nsss(0) <='0';
          end if;
        if(cVar1S9S6N047P024N055N053(0)='1' AND  D(20)='0' )then
          cVar2S9S6P051nsss(0) <='1';
          else
          cVar2S9S6P051nsss(0) <='0';
          end if;
        if(cVar1S10S6N047P024P032P045(0)='1' AND  D(22)='1' )then
          cVar2S10S6P043nsss(0) <='1';
          else
          cVar2S10S6P043nsss(0) <='0';
          end if;
        if(cVar1S11S6N047P024P032N045(0)='1' AND  A(23)='0' AND A(12)='1' AND A(22)='0' )then
          cVar2S11S6P012P015P014nsss(0) <='1';
          else
          cVar2S11S6P012P015P014nsss(0) <='0';
          end if;
        if(cVar1S12S6N047P024P032N045(0)='1' AND  A(23)='0' AND A(12)='0' AND D(13)='1' )then
          cVar2S12S6P012N015P046nsss(0) <='1';
          else
          cVar2S12S6P012N015P046nsss(0) <='0';
          end if;
        if(cVar1S2S7P053P006N028N029(0)='1' AND  B(25)='1' AND A(25)='1' )then
          cVar2S2S7P026P008nsss(0) <='1';
          else
          cVar2S2S7P026P008nsss(0) <='0';
          end if;
        if(cVar1S3S7P053P006N028N029(0)='1' AND  B(25)='1' AND A(25)='0' AND A(10)='0' )then
          cVar2S3S7P026N008P019nsss(0) <='1';
          else
          cVar2S3S7P026N008P019nsss(0) <='0';
          end if;
        if(cVar1S4S7P053P006N028N029(0)='1' AND  B(25)='0' AND B(15)='1' )then
          cVar2S4S7N026P027nsss(0) <='1';
          else
          cVar2S4S7N026P027nsss(0) <='0';
          end if;
        if(cVar1S5S7P053P006P063P017(0)='1' AND  A(10)='1' )then
          cVar2S5S7P019nsss(0) <='1';
          else
          cVar2S5S7P019nsss(0) <='0';
          end if;
        if(cVar1S6S7N053P055P030P057(0)='1' AND  E( 8)='0' )then
          cVar2S6S7P068nsss(0) <='1';
          else
          cVar2S6S7P068nsss(0) <='0';
          end if;
        if(cVar1S7S7N053P055P030P057(0)='1' AND  E( 8)='1' AND A(11)='0' AND B(10)='0' )then
          cVar2S7S7P068P017P037nsss(0) <='1';
          else
          cVar2S7S7P068P017P037nsss(0) <='0';
          end if;
        if(cVar1S8S7N053P055N030P068(0)='1' AND  A(28)='0' AND E(19)='1' )then
          cVar2S8S7P002P057nsss(0) <='1';
          else
          cVar2S8S7P002P057nsss(0) <='0';
          end if;
        if(cVar1S9S7N053P055N030P068(0)='1' AND  A(28)='0' AND E(19)='0' AND A(13)='0' )then
          cVar2S9S7P002N057P013nsss(0) <='1';
          else
          cVar2S9S7P002N057P013nsss(0) <='0';
          end if;
        if(cVar1S10S7N053P055N030P068(0)='1' AND  A(20)='0' AND E(19)='1' )then
          cVar2S10S7P018P057nsss(0) <='1';
          else
          cVar2S10S7P018P057nsss(0) <='0';
          end if;
        if(cVar1S12S7N053N055P047N049(0)='1' AND  B(26)='1' )then
          cVar2S12S7P024nsss(0) <='1';
          else
          cVar2S12S7P024nsss(0) <='0';
          end if;
        if(cVar1S13S7N053N055P047N049(0)='1' AND  B(26)='0' AND A(10)='1' AND A(11)='0' )then
          cVar2S13S7N024P019P017nsss(0) <='1';
          else
          cVar2S13S7N024P019P017nsss(0) <='0';
          end if;
        if(cVar1S14S7N053N055N047P033(0)='1' AND  D(10)='1' AND D(18)='0' )then
          cVar2S14S7P058P059nsss(0) <='1';
          else
          cVar2S14S7P058P059nsss(0) <='0';
          end if;
        if(cVar1S15S7N053N055N047P033(0)='1' AND  D(10)='1' AND D(18)='1' AND A(12)='1' )then
          cVar2S15S7P058P059P015nsss(0) <='1';
          else
          cVar2S15S7P058P059P015nsss(0) <='0';
          end if;
        if(cVar1S16S7N053N055N047P033(0)='1' AND  D(10)='0' AND E(18)='1' AND B(22)='0' )then
          cVar2S16S7N058P061P032nsss(0) <='1';
          else
          cVar2S16S7N058P061P032nsss(0) <='0';
          end if;
        if(cVar1S17S7N053N055N047N033(0)='1' AND  B(17)='1' AND D(14)='1' )then
          cVar2S17S7P023P042nsss(0) <='1';
          else
          cVar2S17S7P023P042nsss(0) <='0';
          end if;
        if(cVar1S18S7N053N055N047N033(0)='1' AND  B(17)='1' AND D(14)='0' AND E(22)='1' )then
          cVar2S18S7P023N042P045nsss(0) <='1';
          else
          cVar2S18S7P023N042P045nsss(0) <='0';
          end if;
        if(cVar1S19S7N053N055N047N033(0)='1' AND  B(17)='0' AND B(27)='1' )then
          cVar2S19S7N023P022nsss(0) <='1';
          else
          cVar2S19S7N023P022nsss(0) <='0';
          end if;
        if(cVar1S1S8P036P053P000N028(0)='1' AND  B(25)='1' )then
          cVar2S1S8P026nsss(0) <='1';
          else
          cVar2S1S8P026nsss(0) <='0';
          end if;
        if(cVar1S2S8P036P053P000N028(0)='1' AND  B(25)='0' AND B(14)='1' )then
          cVar2S2S8N026P029nsss(0) <='1';
          else
          cVar2S2S8N026P029nsss(0) <='0';
          end if;
        if(cVar1S3S8P036P053P000N028(0)='1' AND  B(25)='0' AND B(14)='0' AND E(23)='0' )then
          cVar2S3S8N026N029P041nsss(0) <='1';
          else
          cVar2S3S8N026N029P041nsss(0) <='0';
          end if;
        if(cVar1S5S8P036N053P046N025(0)='1' AND  B(15)='1' )then
          cVar2S5S8P027nsss(0) <='1';
          else
          cVar2S5S8P027nsss(0) <='0';
          end if;
        if(cVar1S6S8P036N053P046N025(0)='1' AND  B(15)='0' AND B(26)='1' )then
          cVar2S6S8N027P024nsss(0) <='1';
          else
          cVar2S6S8N027P024nsss(0) <='0';
          end if;
        if(cVar1S7S8P036N053P046N025(0)='1' AND  B(15)='0' AND B(26)='0' AND A(12)='0' )then
          cVar2S7S8N027N024P015nsss(0) <='1';
          else
          cVar2S7S8N027N024P015nsss(0) <='0';
          end if;
        if(cVar1S8S8P036N053N046P051(0)='1' AND  A(12)='1' )then
          cVar2S8S8P015nsss(0) <='1';
          else
          cVar2S8S8P015nsss(0) <='0';
          end if;
        if(cVar1S9S8P036N053N046P051(0)='1' AND  A(12)='0' AND E(23)='1' AND D(23)='1' )then
          cVar2S9S8N015P041P039nsss(0) <='1';
          else
          cVar2S9S8N015P041P039nsss(0) <='0';
          end if;
        if(cVar1S10S8P036N053N046P051(0)='1' AND  A(12)='0' AND E(23)='0' )then
          cVar2S10S8N015N041psss(0) <='1';
          else
          cVar2S10S8N015N041psss(0) <='0';
          end if;
        if(cVar1S11S8P036N053N046P051(0)='1' AND  E(16)='0' AND A(12)='0' AND A(16)='1' )then
          cVar2S11S8P069P015P007nsss(0) <='1';
          else
          cVar2S11S8P069P015P007nsss(0) <='0';
          end if;
        if(cVar1S12S8P036N053N046P051(0)='1' AND  E(16)='0' AND A(12)='1' AND E(21)='1' )then
          cVar2S12S8P069P015P049nsss(0) <='1';
          else
          cVar2S12S8P069P015P049nsss(0) <='0';
          end if;
        if(cVar1S13S8P036P010P016P008(0)='1' AND  B(26)='0' AND A(20)='0' AND A(29)='0' )then
          cVar2S13S8P024P018P000nsss(0) <='1';
          else
          cVar2S13S8P024P018P000nsss(0) <='0';
          end if;
        if(cVar1S14S8P036P010P016P008(0)='1' AND  B(26)='0' AND A(20)='1' AND A(11)='0' )then
          cVar2S14S8P024P018P017nsss(0) <='1';
          else
          cVar2S14S8P024P018P017nsss(0) <='0';
          end if;
        if(cVar1S15S8P036P010N016P018(0)='1' AND  B(14)='1' )then
          cVar2S15S8P029nsss(0) <='1';
          else
          cVar2S15S8P029nsss(0) <='0';
          end if;
        if(cVar1S16S8P036P010N016P018(0)='1' AND  B(14)='0' AND D( 9)='1' AND E(17)='0' )then
          cVar2S16S8N029P062P065nsss(0) <='1';
          else
          cVar2S16S8N029P062P065nsss(0) <='0';
          end if;
        if(cVar1S17S8P036P010N016P018(0)='1' AND  B(14)='0' AND D( 9)='0' )then
          cVar2S17S8N029N062psss(0) <='1';
          else
          cVar2S17S8N029N062psss(0) <='0';
          end if;
        if(cVar1S18S8P036P010N016N018(0)='1' AND  A(11)='1' AND D( 8)='0' AND B(11)='0' )then
          cVar2S18S8P017P066P035nsss(0) <='1';
          else
          cVar2S18S8P017P066P035nsss(0) <='0';
          end if;
        if(cVar1S19S8P036P010N016N018(0)='1' AND  A(11)='0' AND A(10)='1' AND A(23)='1' )then
          cVar2S19S8N017P019P012nsss(0) <='1';
          else
          cVar2S19S8N017P019P012nsss(0) <='0';
          end if;
        if(cVar1S20S8P036P010P024P004(0)='1' AND  A(20)='1' AND A(22)='0' )then
          cVar2S20S8P018P014nsss(0) <='1';
          else
          cVar2S20S8P018P014nsss(0) <='0';
          end if;
        if(cVar1S3S9P052N029N027N028(0)='1' AND  B(25)='1' AND A(25)='1' )then
          cVar2S3S9P026P008nsss(0) <='1';
          else
          cVar2S3S9P026P008nsss(0) <='0';
          end if;
        if(cVar1S4S9P052N029N027N028(0)='1' AND  B(25)='0' AND D( 9)='1' AND B(11)='0' )then
          cVar2S4S9N026P062P035nsss(0) <='1';
          else
          cVar2S4S9N026P062P035nsss(0) <='0';
          end if;
        if(cVar1S6S9N052P046N025P014(0)='1' AND  B(15)='1' )then
          cVar2S6S9P027nsss(0) <='1';
          else
          cVar2S6S9P027nsss(0) <='0';
          end if;
        if(cVar1S7S9N052P046N025P014(0)='1' AND  B(15)='0' AND B(26)='1' )then
          cVar2S7S9N027P024nsss(0) <='1';
          else
          cVar2S7S9N027P024nsss(0) <='0';
          end if;
        if(cVar1S8S9N052P046N025P014(0)='1' AND  B(15)='0' AND B(26)='0' AND B(12)='1' )then
          cVar2S8S9N027N024P033nsss(0) <='1';
          else
          cVar2S8S9N027N024P033nsss(0) <='0';
          end if;
        if(cVar1S9S9N052N046P041P039(0)='1' AND  B(28)='1' )then
          cVar2S9S9P020nsss(0) <='1';
          else
          cVar2S9S9P020nsss(0) <='0';
          end if;
        if(cVar1S10S9N052N046P041P039(0)='1' AND  B(28)='0' AND B(18)='1' )then
          cVar2S10S9N020P021nsss(0) <='1';
          else
          cVar2S10S9N020P021nsss(0) <='0';
          end if;
        if(cVar1S11S9N052N046P041P039(0)='1' AND  B(28)='0' AND B(18)='0' AND A(23)='0' )then
          cVar2S11S9N020N021P012nsss(0) <='1';
          else
          cVar2S11S9N020N021P012nsss(0) <='0';
          end if;
        if(cVar1S12S9N052N046P041N039(0)='1' AND  E(17)='0' AND D(22)='1' )then
          cVar2S12S9P065P043nsss(0) <='1';
          else
          cVar2S12S9P065P043nsss(0) <='0';
          end if;
        if(cVar1S13S9N052N046N041P039(0)='1' AND  E(20)='1' AND B(24)='1' AND A(23)='0' )then
          cVar2S13S9P053P028P012nsss(0) <='1';
          else
          cVar2S13S9P053P028P012nsss(0) <='0';
          end if;
        if(cVar1S14S9N052N046N041P039(0)='1' AND  E(20)='1' AND B(24)='0' AND B(25)='1' )then
          cVar2S14S9P053N028P026nsss(0) <='1';
          else
          cVar2S14S9P053N028P026nsss(0) <='0';
          end if;
        if(cVar1S15S9N052N046N041P039(0)='1' AND  E(20)='0' AND A(12)='1' AND D(20)='0' )then
          cVar2S15S9N053P015P051nsss(0) <='1';
          else
          cVar2S15S9N053P015P051nsss(0) <='0';
          end if;
        if(cVar1S16S9N052N046N041P039(0)='1' AND  E(20)='0' AND A(12)='0' AND B(17)='1' )then
          cVar2S16S9N053N015P023nsss(0) <='1';
          else
          cVar2S16S9N053N015P023nsss(0) <='0';
          end if;
        if(cVar1S17S9N052N046N041P039(0)='1' AND  A(23)='0' AND E(16)='0' AND A(22)='1' )then
          cVar2S17S9P012P069P014nsss(0) <='1';
          else
          cVar2S17S9P012P069P014nsss(0) <='0';
          end if;
        if(cVar1S1S10P012P053P063N028(0)='1' AND  B(14)='1' )then
          cVar2S1S10P029nsss(0) <='1';
          else
          cVar2S1S10P029nsss(0) <='0';
          end if;
        if(cVar1S2S10P012P053P063N028(0)='1' AND  B(14)='0' AND B(25)='1' )then
          cVar2S2S10N029P026nsss(0) <='1';
          else
          cVar2S2S10N029P026nsss(0) <='0';
          end if;
        if(cVar1S3S10P012P053P063N028(0)='1' AND  B(14)='0' AND B(25)='0' AND E(17)='0' )then
          cVar2S3S10N029N026P065nsss(0) <='1';
          else
          cVar2S3S10N029N026P065nsss(0) <='0';
          end if;
        if(cVar1S4S10P012P053P063P062(0)='1' AND  A(22)='0' AND D(20)='1' )then
          cVar2S4S10P014P051nsss(0) <='1';
          else
          cVar2S4S10P014P051nsss(0) <='0';
          end if;
        if(cVar1S5S10P012N053P041P039(0)='1' AND  B(28)='1' )then
          cVar2S5S10P020nsss(0) <='1';
          else
          cVar2S5S10P020nsss(0) <='0';
          end if;
        if(cVar1S6S10P012N053P041P039(0)='1' AND  B(28)='0' AND B(18)='1' )then
          cVar2S6S10N020P021nsss(0) <='1';
          else
          cVar2S6S10N020P021nsss(0) <='0';
          end if;
        if(cVar1S7S10P012N053P041P039(0)='1' AND  B(28)='0' AND B(18)='0' AND A(20)='0' )then
          cVar2S7S10N020N021P018nsss(0) <='1';
          else
          cVar2S7S10N020N021P018nsss(0) <='0';
          end if;
        if(cVar1S8S10P012N053P041N039(0)='1' AND  E(16)='0' AND A(21)='0' AND D(22)='1' )then
          cVar2S8S10P069P016P043nsss(0) <='1';
          else
          cVar2S8S10P069P016P043nsss(0) <='0';
          end if;
        if(cVar1S9S10P012N053N041P039(0)='1' AND  D(13)='1' )then
          cVar2S9S10P046nsss(0) <='1';
          else
          cVar2S9S10P046nsss(0) <='0';
          end if;
        if(cVar1S10S10P012N053N041P039(0)='1' AND  D(13)='0' AND A(28)='0' AND B(28)='0' )then
          cVar2S10S10N046P002P020nsss(0) <='1';
          else
          cVar2S10S10N046P002P020nsss(0) <='0';
          end if;
        if(cVar1S11S10P012N053N041P039(0)='1' AND  D(13)='0' AND A(28)='1' AND E(15)='1' )then
          cVar2S11S10N046P002P040nsss(0) <='1';
          else
          cVar2S11S10N046P002P040nsss(0) <='0';
          end if;
        if(cVar1S12S10P012N053N041P039(0)='1' AND  D(12)='0' AND A(25)='0' AND B(21)='1' )then
          cVar2S12S10P050P008P034nsss(0) <='1';
          else
          cVar2S12S10P050P008P034nsss(0) <='0';
          end if;
        if(cVar1S13S10P012P030P006P014(0)='1' AND  E(11)='1' )then
          cVar2S13S10P056nsss(0) <='1';
          else
          cVar2S13S10P056nsss(0) <='0';
          end if;
        if(cVar1S14S10P012P030P006P014(0)='1' AND  E(11)='0' AND E(19)='1' )then
          cVar2S14S10N056P057nsss(0) <='1';
          else
          cVar2S14S10N056P057nsss(0) <='0';
          end if;
        if(cVar1S15S10P012P030P006P014(0)='1' AND  E(11)='0' AND E(19)='0' AND A(13)='0' )then
          cVar2S15S10N056N057P013nsss(0) <='1';
          else
          cVar2S15S10N056N057P013nsss(0) <='0';
          end if;
        if(cVar1S16S10P012P030P006P014(0)='1' AND  A(11)='0' AND A(12)='0' )then
          cVar2S16S10P017P015nsss(0) <='1';
          else
          cVar2S16S10P017P015nsss(0) <='0';
          end if;
        if(cVar1S17S10P012N030P008P031(0)='1' AND  D(17)='1' )then
          cVar2S17S10P063nsss(0) <='1';
          else
          cVar2S17S10P063nsss(0) <='0';
          end if;
        if(cVar1S18S10P012N030P008P031(0)='1' AND  D(17)='0' AND D( 8)='1' )then
          cVar2S18S10N063P066nsss(0) <='1';
          else
          cVar2S18S10N063P066nsss(0) <='0';
          end if;
        if(cVar1S19S10P012N030P008P031(0)='1' AND  D(17)='0' AND D( 8)='0' AND A(12)='0' )then
          cVar2S19S10N063N066P015nsss(0) <='1';
          else
          cVar2S19S10N063N066P015nsss(0) <='0';
          end if;
        if(cVar1S20S10P012N030P008N031(0)='1' AND  A(22)='1' AND A(12)='0' AND B(16)='0' )then
          cVar2S20S10P014P015P025nsss(0) <='1';
          else
          cVar2S20S10P014P015P025nsss(0) <='0';
          end if;
        if(cVar1S21S10P012N030P008N031(0)='1' AND  A(22)='1' AND A(12)='1' AND B(22)='1' )then
          cVar2S21S10P014P015P032nsss(0) <='1';
          else
          cVar2S21S10P014P015P032nsss(0) <='0';
          end if;
        if(cVar1S22S10P012N030P008N031(0)='1' AND  A(22)='0' AND D( 8)='1' AND A(10)='1' )then
          cVar2S22S10N014P066P019nsss(0) <='1';
          else
          cVar2S22S10N014P066P019nsss(0) <='0';
          end if;
        if(cVar1S23S10P012N030P008P011(0)='1' AND  E(19)='0' AND B(25)='1' )then
          cVar2S23S10P057P026nsss(0) <='1';
          else
          cVar2S23S10P057P026nsss(0) <='0';
          end if;
        if(cVar1S2S11P053P006N028N029(0)='1' AND  B(25)='1' AND A(25)='1' )then
          cVar2S2S11P026P008nsss(0) <='1';
          else
          cVar2S2S11P026P008nsss(0) <='0';
          end if;
        if(cVar1S3S11P053P006N028N029(0)='1' AND  B(25)='1' AND A(25)='0' AND A(10)='0' )then
          cVar2S3S11P026N008P019nsss(0) <='1';
          else
          cVar2S3S11P026N008P019nsss(0) <='0';
          end if;
        if(cVar1S4S11P053P006N028N029(0)='1' AND  B(25)='0' AND A(15)='1' AND A(24)='0' )then
          cVar2S4S11N026P009P010nsss(0) <='1';
          else
          cVar2S4S11N026P009P010nsss(0) <='0';
          end if;
        if(cVar1S5S11P053P006P063P017(0)='1' AND  A(10)='1' )then
          cVar2S5S11P019nsss(0) <='1';
          else
          cVar2S5S11P019nsss(0) <='0';
          end if;
        if(cVar1S8S11N053P041N020N021(0)='1' AND  A(25)='0' AND E(17)='0' AND E(16)='0' )then
          cVar2S8S11P008P065P069nsss(0) <='1';
          else
          cVar2S8S11P008P065P069nsss(0) <='0';
          end if;
        if(cVar1S9S11N053N041P039P046(0)='1' AND  B(16)='1' )then
          cVar2S9S11P025nsss(0) <='1';
          else
          cVar2S9S11P025nsss(0) <='0';
          end if;
        if(cVar1S10S11N053N041P039P046(0)='1' AND  B(16)='0' AND B(15)='1' )then
          cVar2S10S11N025P027nsss(0) <='1';
          else
          cVar2S10S11N025P027nsss(0) <='0';
          end if;
        if(cVar1S11S11N053N041P039P046(0)='1' AND  B(16)='0' AND B(15)='0' AND B(26)='1' )then
          cVar2S11S11N025N027P024nsss(0) <='1';
          else
          cVar2S11S11N025N027P024nsss(0) <='0';
          end if;
        if(cVar1S12S11N053N041P039N046(0)='1' AND  B(23)='1' AND E(19)='1' )then
          cVar2S12S11P030P057nsss(0) <='1';
          else
          cVar2S12S11P030P057nsss(0) <='0';
          end if;
        if(cVar1S13S11N053N041P039N046(0)='1' AND  B(23)='1' AND E(19)='0' AND D(11)='1' )then
          cVar2S13S11P030N057P054nsss(0) <='1';
          else
          cVar2S13S11P030N057P054nsss(0) <='0';
          end if;
        if(cVar1S14S11N053N041P039N046(0)='1' AND  B(23)='0' AND E(12)='1' AND D(12)='1' )then
          cVar2S14S11N030P052P050nsss(0) <='1';
          else
          cVar2S14S11N030P052P050nsss(0) <='0';
          end if;
        if(cVar1S15S11N053N041P039N046(0)='1' AND  B(23)='0' AND E(12)='0' AND E(22)='1' )then
          cVar2S15S11N030N052P045nsss(0) <='1';
          else
          cVar2S15S11N030N052P045nsss(0) <='0';
          end if;
        if(cVar1S16S11N053N041P039P008(0)='1' AND  A(16)='0' AND A(23)='0' AND A(15)='1' )then
          cVar2S16S11P007P012P009nsss(0) <='1';
          else
          cVar2S16S11P007P012P009nsss(0) <='0';
          end if;
        if(cVar1S0S12P015P016P037P006(0)='1' AND  B(26)='0' AND E( 8)='1' )then
          cVar2S0S12P024P068nsss(0) <='1';
          else
          cVar2S0S12P024P068nsss(0) <='0';
          end if;
        if(cVar1S1S12P015P016P037P006(0)='1' AND  B(26)='0' AND E( 8)='0' AND A(25)='0' )then
          cVar2S1S12P024N068P008nsss(0) <='1';
          else
          cVar2S1S12P024N068P008nsss(0) <='0';
          end if;
        if(cVar1S2S12P015P016P037P006(0)='1' AND  A(20)='1' )then
          cVar2S2S12P018nsss(0) <='1';
          else
          cVar2S2S12P018nsss(0) <='0';
          end if;
        if(cVar1S3S12P015P016N037P063(0)='1' AND  B(21)='1' )then
          cVar2S3S12P034nsss(0) <='1';
          else
          cVar2S3S12P034nsss(0) <='0';
          end if;
        if(cVar1S4S12P015P016N037P063(0)='1' AND  B(21)='0' AND B(20)='1' AND A(22)='0' )then
          cVar2S4S12N034P036P014nsss(0) <='1';
          else
          cVar2S4S12N034P036P014nsss(0) <='0';
          end if;
        if(cVar1S5S12P015P016N037N063(0)='1' AND  E(17)='0' AND B(21)='0' )then
          cVar2S5S12P065P034nsss(0) <='1';
          else
          cVar2S5S12P065P034nsss(0) <='0';
          end if;
        if(cVar1S6S12P015P016N037N063(0)='1' AND  E(17)='1' AND D(16)='1' AND E(16)='0' )then
          cVar2S6S12P065P067P069nsss(0) <='1';
          else
          cVar2S6S12P065P067P069nsss(0) <='0';
          end if;
        if(cVar1S7S12P015N016P065P041(0)='1' AND  B(28)='1' )then
          cVar2S7S12P020nsss(0) <='1';
          else
          cVar2S7S12P020nsss(0) <='0';
          end if;
        if(cVar1S8S12P015N016P065P041(0)='1' AND  B(28)='0' AND A(23)='0' )then
          cVar2S8S12N020P012nsss(0) <='1';
          else
          cVar2S8S12N020P012nsss(0) <='0';
          end if;
        if(cVar1S9S12P015N016P065N041(0)='1' AND  B(15)='1' )then
          cVar2S9S12P027nsss(0) <='1';
          else
          cVar2S9S12P027nsss(0) <='0';
          end if;
        if(cVar1S10S12P015N016P065N041(0)='1' AND  B(15)='0' AND B(21)='0' )then
          cVar2S10S12N027P034nsss(0) <='1';
          else
          cVar2S10S12N027P034nsss(0) <='0';
          end if;
        if(cVar1S11S12P015N016P065N041(0)='1' AND  B(15)='0' AND B(21)='1' AND E(18)='1' )then
          cVar2S11S12N027P034P061nsss(0) <='1';
          else
          cVar2S11S12N027P034P061nsss(0) <='0';
          end if;
        if(cVar1S12S12P015N016P065P004(0)='1' AND  B(21)='1' AND A(22)='1' AND D( 9)='0' )then
          cVar2S12S12P034P014P062nsss(0) <='1';
          else
          cVar2S12S12P034P014P062nsss(0) <='0';
          end if;
        if(cVar1S13S12P015N016P065P004(0)='1' AND  B(21)='1' AND A(22)='0' AND A(11)='1' )then
          cVar2S13S12P034N014P017nsss(0) <='1';
          else
          cVar2S13S12P034N014P017nsss(0) <='0';
          end if;
        if(cVar1S14S12P015N016P065P004(0)='1' AND  B(21)='0' AND A(11)='1' AND A(14)='0' )then
          cVar2S14S12N034P017P011nsss(0) <='1';
          else
          cVar2S14S12N034P017P011nsss(0) <='0';
          end if;
        if(cVar1S15S12P015P016P033P063(0)='1' AND  E(18)='1' )then
          cVar2S15S12P061nsss(0) <='1';
          else
          cVar2S15S12P061nsss(0) <='0';
          end if;
        if(cVar1S16S12P015P016P033P063(0)='1' AND  E(18)='0' AND A(16)='0' )then
          cVar2S16S12N061P007nsss(0) <='1';
          else
          cVar2S16S12N061P007nsss(0) <='0';
          end if;
        if(cVar1S17S12P015P016N033P035(0)='1' AND  D(20)='0' AND A(14)='0' )then
          cVar2S17S12P051P011nsss(0) <='1';
          else
          cVar2S17S12P051P011nsss(0) <='0';
          end if;
        if(cVar1S18S12P015P016N033P035(0)='1' AND  D(20)='0' AND A(14)='1' AND A(13)='0' )then
          cVar2S18S12P051P011P013nsss(0) <='1';
          else
          cVar2S18S12P051P011P013nsss(0) <='0';
          end if;
        if(cVar1S19S12P015P016N033N035(0)='1' AND  E(10)='0' AND E(20)='1' )then
          cVar2S19S12P060P053nsss(0) <='1';
          else
          cVar2S19S12P060P053nsss(0) <='0';
          end if;
        if(cVar1S20S12P015P016N033N035(0)='1' AND  E(10)='0' AND E(20)='0' AND A(22)='1' )then
          cVar2S20S12P060N053P014nsss(0) <='1';
          else
          cVar2S20S12P060N053P014nsss(0) <='0';
          end if;
        if(cVar1S21S12P015P016P006P019(0)='1' AND  D(10)='1' )then
          cVar2S21S12P058nsss(0) <='1';
          else
          cVar2S21S12P058nsss(0) <='0';
          end if;
        if(cVar1S22S12P015P016P006P019(0)='1' AND  D(10)='0' AND E(19)='1' )then
          cVar2S22S12N058P057nsss(0) <='1';
          else
          cVar2S22S12N058P057nsss(0) <='0';
          end if;
        if(cVar1S23S12P015P016P006P019(0)='1' AND  A(11)='0' AND D(10)='0' AND D(11)='0' )then
          cVar2S23S12P017P058P054nsss(0) <='1';
          else
          cVar2S23S12P017P058P054nsss(0) <='0';
          end if;
        if(cVar1S0S13P001P066P011P068(0)='1' AND  E( 9)='1' AND D( 9)='1' )then
          cVar2S0S13P064P062nsss(0) <='1';
          else
          cVar2S0S13P064P062nsss(0) <='0';
          end if;
        if(cVar1S1S13P001P066P011P068(0)='1' AND  E( 9)='1' AND D( 9)='0' AND A(22)='0' )then
          cVar2S1S13P064N062P014nsss(0) <='1';
          else
          cVar2S1S13P064N062P014nsss(0) <='0';
          end if;
        if(cVar1S2S13P001P066P011P068(0)='1' AND  E( 9)='0' AND A(18)='0' AND A(11)='0' )then
          cVar2S2S13N064P003P017nsss(0) <='1';
          else
          cVar2S2S13N064P003P017nsss(0) <='0';
          end if;
        if(cVar1S3S13P001P066P011N068(0)='1' AND  A(25)='0' AND E(10)='1' AND D( 9)='0' )then
          cVar2S3S13P008P060P062nsss(0) <='1';
          else
          cVar2S3S13P008P060P062nsss(0) <='0';
          end if;
        if(cVar1S4S13P001P066P011P002(0)='1' AND  A(20)='1' AND D(16)='1' AND A(25)='0' )then
          cVar2S4S13P018P067P008nsss(0) <='1';
          else
          cVar2S4S13P018P067P008nsss(0) <='0';
          end if;
        if(cVar1S5S13P001P066P011P002(0)='1' AND  A(20)='1' AND D(16)='0' AND E( 8)='1' )then
          cVar2S5S13P018N067P068nsss(0) <='1';
          else
          cVar2S5S13P018N067P068nsss(0) <='0';
          end if;
        if(cVar1S6S13P001P066P011P002(0)='1' AND  A(20)='0' AND A(10)='1' AND D(18)='0' )then
          cVar2S6S13N018P019P059nsss(0) <='1';
          else
          cVar2S6S13N018P019P059nsss(0) <='0';
          end if;
        if(cVar1S7S13P001N066P027P009(0)='1' AND  D(12)='1' )then
          cVar2S7S13P050nsss(0) <='1';
          else
          cVar2S7S13P050nsss(0) <='0';
          end if;
        if(cVar1S8S13P001N066P027P009(0)='1' AND  D(12)='0' AND A(10)='0' )then
          cVar2S8S13N050P019nsss(0) <='1';
          else
          cVar2S8S13N050P019nsss(0) <='0';
          end if;
        if(cVar1S9S13P001N066P027N009(0)='1' AND  E(13)='1' )then
          cVar2S9S13P048nsss(0) <='1';
          else
          cVar2S9S13P048nsss(0) <='0';
          end if;
        if(cVar1S10S13P001N066P027N009(0)='1' AND  E(13)='0' AND D(11)='0' AND D(12)='1' )then
          cVar2S10S13N048P054P050nsss(0) <='1';
          else
          cVar2S10S13N048P054P050nsss(0) <='0';
          end if;
        if(cVar1S11S13P001N066N027P053(0)='1' AND  B(14)='1' )then
          cVar2S11S13P029nsss(0) <='1';
          else
          cVar2S11S13P029nsss(0) <='0';
          end if;
        if(cVar1S12S13P001N066N027P053(0)='1' AND  B(14)='0' AND B(24)='1' )then
          cVar2S12S13N029P028nsss(0) <='1';
          else
          cVar2S12S13N029P028nsss(0) <='0';
          end if;
        if(cVar1S13S13P001N066N027P053(0)='1' AND  B(14)='0' AND B(24)='0' AND B(25)='1' )then
          cVar2S13S13N029N028P026nsss(0) <='1';
          else
          cVar2S13S13N029N028P026nsss(0) <='0';
          end if;
        if(cVar1S14S13P001N066N027N053(0)='1' AND  D(19)='1' AND B(23)='1' )then
          cVar2S14S13P055P030nsss(0) <='1';
          else
          cVar2S14S13P055P030nsss(0) <='0';
          end if;
        if(cVar1S15S13P001N066N027N053(0)='1' AND  D(19)='1' AND B(23)='0' AND B(22)='1' )then
          cVar2S15S13P055N030P032nsss(0) <='1';
          else
          cVar2S15S13P055N030P032nsss(0) <='0';
          end if;
        if(cVar1S16S13P001N066N027N053(0)='1' AND  D(19)='0' AND E(23)='1' AND D(23)='1' )then
          cVar2S16S13N055P041P039nsss(0) <='1';
          else
          cVar2S16S13N055P041P039nsss(0) <='0';
          end if;
        if(cVar1S17S13P001N066N027N053(0)='1' AND  D(19)='0' AND E(23)='0' AND A(12)='1' )then
          cVar2S17S13N055N041P015nsss(0) <='1';
          else
          cVar2S17S13N055N041P015nsss(0) <='0';
          end if;
        if(cVar1S18S13P001P006P051P004(0)='1' AND  A(20)='1' AND A(15)='0' AND A(10)='1' )then
          cVar2S18S13P018P009P019nsss(0) <='1';
          else
          cVar2S18S13P018P009P019nsss(0) <='0';
          end if;
        if(cVar1S19S13P001P006P051P004(0)='1' AND  A(20)='0' AND A(18)='1' AND A(23)='1' )then
          cVar2S19S13N018P003P012nsss(0) <='1';
          else
          cVar2S19S13N018P003P012nsss(0) <='0';
          end if;
        if(cVar1S1S14P015P016P034N063(0)='1' AND  A(14)='0' AND E(17)='0' )then
          cVar2S1S14P011P065nsss(0) <='1';
          else
          cVar2S1S14P011P065nsss(0) <='0';
          end if;
        if(cVar1S2S14P015P016N034P037(0)='1' AND  D(12)='0' AND A(20)='0' )then
          cVar2S2S14P050P018nsss(0) <='1';
          else
          cVar2S2S14P050P018nsss(0) <='0';
          end if;
        if(cVar1S3S14P015P016N034P037(0)='1' AND  D(12)='0' AND A(20)='1' AND B(11)='0' )then
          cVar2S3S14P050P018P035nsss(0) <='1';
          else
          cVar2S3S14P050P018P035nsss(0) <='0';
          end if;
        if(cVar1S4S14P015P016N034N037(0)='1' AND  A(18)='1' AND D( 8)='0' )then
          cVar2S4S14P003P066nsss(0) <='1';
          else
          cVar2S4S14P003P066nsss(0) <='0';
          end if;
        if(cVar1S5S14P015P016N034N037(0)='1' AND  A(18)='0' AND A(15)='1' AND B(26)='0' )then
          cVar2S5S14N003P009P024nsss(0) <='1';
          else
          cVar2S5S14N003P009P024nsss(0) <='0';
          end if;
        if(cVar1S6S14P015P016N034N037(0)='1' AND  A(18)='0' AND A(15)='0' AND D(18)='0' )then
          cVar2S6S14N003N009P059nsss(0) <='1';
          else
          cVar2S6S14N003N009P059nsss(0) <='0';
          end if;
        if(cVar1S8S14P015N016P046N025(0)='1' AND  A(18)='0' AND A(15)='1' )then
          cVar2S8S14P003P009nsss(0) <='1';
          else
          cVar2S8S14P003P009nsss(0) <='0';
          end if;
        if(cVar1S9S14P015N016P046N025(0)='1' AND  A(18)='0' AND A(15)='0' AND B(26)='1' )then
          cVar2S9S14P003N009P024nsss(0) <='1';
          else
          cVar2S9S14P003N009P024nsss(0) <='0';
          end if;
        if(cVar1S10S14P015N016N046P022(0)='1' AND  D(22)='1' )then
          cVar2S10S14P043nsss(0) <='1';
          else
          cVar2S10S14P043nsss(0) <='0';
          end if;
        if(cVar1S11S14P015N016N046P022(0)='1' AND  D(22)='0' AND D(14)='1' )then
          cVar2S11S14N043P042nsss(0) <='1';
          else
          cVar2S11S14N043P042nsss(0) <='0';
          end if;
        if(cVar1S12S14P015N016N046P022(0)='1' AND  D(22)='0' AND D(14)='0' AND A(11)='0' )then
          cVar2S12S14N043N042P017nsss(0) <='1';
          else
          cVar2S12S14N043N042P017nsss(0) <='0';
          end if;
        if(cVar1S13S14P015N016N046N022(0)='1' AND  E(11)='1' AND B(14)='1' )then
          cVar2S13S14P056P029nsss(0) <='1';
          else
          cVar2S13S14P056P029nsss(0) <='0';
          end if;
        if(cVar1S14S14P015N016N046N022(0)='1' AND  E(11)='1' AND B(14)='0' AND A(23)='1' )then
          cVar2S14S14P056N029P012nsss(0) <='1';
          else
          cVar2S14S14P056N029P012nsss(0) <='0';
          end if;
        if(cVar1S15S14P015N016N046N022(0)='1' AND  E(11)='0' AND D(21)='1' AND E(21)='1' )then
          cVar2S15S14N056P047P049nsss(0) <='1';
          else
          cVar2S15S14N056P047P049nsss(0) <='0';
          end if;
        if(cVar1S16S14P015N016N046N022(0)='1' AND  E(11)='0' AND D(21)='0' AND E(17)='0' )then
          cVar2S16S14N056N047P065nsss(0) <='1';
          else
          cVar2S16S14N056N047P065nsss(0) <='0';
          end if;
        if(cVar1S17S14P015P009P016P033(0)='1' AND  E(18)='1' )then
          cVar2S17S14P061nsss(0) <='1';
          else
          cVar2S17S14P061nsss(0) <='0';
          end if;
        if(cVar1S18S14P015P009P016P033(0)='1' AND  E(18)='0' AND B(20)='0' )then
          cVar2S18S14N061P036nsss(0) <='1';
          else
          cVar2S18S14N061P036nsss(0) <='0';
          end if;
        if(cVar1S19S14P015P009P016N033(0)='1' AND  D(12)='0' AND B(11)='1' AND B(21)='0' )then
          cVar2S19S14P050P035P034nsss(0) <='1';
          else
          cVar2S19S14P050P035P034nsss(0) <='0';
          end if;
        if(cVar1S20S14P015P009P016N033(0)='1' AND  D(12)='0' AND B(11)='0' AND E(10)='0' )then
          cVar2S20S14P050N035P060nsss(0) <='1';
          else
          cVar2S20S14P050N035P060nsss(0) <='0';
          end if;
        if(cVar1S21S14P015P009P016P019(0)='1' AND  B(12)='1' AND E(18)='1' )then
          cVar2S21S14P033P061nsss(0) <='1';
          else
          cVar2S21S14P033P061nsss(0) <='0';
          end if;
        if(cVar1S22S14P015P009P016P019(0)='1' AND  B(12)='1' AND E(18)='0' AND E(10)='1' )then
          cVar2S22S14P033N061P060nsss(0) <='1';
          else
          cVar2S22S14P033N061P060nsss(0) <='0';
          end if;
        if(cVar1S23S14P015P009P016P019(0)='1' AND  B(12)='0' AND B(11)='1' AND A(20)='0' )then
          cVar2S23S14N033P035P018nsss(0) <='1';
          else
          cVar2S23S14N033P035P018nsss(0) <='0';
          end if;
        if(cVar1S24S14P015P009P016P019(0)='1' AND  E( 8)='1' AND D( 9)='1' )then
          cVar2S24S14P068P062nsss(0) <='1';
          else
          cVar2S24S14P068P062nsss(0) <='0';
          end if;
        if(cVar1S25S14P015P009P016P019(0)='1' AND  E( 8)='0' AND A(11)='0' AND A(29)='1' )then
          cVar2S25S14N068P017P000nsss(0) <='1';
          else
          cVar2S25S14N068P017P000nsss(0) <='0';
          end if;
        if(cVar1S1S15P046N025P032P014(0)='1' AND  D(21)='1' )then
          cVar2S1S15P047nsss(0) <='1';
          else
          cVar2S1S15P047nsss(0) <='0';
          end if;
        if(cVar1S2S15P046N025P032P014(0)='1' AND  D(21)='0' AND A(21)='0' )then
          cVar2S2S15N047P016nsss(0) <='1';
          else
          cVar2S2S15N047P016nsss(0) <='0';
          end if;
        if(cVar1S3S15P046N025P032P014(0)='1' AND  D(21)='0' AND A(21)='1' AND A(23)='1' )then
          cVar2S3S15N047P016P012nsss(0) <='1';
          else
          cVar2S3S15N047P016P012nsss(0) <='0';
          end if;
        if(cVar1S4S15P046N025P032P014(0)='1' AND  B(11)='0' AND A(13)='0' AND A(12)='0' )then
          cVar2S4S15P035P013P015nsss(0) <='1';
          else
          cVar2S4S15P035P013P015nsss(0) <='0';
          end if;
        if(cVar1S5S15N046P016P018P034(0)='1' AND  A(29)='0' AND D(17)='1' AND A(25)='0' )then
          cVar2S5S15P000P063P008nsss(0) <='1';
          else
          cVar2S5S15P000P063P008nsss(0) <='0';
          end if;
        if(cVar1S6S15N046P016P018P034(0)='1' AND  A(29)='0' AND D(17)='0' AND A(14)='0' )then
          cVar2S6S15P000N063P011nsss(0) <='1';
          else
          cVar2S6S15P000N063P011nsss(0) <='0';
          end if;
        if(cVar1S7S15N046P016P018N034(0)='1' AND  B(11)='1' AND D(20)='0' AND D( 9)='1' )then
          cVar2S7S15P035P051P062nsss(0) <='1';
          else
          cVar2S7S15P035P051P062nsss(0) <='0';
          end if;
        if(cVar1S8S15N046P016P018N034(0)='1' AND  B(11)='0' AND B(20)='1' AND B(26)='0' )then
          cVar2S8S15N035P036P024nsss(0) <='1';
          else
          cVar2S8S15N035P036P024nsss(0) <='0';
          end if;
        if(cVar1S9S15N046P016P018N034(0)='1' AND  B(11)='0' AND B(20)='0' AND E(17)='0' )then
          cVar2S9S15N035N036P065nsss(0) <='1';
          else
          cVar2S9S15N035N036P065nsss(0) <='0';
          end if;
        if(cVar1S10S15N046P016P018P019(0)='1' AND  B(27)='0' AND A(25)='0' AND E(23)='0' )then
          cVar2S10S15P022P008P041nsss(0) <='1';
          else
          cVar2S10S15P022P008P041nsss(0) <='0';
          end if;
        if(cVar1S11S15N046P016P018P019(0)='1' AND  B(27)='0' AND A(25)='1' AND B(10)='1' )then
          cVar2S11S15P022P008P037nsss(0) <='1';
          else
          cVar2S11S15P022P008P037nsss(0) <='0';
          end if;
        if(cVar1S12S15N046P016P018P019(0)='1' AND  E(19)='0' AND E( 8)='1' AND B(21)='1' )then
          cVar2S12S15P057P068P034nsss(0) <='1';
          else
          cVar2S12S15P057P068P034nsss(0) <='0';
          end if;
        if(cVar1S14S15N046N016P056N057(0)='1' AND  B(14)='1' )then
          cVar2S14S15P029nsss(0) <='1';
          else
          cVar2S14S15P029nsss(0) <='0';
          end if;
        if(cVar1S15S15N046N016P056N057(0)='1' AND  B(14)='0' AND A(23)='1' )then
          cVar2S15S15N029P012nsss(0) <='1';
          else
          cVar2S15S15N029P012nsss(0) <='0';
          end if;
        if(cVar1S16S15N046N016N056P054(0)='1' AND  D(21)='1' AND E(21)='1' )then
          cVar2S16S15P047P049nsss(0) <='1';
          else
          cVar2S16S15P047P049nsss(0) <='0';
          end if;
        if(cVar1S17S15N046N016N056P054(0)='1' AND  D(21)='0' AND E(23)='1' AND B(28)='1' )then
          cVar2S17S15N047P041P020nsss(0) <='1';
          else
          cVar2S17S15N047P041P020nsss(0) <='0';
          end if;
        if(cVar1S18S15N046N016N056P054(0)='1' AND  D(21)='0' AND E(23)='0' AND D(15)='1' )then
          cVar2S18S15N047N041P038nsss(0) <='1';
          else
          cVar2S18S15N047N041P038nsss(0) <='0';
          end if;
        if(cVar1S19S15N046N016N056P054(0)='1' AND  B(14)='1' )then
          cVar2S19S15P029nsss(0) <='1';
          else
          cVar2S19S15P029nsss(0) <='0';
          end if;
        if(cVar1S1S16P016P000P023N042(0)='1' AND  E(22)='1' )then
          cVar2S1S16P045nsss(0) <='1';
          else
          cVar2S1S16P045nsss(0) <='0';
          end if;
        if(cVar1S2S16P016P000N023P022(0)='1' AND  D(22)='1' )then
          cVar2S2S16P043nsss(0) <='1';
          else
          cVar2S2S16P043nsss(0) <='0';
          end if;
        if(cVar1S3S16P016P000N023P022(0)='1' AND  D(22)='0' AND A(22)='0' AND D(14)='1' )then
          cVar2S3S16N043P014P042nsss(0) <='1';
          else
          cVar2S3S16N043P014P042nsss(0) <='0';
          end if;
        if(cVar1S4S16P016P000N023N022(0)='1' AND  D(14)='0' )then
          cVar2S4S16P042nsss(0) <='1';
          else
          cVar2S4S16P042nsss(0) <='0';
          end if;
        if(cVar1S5S16P016P000N023N022(0)='1' AND  D(14)='1' AND E(15)='0' AND E(16)='1' )then
          cVar2S5S16P042N040P069nsss(0) <='1';
          else
          cVar2S5S16P042N040P069nsss(0) <='0';
          end if;
        if(cVar1S6S16P016P000P053P062(0)='1' AND  E(10)='0' AND E(11)='0' AND A(28)='0' )then
          cVar2S6S16P060P056P002nsss(0) <='1';
          else
          cVar2S6S16P060P056P002nsss(0) <='0';
          end if;
        if(cVar1S7S16P016P015P034P063(0)='1' AND  A(14)='0' AND A(20)='0' )then
          cVar2S7S16P011P018nsss(0) <='1';
          else
          cVar2S7S16P011P018nsss(0) <='0';
          end if;
        if(cVar1S8S16P016P015P034P063(0)='1' AND  A(14)='0' AND A(20)='1' AND A(11)='1' )then
          cVar2S8S16P011P018P017nsss(0) <='1';
          else
          cVar2S8S16P011P018P017nsss(0) <='0';
          end if;
        if(cVar1S9S16P016P015P034P063(0)='1' AND  A(14)='1' AND A(11)='0' )then
          cVar2S9S16P011P017nsss(0) <='1';
          else
          cVar2S9S16P011P017nsss(0) <='0';
          end if;
        if(cVar1S10S16P016P015P034N063(0)='1' AND  A(29)='0' AND E(17)='0' AND E( 8)='1' )then
          cVar2S10S16P000P065P068nsss(0) <='1';
          else
          cVar2S10S16P000P065P068nsss(0) <='0';
          end if;
        if(cVar1S11S16P016P015N034P037(0)='1' AND  D(12)='0' )then
          cVar2S11S16P050nsss(0) <='1';
          else
          cVar2S11S16P050nsss(0) <='0';
          end if;
        if(cVar1S12S16P016P015N034N037(0)='1' AND  A(18)='1' AND D( 8)='0' AND A(13)='0' )then
          cVar2S12S16P003P066P013nsss(0) <='1';
          else
          cVar2S12S16P003P066P013nsss(0) <='0';
          end if;
        if(cVar1S13S16P016P015N034N037(0)='1' AND  A(18)='0' AND A(15)='1' AND D( 8)='0' )then
          cVar2S13S16N003P009P066nsss(0) <='1';
          else
          cVar2S13S16N003P009P066nsss(0) <='0';
          end if;
        if(cVar1S14S16P016P015N034N037(0)='1' AND  A(18)='0' AND A(15)='0' AND B(20)='1' )then
          cVar2S14S16N003N009P036nsss(0) <='1';
          else
          cVar2S14S16N003N009P036nsss(0) <='0';
          end if;
        if(cVar1S15S16P016P015P006P019(0)='1' AND  E(22)='0' AND B(11)='1' )then
          cVar2S15S16P045P035nsss(0) <='1';
          else
          cVar2S15S16P045P035nsss(0) <='0';
          end if;
        if(cVar1S16S16P016P015P006P019(0)='1' AND  E(22)='0' AND B(11)='0' AND E(18)='1' )then
          cVar2S16S16P045N035P061nsss(0) <='1';
          else
          cVar2S16S16P045N035P061nsss(0) <='0';
          end if;
        if(cVar1S17S16P016P015P006P019(0)='1' AND  B(26)='0' AND E(19)='0' AND E( 8)='1' )then
          cVar2S17S16P024P057P068nsss(0) <='1';
          else
          cVar2S17S16P024P057P068nsss(0) <='0';
          end if;
        if(cVar1S18S16P016P015P006P011(0)='1' AND  B(20)='0' AND A(23)='1' AND A(11)='0' )then
          cVar2S18S16P036P012P017nsss(0) <='1';
          else
          cVar2S18S16P036P012P017nsss(0) <='0';
          end if;
        if(cVar1S2S17P023N042N005P067(0)='1' AND  D( 9)='0' AND B(27)='0' AND D( 8)='0' )then
          cVar2S2S17P062P022P066nsss(0) <='1';
          else
          cVar2S2S17P062P022P066nsss(0) <='0';
          end if;
        if(cVar1S3S17N023P005P053P006(0)='1' AND  B(26)='0' AND B(24)='1' )then
          cVar2S3S17P024P028nsss(0) <='1';
          else
          cVar2S3S17P024P028nsss(0) <='0';
          end if;
        if(cVar1S4S17N023P005P053P006(0)='1' AND  B(26)='0' AND B(24)='0' AND D(23)='0' )then
          cVar2S4S17P024N028P039nsss(0) <='1';
          else
          cVar2S4S17P024N028P039nsss(0) <='0';
          end if;
        if(cVar1S5S17N023P005P053P006(0)='1' AND  D( 9)='0' AND A(11)='0' AND A(23)='1' )then
          cVar2S5S17P062P017P012nsss(0) <='1';
          else
          cVar2S5S17P062P017P012nsss(0) <='0';
          end if;
        if(cVar1S6S17N023P005N053P058(0)='1' AND  A(14)='0' AND B(12)='1' AND A(10)='0' )then
          cVar2S6S17P011P033P019nsss(0) <='1';
          else
          cVar2S6S17P011P033P019nsss(0) <='0';
          end if;
        if(cVar1S7S17N023P005N053P058(0)='1' AND  A(14)='0' AND B(12)='0' AND B(22)='1' )then
          cVar2S7S17P011N033P032nsss(0) <='1';
          else
          cVar2S7S17P011N033P032nsss(0) <='0';
          end if;
        if(cVar1S8S17N023P005N053P058(0)='1' AND  A(14)='1' AND A(13)='0' AND A(12)='1' )then
          cVar2S8S17P011P013P015nsss(0) <='1';
          else
          cVar2S8S17P011P013P015nsss(0) <='0';
          end if;
        if(cVar1S9S17N023P005N053N058(0)='1' AND  B(27)='1' AND A(27)='1' )then
          cVar2S9S17P022P004nsss(0) <='1';
          else
          cVar2S9S17P022P004nsss(0) <='0';
          end if;
        if(cVar1S10S17N023P005N053N058(0)='1' AND  B(27)='1' AND A(27)='0' AND B(11)='0' )then
          cVar2S10S17P022N004P035nsss(0) <='1';
          else
          cVar2S10S17P022N004P035nsss(0) <='0';
          end if;
        if(cVar1S11S17N023P005N053N058(0)='1' AND  B(27)='0' AND D(22)='0' AND B(21)='1' )then
          cVar2S11S17N022P043P034nsss(0) <='1';
          else
          cVar2S11S17N022P043P034nsss(0) <='0';
          end if;
        if(cVar1S12S17N023P005N053N058(0)='1' AND  B(27)='0' AND D(22)='1' AND B(26)='1' )then
          cVar2S12S17N022P043P024nsss(0) <='1';
          else
          cVar2S12S17N022P043P024nsss(0) <='0';
          end if;
        if(cVar1S14S17N023P005P006N041(0)='1' AND  D(21)='1' )then
          cVar2S14S17P047nsss(0) <='1';
          else
          cVar2S14S17P047nsss(0) <='0';
          end if;
        if(cVar1S15S17N023P005P006N041(0)='1' AND  D(21)='0' AND D(22)='1' )then
          cVar2S15S17N047P043nsss(0) <='1';
          else
          cVar2S15S17N047P043nsss(0) <='0';
          end if;
        if(cVar1S0S18P011P058P039P024(0)='1' AND  B(22)='1' )then
          cVar2S0S18P032nsss(0) <='1';
          else
          cVar2S0S18P032nsss(0) <='0';
          end if;
        if(cVar1S1S18P011P058P039P024(0)='1' AND  B(22)='0' AND B(12)='1' )then
          cVar2S1S18N032P033nsss(0) <='1';
          else
          cVar2S1S18N032P033nsss(0) <='0';
          end if;
        if(cVar1S2S18P011P058P039P024(0)='1' AND  B(22)='0' AND B(12)='0' AND B(11)='1' )then
          cVar2S2S18N032N033P035nsss(0) <='1';
          else
          cVar2S2S18N032N033P035nsss(0) <='0';
          end if;
        if(cVar1S3S18P011P058P039P024(0)='1' AND  A(21)='1' )then
          cVar2S3S18P016nsss(0) <='1';
          else
          cVar2S3S18P016nsss(0) <='0';
          end if;
        if(cVar1S5S18P011N058P046N025(0)='1' AND  D(21)='1' )then
          cVar2S5S18P047nsss(0) <='1';
          else
          cVar2S5S18P047nsss(0) <='0';
          end if;
        if(cVar1S6S18P011N058P046N025(0)='1' AND  D(21)='0' AND A(22)='0' )then
          cVar2S6S18N047P014nsss(0) <='1';
          else
          cVar2S6S18N047P014nsss(0) <='0';
          end if;
        if(cVar1S7S18P011N058N046P021(0)='1' AND  E(15)='1' )then
          cVar2S7S18P040nsss(0) <='1';
          else
          cVar2S7S18P040nsss(0) <='0';
          end if;
        if(cVar1S8S18P011N058N046P021(0)='1' AND  E(15)='0' AND D(23)='1' )then
          cVar2S8S18N040P039nsss(0) <='1';
          else
          cVar2S8S18N040P039nsss(0) <='0';
          end if;
        if(cVar1S9S18P011N058N046N021(0)='1' AND  B(28)='1' AND D(23)='1' )then
          cVar2S9S18P020P039nsss(0) <='1';
          else
          cVar2S9S18P020P039nsss(0) <='0';
          end if;
        if(cVar1S10S18P011N058N046N021(0)='1' AND  B(28)='1' AND D(23)='0' AND E(15)='1' )then
          cVar2S10S18P020N039P040nsss(0) <='1';
          else
          cVar2S10S18P020N039P040nsss(0) <='0';
          end if;
        if(cVar1S11S18P011N058N046N021(0)='1' AND  B(28)='0' AND D(23)='0' AND D(15)='0' )then
          cVar2S11S18N020P039P038nsss(0) <='1';
          else
          cVar2S11S18N020P039P038nsss(0) <='0';
          end if;
        if(cVar1S13S18P011P029P066N054(0)='1' AND  D(20)='1' )then
          cVar2S13S18P051nsss(0) <='1';
          else
          cVar2S13S18P051nsss(0) <='0';
          end if;
        if(cVar1S14S18P011P029P066N054(0)='1' AND  D(20)='0' AND E(12)='1' )then
          cVar2S14S18N051P052nsss(0) <='1';
          else
          cVar2S14S18N051P052nsss(0) <='0';
          end if;
        if(cVar1S15S18P011P029P066N054(0)='1' AND  D(20)='0' AND E(12)='0' AND A(22)='0' )then
          cVar2S15S18N051N052P014nsss(0) <='1';
          else
          cVar2S15S18N051N052P014nsss(0) <='0';
          end if;
        if(cVar1S16S18P011N029P013P032(0)='1' AND  A(18)='0' AND B(24)='1' )then
          cVar2S16S18P003P028nsss(0) <='1';
          else
          cVar2S16S18P003P028nsss(0) <='0';
          end if;
        if(cVar1S17S18P011N029P013P032(0)='1' AND  A(18)='0' AND B(24)='0' AND B(15)='1' )then
          cVar2S17S18P003N028P027nsss(0) <='1';
          else
          cVar2S17S18P003N028P027nsss(0) <='0';
          end if;
        if(cVar1S18S18P011N029P013P032(0)='1' AND  A(18)='1' AND A(12)='1' AND A(20)='0' )then
          cVar2S18S18P003P015P018nsss(0) <='1';
          else
          cVar2S18S18P003P015P018nsss(0) <='0';
          end if;
        if(cVar1S19S18P011N029P013P032(0)='1' AND  A(25)='0' AND A(12)='0' AND A(23)='1' )then
          cVar2S19S18P008P015P012nsss(0) <='1';
          else
          cVar2S19S18P008P015P012nsss(0) <='0';
          end if;
        if(cVar1S2S19P021N040N041P056(0)='1' AND  D(16)='0' AND A(26)='1' )then
          cVar2S2S19P067P006nsss(0) <='1';
          else
          cVar2S2S19P067P006nsss(0) <='0';
          end if;
        if(cVar1S3S19P021N040N041P056(0)='1' AND  D(16)='0' AND A(26)='0' AND A(14)='0' )then
          cVar2S3S19P067N006P011nsss(0) <='1';
          else
          cVar2S3S19P067N006P011nsss(0) <='0';
          end if;
        if(cVar1S4S19N021P001P058P039(0)='1' AND  A(14)='0' AND A(13)='1' )then
          cVar2S4S19P011P013nsss(0) <='1';
          else
          cVar2S4S19P011P013nsss(0) <='0';
          end if;
        if(cVar1S5S19N021P001P058P039(0)='1' AND  A(14)='0' AND A(13)='0' AND B(25)='0' )then
          cVar2S5S19P011N013P026nsss(0) <='1';
          else
          cVar2S5S19P011N013P026nsss(0) <='0';
          end if;
        if(cVar1S6S19N021P001N058P020(0)='1' AND  D(23)='1' )then
          cVar2S6S19P039nsss(0) <='1';
          else
          cVar2S6S19P039nsss(0) <='0';
          end if;
        if(cVar1S7S19N021P001N058P020(0)='1' AND  D(23)='0' AND E(15)='1' )then
          cVar2S7S19N039P040nsss(0) <='1';
          else
          cVar2S7S19N039P040nsss(0) <='0';
          end if;
        if(cVar1S8S19N021P001N058P020(0)='1' AND  D(23)='0' AND E(15)='0' AND E( 9)='0' )then
          cVar2S8S19N039N040P064nsss(0) <='1';
          else
          cVar2S8S19N039N040P064nsss(0) <='0';
          end if;
        if(cVar1S9S19N021P001N058N020(0)='1' AND  D(23)='0' AND D(13)='1' )then
          cVar2S9S19P039P046nsss(0) <='1';
          else
          cVar2S9S19P039P046nsss(0) <='0';
          end if;
        if(cVar1S10S19N021P001P051P004(0)='1' AND  E(10)='0' AND A(20)='1' AND B(11)='1' )then
          cVar2S10S19P060P018P035nsss(0) <='1';
          else
          cVar2S10S19P060P018P035nsss(0) <='0';
          end if;
        if(cVar1S2S20P032P023N042N005(0)='1' AND  D(16)='0' AND D(22)='1' )then
          cVar2S2S20P067P043nsss(0) <='1';
          else
          cVar2S2S20P067P043nsss(0) <='0';
          end if;
        if(cVar1S3S20P032N023P005P056(0)='1' AND  A(29)='0' AND D(23)='0' )then
          cVar2S3S20P000P039nsss(0) <='1';
          else
          cVar2S3S20P000P039nsss(0) <='0';
          end if;
        if(cVar1S4S20P032N023P005N056(0)='1' AND  D(11)='0' AND B(11)='1' AND E(22)='0' )then
          cVar2S4S20P054P035P045nsss(0) <='1';
          else
          cVar2S4S20P054P035P045nsss(0) <='0';
          end if;
        if(cVar1S5S20P032N023P005N056(0)='1' AND  D(11)='0' AND B(11)='0' )then
          cVar2S5S20P054N035psss(0) <='1';
          else
          cVar2S5S20P054N035psss(0) <='0';
          end if;
        if(cVar1S6S20P032N023P005N056(0)='1' AND  D(11)='1' AND E(12)='1' AND A(24)='1' )then
          cVar2S6S20P054P052P010nsss(0) <='1';
          else
          cVar2S6S20P054P052P010nsss(0) <='0';
          end if;
        if(cVar1S7S20P032N023P005P031(0)='1' AND  A(26)='0' AND D(23)='1' )then
          cVar2S7S20P006P039nsss(0) <='1';
          else
          cVar2S7S20P006P039nsss(0) <='0';
          end if;
        if(cVar1S8S20P032N023P005P031(0)='1' AND  A(26)='0' AND D(23)='0' AND D(22)='1' )then
          cVar2S8S20P006N039P043nsss(0) <='1';
          else
          cVar2S8S20P006N039P043nsss(0) <='0';
          end if;
        if(cVar1S9S20P032P008P014P051(0)='1' AND  E(10)='1' )then
          cVar2S9S20P060nsss(0) <='1';
          else
          cVar2S9S20P060nsss(0) <='0';
          end if;
        if(cVar1S10S20P032P008P014P051(0)='1' AND  E(10)='0' AND B(21)='0' AND D(17)='0' )then
          cVar2S10S20N060P034P063nsss(0) <='1';
          else
          cVar2S10S20N060P034P063nsss(0) <='0';
          end if;
        if(cVar1S11S20P032P008N014P012(0)='1' AND  E( 9)='1' )then
          cVar2S11S20P064nsss(0) <='1';
          else
          cVar2S11S20P064nsss(0) <='0';
          end if;
        if(cVar1S12S20P032P008N014P012(0)='1' AND  E( 9)='0' AND B(20)='0' AND D( 8)='1' )then
          cVar2S12S20N064P036P066nsss(0) <='1';
          else
          cVar2S12S20N064P036P066nsss(0) <='0';
          end if;
        if(cVar1S13S20P032P008N014N012(0)='1' AND  D(18)='0' AND E(16)='0' AND A(21)='1' )then
          cVar2S13S20P059P069P016nsss(0) <='1';
          else
          cVar2S13S20P059P069P016nsss(0) <='0';
          end if;
        if(cVar1S14S20P032P008N014N012(0)='1' AND  D(18)='1' AND A(12)='1' )then
          cVar2S14S20P059P015nsss(0) <='1';
          else
          cVar2S14S20P059P015nsss(0) <='0';
          end if;
        if(cVar1S15S20P032P008P006P068(0)='1' AND  A(11)='1' )then
          cVar2S15S20P017nsss(0) <='1';
          else
          cVar2S15S20P017nsss(0) <='0';
          end if;
        if(cVar1S2S21P023N042P024N005(0)='1' AND  D(16)='0' AND A(12)='0' AND E( 8)='1' )then
          cVar2S2S21P067P015P068nsss(0) <='1';
          else
          cVar2S2S21P067P015P068nsss(0) <='0';
          end if;
        if(cVar1S3S21N023P001P047P024(0)='1' AND  A(24)='0' )then
          cVar2S3S21P010nsss(0) <='1';
          else
          cVar2S3S21P010nsss(0) <='0';
          end if;
        if(cVar1S4S21N023P001P047N024(0)='1' AND  B(25)='1' )then
          cVar2S4S21P026nsss(0) <='1';
          else
          cVar2S4S21P026nsss(0) <='0';
          end if;
        if(cVar1S5S21N023P001P047N024(0)='1' AND  B(25)='0' AND B(16)='1' )then
          cVar2S5S21N026P025nsss(0) <='1';
          else
          cVar2S5S21N026P025nsss(0) <='0';
          end if;
        if(cVar1S6S21N023P001P047N024(0)='1' AND  B(25)='0' AND B(16)='0' AND B(15)='1' )then
          cVar2S6S21N026N025P027nsss(0) <='1';
          else
          cVar2S6S21N026N025P027nsss(0) <='0';
          end if;
        if(cVar1S7S21N023P001N047P024(0)='1' AND  E(11)='1' AND D(23)='0' AND A(27)='0' )then
          cVar2S7S21P056P039P004nsss(0) <='1';
          else
          cVar2S7S21P056P039P004nsss(0) <='0';
          end if;
        if(cVar1S8S21N023P001N047P024(0)='1' AND  E(11)='0' AND E(12)='1' AND B(14)='1' )then
          cVar2S8S21N056P052P029nsss(0) <='1';
          else
          cVar2S8S21N056P052P029nsss(0) <='0';
          end if;
        if(cVar1S9S21N023P001N047P024(0)='1' AND  B(22)='0' AND D(22)='1' AND A(12)='0' )then
          cVar2S9S21P032P043P015nsss(0) <='1';
          else
          cVar2S9S21P032P043P015nsss(0) <='0';
          end if;
        if(cVar1S10S21N023P001P006P028(0)='1' AND  D(20)='0' AND A(20)='1' AND A(15)='0' )then
          cVar2S10S21P051P018P009nsss(0) <='1';
          else
          cVar2S10S21P051P018P009nsss(0) <='0';
          end if;
        if(cVar1S0S22P001P010P028P027(0)='1' AND  D(12)='1' )then
          cVar2S0S22P050nsss(0) <='1';
          else
          cVar2S0S22P050nsss(0) <='0';
          end if;
        if(cVar1S1S22P001P010P028P027(0)='1' AND  D(12)='0' AND A(15)='1' AND A(22)='0' )then
          cVar2S1S22N050P009P014nsss(0) <='1';
          else
          cVar2S1S22N050P009P014nsss(0) <='0';
          end if;
        if(cVar1S2S22P001P010P028N027(0)='1' AND  D(12)='0' )then
          cVar2S2S22P050nsss(0) <='1';
          else
          cVar2S2S22P050nsss(0) <='0';
          end if;
        if(cVar1S3S22P001P010P028N027(0)='1' AND  D(12)='1' AND B(14)='1' )then
          cVar2S3S22P050P029nsss(0) <='1';
          else
          cVar2S3S22P050P029nsss(0) <='0';
          end if;
        if(cVar1S4S22P001P010P028N027(0)='1' AND  D(12)='1' AND B(14)='0' AND B(25)='1' )then
          cVar2S4S22P050N029P026nsss(0) <='1';
          else
          cVar2S4S22P050N029P026nsss(0) <='0';
          end if;
        if(cVar1S5S22P001P010P028P000(0)='1' AND  A(14)='1' AND D( 8)='0' )then
          cVar2S5S22P011P066nsss(0) <='1';
          else
          cVar2S5S22P011P066nsss(0) <='0';
          end if;
        if(cVar1S6S22P001P010P028P000(0)='1' AND  A(14)='0' AND A(25)='1' )then
          cVar2S6S22N011P008nsss(0) <='1';
          else
          cVar2S6S22N011P008nsss(0) <='0';
          end if;
        if(cVar1S8S22P001P010N028P045(0)='1' AND  B(26)='0' AND B(14)='1' )then
          cVar2S8S22P024P029nsss(0) <='1';
          else
          cVar2S8S22P024P029nsss(0) <='0';
          end if;
        if(cVar1S9S22P001P010N028P045(0)='1' AND  B(26)='0' AND B(14)='0' AND D(10)='1' )then
          cVar2S9S22P024N029P058nsss(0) <='1';
          else
          cVar2S9S22P024N029P058nsss(0) <='0';
          end if;
        if(cVar1S10S22P001P010N028P045(0)='1' AND  B(21)='0' AND A(23)='1' )then
          cVar2S10S22P034P012nsss(0) <='1';
          else
          cVar2S10S22P034P012nsss(0) <='0';
          end if;
        if(cVar1S11S22P001P004P051P024(0)='1' AND  A(21)='1' AND B(11)='1' )then
          cVar2S11S22P016P035nsss(0) <='1';
          else
          cVar2S11S22P016P035nsss(0) <='0';
          end if;
        if(cVar1S12S22P001P004P051P024(0)='1' AND  A(21)='1' AND B(11)='0' AND A(10)='1' )then
          cVar2S12S22P016N035P019nsss(0) <='1';
          else
          cVar2S12S22P016N035P019nsss(0) <='0';
          end if;
        if(cVar1S1S23P027P000N048P035(0)='1' AND  D( 9)='0' AND A(15)='1' )then
          cVar2S1S23P062P009nsss(0) <='1';
          else
          cVar2S1S23P062P009nsss(0) <='0';
          end if;
        if(cVar1S2S23P027P000N048P035(0)='1' AND  D( 9)='0' AND A(15)='0' AND A(22)='0' )then
          cVar2S2S23P062N009P014nsss(0) <='1';
          else
          cVar2S2S23P062N009P014nsss(0) <='0';
          end if;
        if(cVar1S4S23N027P009P023N042(0)='1' AND  E(22)='1' )then
          cVar2S4S23P045nsss(0) <='1';
          else
          cVar2S4S23P045nsss(0) <='0';
          end if;
        if(cVar1S5S23N027P009P023N042(0)='1' AND  E(22)='0' AND E(16)='0' AND B(20)='1' )then
          cVar2S5S23N045P069P036nsss(0) <='1';
          else
          cVar2S5S23N045P069P036nsss(0) <='0';
          end if;
        if(cVar1S6S23N027P009N023P035(0)='1' AND  D( 9)='1' AND D(20)='0' )then
          cVar2S6S23P062P051nsss(0) <='1';
          else
          cVar2S6S23P062P051nsss(0) <='0';
          end if;
        if(cVar1S7S23N027P009N023P035(0)='1' AND  D( 9)='0' AND D(17)='1' AND E(17)='1' )then
          cVar2S7S23N062P063P065nsss(0) <='1';
          else
          cVar2S7S23N062P063P065nsss(0) <='0';
          end if;
        if(cVar1S8S23N027P009N023N035(0)='1' AND  B(27)='1' AND D(22)='1' )then
          cVar2S8S23P022P043nsss(0) <='1';
          else
          cVar2S8S23P022P043nsss(0) <='0';
          end if;
        if(cVar1S9S23N027P009N023N035(0)='1' AND  B(27)='1' AND D(22)='0' AND A(22)='0' )then
          cVar2S9S23P022N043P014nsss(0) <='1';
          else
          cVar2S9S23P022N043P014nsss(0) <='0';
          end if;
        if(cVar1S10S23N027P009N023N035(0)='1' AND  B(27)='0' AND D(22)='0' AND B(18)='1' )then
          cVar2S10S23N022P043P021nsss(0) <='1';
          else
          cVar2S10S23N022P043P021nsss(0) <='0';
          end if;
        if(cVar1S11S23N027P009P068P062(0)='1' AND  D( 8)='0' AND B(20)='1' AND A(10)='1' )then
          cVar2S11S23P066P036P019nsss(0) <='1';
          else
          cVar2S11S23P066P036P019nsss(0) <='0';
          end if;
        if(cVar1S12S23N027P009P068P062(0)='1' AND  D( 8)='0' AND B(20)='0' AND D(21)='1' )then
          cVar2S12S23P066N036P047nsss(0) <='1';
          else
          cVar2S12S23P066N036P047nsss(0) <='0';
          end if;
        if(cVar1S13S23N027P009P068P062(0)='1' AND  A(22)='1' AND E( 9)='1' AND A(10)='0' )then
          cVar2S13S23P014P064P019nsss(0) <='1';
          else
          cVar2S13S23P014P064P019nsss(0) <='0';
          end if;
        if(cVar1S14S23N027P009P068P002(0)='1' AND  D( 8)='1' AND D(18)='1' )then
          cVar2S14S23P066P059nsss(0) <='1';
          else
          cVar2S14S23P066P059nsss(0) <='0';
          end if;
        if(cVar1S0S24P008P026P055P057(0)='1' AND  B(23)='1' )then
          cVar2S0S24P030nsss(0) <='1';
          else
          cVar2S0S24P030nsss(0) <='0';
          end if;
        if(cVar1S1S24P008P026P055P057(0)='1' AND  B(23)='0' AND B(13)='1' )then
          cVar2S1S24N030P031nsss(0) <='1';
          else
          cVar2S1S24N030P031nsss(0) <='0';
          end if;
        if(cVar1S2S24P008P026P055P057(0)='1' AND  B(23)='0' AND B(13)='0' AND E( 8)='0' )then
          cVar2S2S24N030N031P068nsss(0) <='1';
          else
          cVar2S2S24N030N031P068nsss(0) <='0';
          end if;
        if(cVar1S3S24P008P026P055N057(0)='1' AND  A(13)='0' AND A(21)='1' )then
          cVar2S3S24P013P016nsss(0) <='1';
          else
          cVar2S3S24P013P016nsss(0) <='0';
          end if;
        if(cVar1S4S24P008P026P055N057(0)='1' AND  A(13)='0' AND A(21)='0' AND A(22)='1' )then
          cVar2S4S24P013N016P014nsss(0) <='1';
          else
          cVar2S4S24P013N016P014nsss(0) <='0';
          end if;
        if(cVar1S5S24P008P026N055P041(0)='1' AND  B(28)='1' )then
          cVar2S5S24P020nsss(0) <='1';
          else
          cVar2S5S24P020nsss(0) <='0';
          end if;
        if(cVar1S6S24P008P026N055P041(0)='1' AND  B(28)='0' AND B(18)='1' )then
          cVar2S6S24N020P021nsss(0) <='1';
          else
          cVar2S6S24N020P021nsss(0) <='0';
          end if;
        if(cVar1S7S24P008P026N055P041(0)='1' AND  B(28)='0' AND B(18)='0' AND A(27)='1' )then
          cVar2S7S24N020N021P004nsss(0) <='1';
          else
          cVar2S7S24N020N021P004nsss(0) <='0';
          end if;
        if(cVar1S8S24P008P026N055N041(0)='1' AND  D(23)='0' )then
          cVar2S8S24P039nsss(0) <='1';
          else
          cVar2S8S24P039nsss(0) <='0';
          end if;
        if(cVar1S10S24P008P026P045N047(0)='1' AND  D(19)='0' AND A(27)='0' AND A(24)='1' )then
          cVar2S10S24P055P004P010nsss(0) <='1';
          else
          cVar2S10S24P055P004P010nsss(0) <='0';
          end if;
        if(cVar1S12S24P008P026P004N051(0)='1' AND  D(12)='1' )then
          cVar2S12S24P050nsss(0) <='1';
          else
          cVar2S12S24P050nsss(0) <='0';
          end if;
        if(cVar1S13S24P008P026P004N051(0)='1' AND  D(12)='0' AND D( 9)='0' AND D(16)='0' )then
          cVar2S13S24N050P062P067nsss(0) <='1';
          else
          cVar2S13S24N050P062P067nsss(0) <='0';
          end if;
        if(cVar1S14S24P008N026P032P039(0)='1' AND  E( 8)='1' AND E(17)='1' AND D(17)='1' )then
          cVar2S14S24P068P065P063nsss(0) <='1';
          else
          cVar2S14S24P068P065P063nsss(0) <='0';
          end if;
        if(cVar1S15S24P008N026P032P039(0)='1' AND  E( 8)='1' AND E(17)='0' AND D(16)='1' )then
          cVar2S15S24P068N065P067nsss(0) <='1';
          else
          cVar2S15S24P068N065P067nsss(0) <='0';
          end if;
        if(cVar1S16S24P008N026P032P039(0)='1' AND  E( 8)='0' AND B(20)='0' AND B(24)='1' )then
          cVar2S16S24N068P036P028nsss(0) <='1';
          else
          cVar2S16S24N068P036P028nsss(0) <='0';
          end if;
        if(cVar1S17S24P008N026P032P039(0)='1' AND  E( 8)='0' AND B(20)='1' AND B(12)='1' )then
          cVar2S17S24N068P036P033nsss(0) <='1';
          else
          cVar2S17S24N068P036P033nsss(0) <='0';
          end if;
        if(cVar1S0S25P055P026P030P057(0)='1' AND  A(22)='0' )then
          cVar2S0S25P014nsss(0) <='1';
          else
          cVar2S0S25P014nsss(0) <='0';
          end if;
        if(cVar1S1S25P055P026P030P057(0)='1' AND  A(22)='1' AND A(10)='0' )then
          cVar2S1S25P014P019nsss(0) <='1';
          else
          cVar2S1S25P014P019nsss(0) <='0';
          end if;
        if(cVar1S2S25P055P026N030P031(0)='1' AND  A(13)='1' )then
          cVar2S2S25P013nsss(0) <='1';
          else
          cVar2S2S25P013nsss(0) <='0';
          end if;
        if(cVar1S3S25P055P026N030N031(0)='1' AND  A(27)='0' AND A(24)='1' AND E(16)='0' )then
          cVar2S3S25P004P010P069nsss(0) <='1';
          else
          cVar2S3S25P004P010P069nsss(0) <='0';
          end if;
        if(cVar1S4S25P055P026N030N031(0)='1' AND  A(27)='0' AND A(24)='0' AND B(22)='1' )then
          cVar2S4S25P004N010P032nsss(0) <='1';
          else
          cVar2S4S25P004N010P032nsss(0) <='0';
          end if;
        if(cVar1S6S25N055P057P041N020(0)='1' AND  B(18)='1' )then
          cVar2S6S25P021nsss(0) <='1';
          else
          cVar2S6S25P021nsss(0) <='0';
          end if;
        if(cVar1S7S25N055P057P041N020(0)='1' AND  B(18)='0' AND A(25)='0' AND B(11)='0' )then
          cVar2S7S25N021P008P035nsss(0) <='1';
          else
          cVar2S7S25N021P008P035nsss(0) <='0';
          end if;
        if(cVar1S8S25N055P057N041P053(0)='1' AND  B(24)='1' AND A(23)='0' )then
          cVar2S8S25P028P012nsss(0) <='1';
          else
          cVar2S8S25P028P012nsss(0) <='0';
          end if;
        if(cVar1S9S25N055P057N041P053(0)='1' AND  B(24)='0' AND B(14)='1' )then
          cVar2S9S25N028P029nsss(0) <='1';
          else
          cVar2S9S25N028P029nsss(0) <='0';
          end if;
        if(cVar1S10S25N055P057N041P053(0)='1' AND  B(24)='0' AND B(14)='0' AND E(16)='0' )then
          cVar2S10S25N028N029P069nsss(0) <='1';
          else
          cVar2S10S25N028N029P069nsss(0) <='0';
          end if;
        if(cVar1S11S25N055P057N041N053(0)='1' AND  E(15)='1' AND B(18)='1' )then
          cVar2S11S25P040P021nsss(0) <='1';
          else
          cVar2S11S25P040P021nsss(0) <='0';
          end if;
        if(cVar1S12S25N055P057N041N053(0)='1' AND  E(15)='1' AND B(18)='0' AND B(28)='1' )then
          cVar2S12S25P040N021P020nsss(0) <='1';
          else
          cVar2S12S25P040N021P020nsss(0) <='0';
          end if;
        if(cVar1S13S25N055P057P053P037(0)='1' AND  E(18)='0' AND E(16)='0' AND D(18)='1' )then
          cVar2S13S25P061P069P059nsss(0) <='1';
          else
          cVar2S13S25P061P069P059nsss(0) <='0';
          end if;
        if(cVar1S0S26P017P019P037P002(0)='1' AND  D( 9)='1' AND E( 9)='1' )then
          cVar2S0S26P062P064nsss(0) <='1';
          else
          cVar2S0S26P062P064nsss(0) <='0';
          end if;
        if(cVar1S1S26P017P019P037P002(0)='1' AND  D( 9)='1' AND E( 9)='0' AND D( 8)='1' )then
          cVar2S1S26P062N064P066nsss(0) <='1';
          else
          cVar2S1S26P062N064P066nsss(0) <='0';
          end if;
        if(cVar1S2S26P017P019P037P002(0)='1' AND  D( 9)='0' AND D(16)='1' )then
          cVar2S2S26N062P067nsss(0) <='1';
          else
          cVar2S2S26N062P067nsss(0) <='0';
          end if;
        if(cVar1S3S26P017P019P037P002(0)='1' AND  D( 9)='0' AND D(16)='0' AND E( 9)='0' )then
          cVar2S3S26N062N067P064nsss(0) <='1';
          else
          cVar2S3S26N062N067P064nsss(0) <='0';
          end if;
        if(cVar1S4S26P017P019P037P002(0)='1' AND  D( 8)='0' )then
          cVar2S4S26P066nsss(0) <='1';
          else
          cVar2S4S26P066nsss(0) <='0';
          end if;
        if(cVar1S5S26P017P019N037P018(0)='1' AND  D(16)='1' AND A(12)='0' AND A(14)='0' )then
          cVar2S5S26P067P015P011nsss(0) <='1';
          else
          cVar2S5S26P067P015P011nsss(0) <='0';
          end if;
        if(cVar1S6S26P017P019N037P018(0)='1' AND  D(16)='0' AND B(25)='1' )then
          cVar2S6S26N067P026nsss(0) <='1';
          else
          cVar2S6S26N067P026nsss(0) <='0';
          end if;
        if(cVar1S7S26P017P019N037P018(0)='1' AND  D(16)='0' AND B(25)='0' AND B(20)='0' )then
          cVar2S7S26N067N026P036nsss(0) <='1';
          else
          cVar2S7S26N067N026P036nsss(0) <='0';
          end if;
        if(cVar1S8S26P017P019N037P018(0)='1' AND  B(26)='0' AND B(28)='0' AND B(21)='0' )then
          cVar2S8S26P024P020P034nsss(0) <='1';
          else
          cVar2S8S26P024P020P034nsss(0) <='0';
          end if;
        if(cVar1S9S26P017P019N037P018(0)='1' AND  B(26)='1' AND A(25)='1' )then
          cVar2S9S26P024P008nsss(0) <='1';
          else
          cVar2S9S26P024P008nsss(0) <='0';
          end if;
        if(cVar1S11S26P017N019P037P064(0)='1' AND  B(11)='1' AND A(12)='1' )then
          cVar2S11S26P035P015nsss(0) <='1';
          else
          cVar2S11S26P035P015nsss(0) <='0';
          end if;
        if(cVar1S12S26P017N019P037P064(0)='1' AND  B(11)='0' AND D( 8)='1' AND A(13)='0' )then
          cVar2S12S26N035P066P013nsss(0) <='1';
          else
          cVar2S12S26N035P066P013nsss(0) <='0';
          end if;
        if(cVar1S13S26P017N019P037P064(0)='1' AND  B(11)='0' AND D( 8)='0' AND D(10)='1' )then
          cVar2S13S26N035N066P058nsss(0) <='1';
          else
          cVar2S13S26N035N066P058nsss(0) <='0';
          end if;
        if(cVar1S14S26P017N019P037P003(0)='1' AND  A(20)='1' AND A(12)='1' AND D( 8)='0' )then
          cVar2S14S26P018P015P066nsss(0) <='1';
          else
          cVar2S14S26P018P015P066nsss(0) <='0';
          end if;
        if(cVar1S15S26P017N019P037P003(0)='1' AND  A(20)='1' AND A(12)='0' AND A(13)='1' )then
          cVar2S15S26P018N015P013nsss(0) <='1';
          else
          cVar2S15S26P018N015P013nsss(0) <='0';
          end if;
        if(cVar1S16S26P017N019P037P003(0)='1' AND  A(20)='0' AND A(21)='1' AND A(12)='0' )then
          cVar2S16S26N018P016P015nsss(0) <='1';
          else
          cVar2S16S26N018P016P015nsss(0) <='0';
          end if;
        if(cVar1S17S26P017P037P019P064(0)='1' AND  A(20)='1' )then
          cVar2S17S26P018nsss(0) <='1';
          else
          cVar2S17S26P018nsss(0) <='0';
          end if;
        if(cVar1S18S26P017P037P019P064(0)='1' AND  A(20)='0' AND A(12)='0' )then
          cVar2S18S26N018P015nsss(0) <='1';
          else
          cVar2S18S26N018P015nsss(0) <='0';
          end if;
        if(cVar1S19S26P017P037P019N064(0)='1' AND  A(26)='0' AND A(18)='0' )then
          cVar2S19S26P006P003nsss(0) <='1';
          else
          cVar2S19S26P006P003nsss(0) <='0';
          end if;
        if(cVar1S20S26P017P037P019P013(0)='1' AND  A(15)='0' AND D(19)='1' )then
          cVar2S20S26P009P055nsss(0) <='1';
          else
          cVar2S20S26P009P055nsss(0) <='0';
          end if;
        if(cVar1S21S26P017P037P019P013(0)='1' AND  A(15)='0' AND D(19)='0' AND D( 8)='1' )then
          cVar2S21S26P009N055P066nsss(0) <='1';
          else
          cVar2S21S26P009N055P066nsss(0) <='0';
          end if;
        if(cVar1S22S26P017P037P019P013(0)='1' AND  A(15)='1' AND B(20)='1' )then
          cVar2S22S26P009P036nsss(0) <='1';
          else
          cVar2S22S26P009P036nsss(0) <='0';
          end if;
        if(cVar1S23S26P017P037P019P013(0)='1' AND  D( 9)='0' AND B(11)='1' )then
          cVar2S23S26P062P035nsss(0) <='1';
          else
          cVar2S23S26P062P035nsss(0) <='0';
          end if;
        if(cVar1S24S26P017P037P019P013(0)='1' AND  D( 9)='0' AND B(11)='0' AND A(12)='0' )then
          cVar2S24S26P062N035P015nsss(0) <='1';
          else
          cVar2S24S26P062N035P015nsss(0) <='0';
          end if;
        if(cVar1S25S26P017N037P035P019(0)='1' AND  A(12)='0' AND D( 8)='0' )then
          cVar2S25S26P015P066nsss(0) <='1';
          else
          cVar2S25S26P015P066nsss(0) <='0';
          end if;
        if(cVar1S26S26P017N037P035P019(0)='1' AND  A(12)='0' AND D( 8)='1' AND E( 8)='1' )then
          cVar2S26S26P015P066P068nsss(0) <='1';
          else
          cVar2S26S26P015P066P068nsss(0) <='0';
          end if;
        if(cVar1S27S26P017N037P035P019(0)='1' AND  A(12)='1' AND A(21)='0' )then
          cVar2S27S26P015P016nsss(0) <='1';
          else
          cVar2S27S26P015P016nsss(0) <='0';
          end if;
        if(cVar1S28S26P017N037P035P019(0)='1' AND  D(20)='0' AND A(28)='0' AND D(11)='0' )then
          cVar2S28S26P051P002P054nsss(0) <='1';
          else
          cVar2S28S26P051P002P054nsss(0) <='0';
          end if;
        if(cVar1S29S26P017N037N035P064(0)='1' AND  A(18)='1' AND E( 8)='0' AND A(25)='0' )then
          cVar2S29S26P003P068P008nsss(0) <='1';
          else
          cVar2S29S26P003P068P008nsss(0) <='0';
          end if;
        if(cVar1S30S26P017N037N035P064(0)='1' AND  A(14)='1' AND A(20)='1' )then
          cVar2S30S26P011P018nsss(0) <='1';
          else
          cVar2S30S26P011P018nsss(0) <='0';
          end if;
        if(cVar1S31S26P017N037N035P064(0)='1' AND  A(14)='0' AND E(16)='0' AND E( 8)='1' )then
          cVar2S31S26N011P069P068nsss(0) <='1';
          else
          cVar2S31S26N011P069P068nsss(0) <='0';
          end if;
        if(cVar1S0S27P017P051P048P025(0)='1' AND  E(22)='0' AND B(27)='0' )then
          cVar2S0S27P045P022nsss(0) <='1';
          else
          cVar2S0S27P045P022nsss(0) <='0';
          end if;
        if(cVar1S2S27P017P051P058P041(0)='1' AND  A(10)='0' AND A(20)='1' AND A(12)='0' )then
          cVar2S2S27P019P018P015nsss(0) <='1';
          else
          cVar2S2S27P019P018P015nsss(0) <='0';
          end if;
        if(cVar1S3S27P017P051P058P041(0)='1' AND  A(10)='0' AND A(20)='0' AND E(20)='1' )then
          cVar2S3S27P019N018P053nsss(0) <='1';
          else
          cVar2S3S27P019N018P053nsss(0) <='0';
          end if;
        if(cVar1S4S27P017P051P058P041(0)='1' AND  A(10)='1' AND A(22)='0' AND B(10)='1' )then
          cVar2S4S27P019P014P037nsss(0) <='1';
          else
          cVar2S4S27P019P014P037nsss(0) <='0';
          end if;
        if(cVar1S5S27N017P019P067P024(0)='1' AND  A(29)='0' AND A(16)='0' )then
          cVar2S5S27P000P007nsss(0) <='1';
          else
          cVar2S5S27P000P007nsss(0) <='0';
          end if;
        if(cVar1S6S27N017P019P067P024(0)='1' AND  A(29)='0' AND A(16)='1' AND A(23)='1' )then
          cVar2S6S27P000P007P012nsss(0) <='1';
          else
          cVar2S6S27P000P007P012nsss(0) <='0';
          end if;
        if(cVar1S7S27N017P019N067P037(0)='1' AND  D( 9)='1' AND A(12)='0' )then
          cVar2S7S27P062P015nsss(0) <='1';
          else
          cVar2S7S27P062P015nsss(0) <='0';
          end if;
        if(cVar1S8S27N017P019N067P037(0)='1' AND  D( 9)='1' AND A(12)='1' AND D( 8)='1' )then
          cVar2S8S27P062P015P066nsss(0) <='1';
          else
          cVar2S8S27P062P015P066nsss(0) <='0';
          end if;
        if(cVar1S9S27N017P019N067P037(0)='1' AND  D( 9)='0' AND A(16)='1' )then
          cVar2S9S27N062P007nsss(0) <='1';
          else
          cVar2S9S27N062P007nsss(0) <='0';
          end if;
        if(cVar1S10S27N017P019N067P037(0)='1' AND  D( 9)='0' AND A(16)='0' AND E( 9)='0' )then
          cVar2S10S27N062N007P064nsss(0) <='1';
          else
          cVar2S10S27N062N007P064nsss(0) <='0';
          end if;
        if(cVar1S11S27N017P019N067N037(0)='1' AND  A(25)='1' AND B(22)='0' )then
          cVar2S11S27P008P032nsss(0) <='1';
          else
          cVar2S11S27P008P032nsss(0) <='0';
          end if;
        if(cVar1S12S27N017N019P068P027(0)='1' AND  E(13)='1' )then
          cVar2S12S27P048nsss(0) <='1';
          else
          cVar2S12S27P048nsss(0) <='0';
          end if;
        if(cVar1S13S27N017N019P068P027(0)='1' AND  E(13)='0' AND A(15)='1' )then
          cVar2S13S27N048P009nsss(0) <='1';
          else
          cVar2S13S27N048P009nsss(0) <='0';
          end if;
        if(cVar1S14S27N017N019P068P027(0)='1' AND  E(13)='0' AND A(15)='0' AND B(25)='0' )then
          cVar2S14S27N048N009P026nsss(0) <='1';
          else
          cVar2S14S27N048N009P026nsss(0) <='0';
          end if;
        if(cVar1S15S27N017N019P068N027(0)='1' AND  B(14)='1' AND A(14)='1' )then
          cVar2S15S27P029P011nsss(0) <='1';
          else
          cVar2S15S27P029P011nsss(0) <='0';
          end if;
        if(cVar1S16S27N017N019P068N027(0)='1' AND  B(14)='1' AND A(14)='0' AND A(15)='1' )then
          cVar2S16S27P029N011P009nsss(0) <='1';
          else
          cVar2S16S27P029N011P009nsss(0) <='0';
          end if;
        if(cVar1S17S27N017N019P068N027(0)='1' AND  B(14)='0' AND B(17)='1' )then
          cVar2S17S27N029P023nsss(0) <='1';
          else
          cVar2S17S27N029P023nsss(0) <='0';
          end if;
        if(cVar1S18S27N017N019P068N027(0)='1' AND  B(14)='0' AND B(17)='0' AND B(16)='1' )then
          cVar2S18S27N029N023P025nsss(0) <='1';
          else
          cVar2S18S27N029N023P025nsss(0) <='0';
          end if;
        if(cVar1S19S27N017N019P068P018(0)='1' AND  D(19)='0' AND E(17)='0' AND A(18)='0' )then
          cVar2S19S27P055P065P003nsss(0) <='1';
          else
          cVar2S19S27P055P065P003nsss(0) <='0';
          end if;
        if(cVar1S20S27N017N019P068N018(0)='1' AND  D(16)='0' AND B(28)='0' AND E(19)='1' )then
          cVar2S20S27P067P020P057nsss(0) <='1';
          else
          cVar2S20S27P067P020P057nsss(0) <='0';
          end if;
        if(cVar1S0S28P017P068P064P044(0)='1' AND  B(17)='1' )then
          cVar2S0S28P023nsss(0) <='1';
          else
          cVar2S0S28P023nsss(0) <='0';
          end if;
        if(cVar1S1S28P017P068P064P044(0)='1' AND  B(17)='0' AND B(27)='1' )then
          cVar2S1S28N023P022nsss(0) <='1';
          else
          cVar2S1S28N023P022nsss(0) <='0';
          end if;
        if(cVar1S2S28P017P068P064P044(0)='1' AND  B(17)='0' AND B(27)='0' AND A(16)='1' )then
          cVar2S2S28N023N022P007nsss(0) <='1';
          else
          cVar2S2S28N023N022P007nsss(0) <='0';
          end if;
        if(cVar1S3S28P017P068P064N044(0)='1' AND  D(14)='0' )then
          cVar2S3S28P042nsss(0) <='1';
          else
          cVar2S3S28P042nsss(0) <='0';
          end if;
        if(cVar1S4S28P017P068P064N044(0)='1' AND  D(14)='1' AND E(15)='1' )then
          cVar2S4S28P042P040nsss(0) <='1';
          else
          cVar2S4S28P042P040nsss(0) <='0';
          end if;
        if(cVar1S6S28P017P068P064N055(0)='1' AND  D(16)='1' AND E(17)='0' AND A(22)='0' )then
          cVar2S6S28P067P065P014nsss(0) <='1';
          else
          cVar2S6S28P067P065P014nsss(0) <='0';
          end if;
        if(cVar1S7S28P017P068P064N055(0)='1' AND  D(16)='0' AND D( 9)='1' AND D(10)='1' )then
          cVar2S7S28N067P062P058nsss(0) <='1';
          else
          cVar2S7S28N067P062P058nsss(0) <='0';
          end if;
        if(cVar1S8S28P017P068P019P064(0)='1' AND  A(15)='0' AND B(21)='1' )then
          cVar2S8S28P009P034nsss(0) <='1';
          else
          cVar2S8S28P009P034nsss(0) <='0';
          end if;
        if(cVar1S9S28P017P068P019P064(0)='1' AND  A(15)='0' AND B(21)='0' AND A(13)='0' )then
          cVar2S9S28P009N034P013nsss(0) <='1';
          else
          cVar2S9S28P009N034P013nsss(0) <='0';
          end if;
        if(cVar1S10S28P017P068P019N064(0)='1' AND  B(11)='0' AND A(28)='0' )then
          cVar2S10S28P035P002nsss(0) <='1';
          else
          cVar2S10S28P035P002nsss(0) <='0';
          end if;
        if(cVar1S11S28P017P068N019P067(0)='1' AND  D(17)='0' AND B(10)='0' AND A(23)='0' )then
          cVar2S11S28P063P037P012nsss(0) <='1';
          else
          cVar2S11S28P063P037P012nsss(0) <='0';
          end if;
        if(cVar1S12S28P017P068N019P067(0)='1' AND  D(17)='0' AND B(10)='1' AND A(21)='1' )then
          cVar2S12S28P063P037P016nsss(0) <='1';
          else
          cVar2S12S28P063P037P016nsss(0) <='0';
          end if;
        if(cVar1S13S28P017P068N019P067(0)='1' AND  D(17)='1' AND A(12)='1' )then
          cVar2S13S28P063P015nsss(0) <='1';
          else
          cVar2S13S28P063P015nsss(0) <='0';
          end if;
        if(cVar1S14S28P017P019P016P067(0)='1' AND  E(14)='0' AND A(23)='1' AND A(27)='0' )then
          cVar2S14S28P044P012P004nsss(0) <='1';
          else
          cVar2S14S28P044P012P004nsss(0) <='0';
          end if;
        if(cVar1S15S28P017P019P016P067(0)='1' AND  E(14)='0' AND A(23)='0' AND E(17)='0' )then
          cVar2S15S28P044N012P065nsss(0) <='1';
          else
          cVar2S15S28P044N012P065nsss(0) <='0';
          end if;
        if(cVar1S16S28P017P019P016P067(0)='1' AND  E(17)='1' )then
          cVar2S16S28P065nsss(0) <='1';
          else
          cVar2S16S28P065nsss(0) <='0';
          end if;
        if(cVar1S17S28P017P019P016P067(0)='1' AND  E(17)='0' AND B(10)='1' AND A(20)='1' )then
          cVar2S17S28N065P037P018nsss(0) <='1';
          else
          cVar2S17S28N065P037P018nsss(0) <='0';
          end if;
        if(cVar1S18S28P017P019N016P010(0)='1' AND  A(29)='0' AND A(15)='0' )then
          cVar2S18S28P000P009nsss(0) <='1';
          else
          cVar2S18S28P000P009nsss(0) <='0';
          end if;
        if(cVar1S19S28P017P019N016N010(0)='1' AND  A(13)='0' AND D(17)='1' AND E( 9)='0' )then
          cVar2S19S28P013P063P064nsss(0) <='1';
          else
          cVar2S19S28P013P063P064nsss(0) <='0';
          end if;
        if(cVar1S20S28P017P019N016N010(0)='1' AND  A(13)='0' AND D(17)='0' AND D( 9)='1' )then
          cVar2S20S28P013N063P062nsss(0) <='1';
          else
          cVar2S20S28P013N063P062nsss(0) <='0';
          end if;
        if(cVar1S21S28P017P019N016N010(0)='1' AND  A(13)='1' AND E(17)='0' AND A(22)='1' )then
          cVar2S21S28P013P065P014nsss(0) <='1';
          else
          cVar2S21S28P013P065P014nsss(0) <='0';
          end if;
        if(cVar1S22S28P017P019P064P057(0)='1' AND  A(22)='1' AND D(20)='0' AND E(16)='0' )then
          cVar2S22S28P014P051P069nsss(0) <='1';
          else
          cVar2S22S28P014P051P069nsss(0) <='0';
          end if;
        if(cVar1S23S28P017P019P064P057(0)='1' AND  A(22)='0' AND A(20)='0' AND A(12)='1' )then
          cVar2S23S28P014P018P015nsss(0) <='1';
          else
          cVar2S23S28P014P018P015nsss(0) <='0';
          end if;
        if(cVar1S24S28P017P019P064P068(0)='1' AND  E(17)='1' )then
          cVar2S24S28P065nsss(0) <='1';
          else
          cVar2S24S28P065nsss(0) <='0';
          end if;
        if(cVar1S25S28P017P019P064P068(0)='1' AND  E(17)='0' AND E(16)='0' AND A(23)='0' )then
          cVar2S25S28N065P069P012nsss(0) <='1';
          else
          cVar2S25S28N065P069P012nsss(0) <='0';
          end if;
        if(cVar1S26S28P017P019P064N068(0)='1' AND  A(14)='1' AND B(20)='1' )then
          cVar2S26S28P011P036nsss(0) <='1';
          else
          cVar2S26S28P011P036nsss(0) <='0';
          end if;
        if(cVar1S27S28P017P019P064N068(0)='1' AND  A(14)='1' AND B(20)='0' AND A(21)='0' )then
          cVar2S27S28P011N036P016nsss(0) <='1';
          else
          cVar2S27S28P011N036P016nsss(0) <='0';
          end if;
        if(cVar1S0S29P017P013P011P032(0)='1' AND  B(21)='0' AND B(28)='0' )then
          cVar2S0S29P034P020nsss(0) <='1';
          else
          cVar2S0S29P034P020nsss(0) <='0';
          end if;
        if(cVar1S1S29P017P013P011P032(0)='1' AND  B(21)='1' AND A(12)='1' AND A(10)='1' )then
          cVar2S1S29P034P015P019nsss(0) <='1';
          else
          cVar2S1S29P034P015P019nsss(0) <='0';
          end if;
        if(cVar1S2S29P017P013N011P029(0)='1' AND  D(17)='1' AND B(21)='1' AND E(10)='0' )then
          cVar2S2S29P063P034P060nsss(0) <='1';
          else
          cVar2S2S29P063P034P060nsss(0) <='0';
          end if;
        if(cVar1S3S29P017P013N011P029(0)='1' AND  D(17)='1' AND B(21)='0' AND B(23)='1' )then
          cVar2S3S29P063N034P030nsss(0) <='1';
          else
          cVar2S3S29P063N034P030nsss(0) <='0';
          end if;
        if(cVar1S4S29P017P013N011P029(0)='1' AND  D(17)='0' AND E(17)='0' AND B(13)='0' )then
          cVar2S4S29N063P065P031nsss(0) <='1';
          else
          cVar2S4S29N063P065P031nsss(0) <='0';
          end if;
        if(cVar1S5S29P017P013N011P029(0)='1' AND  A(24)='1' )then
          cVar2S5S29P010nsss(0) <='1';
          else
          cVar2S5S29P010nsss(0) <='0';
          end if;
        if(cVar1S6S29P017P013P067P027(0)='1' AND  B(28)='0' AND A(21)='1' AND B(26)='0' )then
          cVar2S6S29P020P016P024nsss(0) <='1';
          else
          cVar2S6S29P020P016P024nsss(0) <='0';
          end if;
        if(cVar1S7S29P017P013P067P051(0)='1' AND  A(20)='1' AND E(16)='1' AND A(23)='1' )then
          cVar2S7S29P018P069P012nsss(0) <='1';
          else
          cVar2S7S29P018P069P012nsss(0) <='0';
          end if;
        if(cVar1S10S29N017P044N023N025(0)='1' AND  A(16)='0' AND B(27)='1' )then
          cVar2S10S29P007P022nsss(0) <='1';
          else
          cVar2S10S29P007P022nsss(0) <='0';
          end if;
        if(cVar1S11S29N017N044P055P057(0)='1' AND  B(23)='1' AND E( 8)='0' )then
          cVar2S11S29P030P068nsss(0) <='1';
          else
          cVar2S11S29P030P068nsss(0) <='0';
          end if;
        if(cVar1S12S29N017N044P055P057(0)='1' AND  B(23)='1' AND E( 8)='1' AND B(10)='0' )then
          cVar2S12S29P030P068P037nsss(0) <='1';
          else
          cVar2S12S29P030P068P037nsss(0) <='0';
          end if;
        if(cVar1S13S29N017N044P055P057(0)='1' AND  B(23)='0' AND B(13)='1' )then
          cVar2S13S29N030P031nsss(0) <='1';
          else
          cVar2S13S29N030P031nsss(0) <='0';
          end if;
        if(cVar1S14S29N017N044P055P057(0)='1' AND  B(23)='0' AND B(13)='0' AND B(22)='1' )then
          cVar2S14S29N030N031P032nsss(0) <='1';
          else
          cVar2S14S29N030N031P032nsss(0) <='0';
          end if;
        if(cVar1S15S29N017N044P055N057(0)='1' AND  E(17)='1' )then
          cVar2S15S29P065nsss(0) <='1';
          else
          cVar2S15S29P065nsss(0) <='0';
          end if;
        if(cVar1S16S29N017N044N055P041(0)='1' AND  B(28)='1' )then
          cVar2S16S29P020nsss(0) <='1';
          else
          cVar2S16S29P020nsss(0) <='0';
          end if;
        if(cVar1S17S29N017N044N055P041(0)='1' AND  B(28)='0' AND E(18)='0' AND B(18)='1' )then
          cVar2S17S29N020P061P021nsss(0) <='1';
          else
          cVar2S17S29N020P061P021nsss(0) <='0';
          end if;
        if(cVar1S18S29N017N044N055N041(0)='1' AND  B(20)='0' AND D(21)='1' )then
          cVar2S18S29P036P047nsss(0) <='1';
          else
          cVar2S18S29P036P047nsss(0) <='0';
          end if;
        if(cVar1S19S29N017N044N055N041(0)='1' AND  B(20)='1' AND A(21)='1' AND A(28)='0' )then
          cVar2S19S29P036P016P002nsss(0) <='1';
          else
          cVar2S19S29P036P016P002nsss(0) <='0';
          end if;
        if(cVar1S0S30P017P036P044P032(0)='1' AND  B(17)='1' )then
          cVar2S0S30P023nsss(0) <='1';
          else
          cVar2S0S30P023nsss(0) <='0';
          end if;
        if(cVar1S1S30P017P036P044P032(0)='1' AND  B(17)='0' AND B(27)='1' )then
          cVar2S1S30N023P022nsss(0) <='1';
          else
          cVar2S1S30N023P022nsss(0) <='0';
          end if;
        if(cVar1S2S30P017P036P044P032(0)='1' AND  B(17)='0' AND B(27)='0' AND D( 9)='0' )then
          cVar2S2S30N023N022P062nsss(0) <='1';
          else
          cVar2S2S30N023N022P062nsss(0) <='0';
          end if;
        if(cVar1S3S30P017P036N044P041(0)='1' AND  B(28)='1' )then
          cVar2S3S30P020nsss(0) <='1';
          else
          cVar2S3S30P020nsss(0) <='0';
          end if;
        if(cVar1S4S30P017P036N044P041(0)='1' AND  B(28)='0' AND D(18)='0' AND A(21)='0' )then
          cVar2S4S30N020P059P016nsss(0) <='1';
          else
          cVar2S4S30N020P059P016nsss(0) <='0';
          end if;
        if(cVar1S5S30P017P036N044N041(0)='1' AND  E( 9)='1' AND D( 9)='1' )then
          cVar2S5S30P064P062nsss(0) <='1';
          else
          cVar2S5S30P064P062nsss(0) <='0';
          end if;
        if(cVar1S6S30P017P036N044N041(0)='1' AND  E( 9)='1' AND D( 9)='0' AND D( 8)='1' )then
          cVar2S6S30P064N062P066nsss(0) <='1';
          else
          cVar2S6S30P064N062P066nsss(0) <='0';
          end if;
        if(cVar1S7S30P017P036N044N041(0)='1' AND  E( 9)='0' AND D( 9)='0' )then
          cVar2S7S30N064P062nsss(0) <='1';
          else
          cVar2S7S30N064P062nsss(0) <='0';
          end if;
        if(cVar1S8S30P017P036P004P013(0)='1' AND  B(13)='1' )then
          cVar2S8S30P031nsss(0) <='1';
          else
          cVar2S8S30P031nsss(0) <='0';
          end if;
        if(cVar1S9S30P017P036P004P013(0)='1' AND  B(13)='0' AND D( 9)='0' AND B(12)='1' )then
          cVar2S9S30N031P062P033nsss(0) <='1';
          else
          cVar2S9S30N031P062P033nsss(0) <='0';
          end if;
        if(cVar1S10S30P017P036P004N013(0)='1' AND  E(12)='1' AND D(12)='1' )then
          cVar2S10S30P052P050nsss(0) <='1';
          else
          cVar2S10S30P052P050nsss(0) <='0';
          end if;
        if(cVar1S11S30P017P036P004N013(0)='1' AND  E(12)='0' AND D( 9)='1' AND A(15)='0' )then
          cVar2S11S30N052P062P009nsss(0) <='1';
          else
          cVar2S11S30N052P062P009nsss(0) <='0';
          end if;
        if(cVar1S12S30P017P036P004P006(0)='1' AND  A(22)='0' AND D(16)='0' )then
          cVar2S12S30P014P067nsss(0) <='1';
          else
          cVar2S12S30P014P067nsss(0) <='0';
          end if;
        if(cVar1S13S30P017P044P063P043(0)='1' AND  A(17)='0' AND A(14)='0' AND A(27)='0' )then
          cVar2S13S30P005P011P004nsss(0) <='1';
          else
          cVar2S13S30P005P011P004nsss(0) <='0';
          end if;
        if(cVar1S14S30P017P044P063P043(0)='1' AND  A(17)='0' AND A(14)='1' AND A(23)='1' )then
          cVar2S14S30P005P011P012nsss(0) <='1';
          else
          cVar2S14S30P005P011P012nsss(0) <='0';
          end if;
        if(cVar1S15S30P017P044N063P065(0)='1' AND  A(14)='1' AND A(28)='0' AND B(11)='0' )then
          cVar2S15S30P011P002P035nsss(0) <='1';
          else
          cVar2S15S30P011P002P035nsss(0) <='0';
          end if;
        if(cVar1S16S30P017P044N063P065(0)='1' AND  A(14)='0' AND B(25)='1' AND E( 8)='0' )then
          cVar2S16S30N011P026P068nsss(0) <='1';
          else
          cVar2S16S30N011P026P068nsss(0) <='0';
          end if;
        if(cVar1S17S30P017P044N063P065(0)='1' AND  A(14)='0' AND B(25)='0' AND D(10)='1' )then
          cVar2S17S30N011N026P058nsss(0) <='1';
          else
          cVar2S17S30N011N026P058nsss(0) <='0';
          end if;
        if(cVar1S18S30P017P044N063P065(0)='1' AND  B(21)='0' AND A(25)='0' AND D( 9)='1' )then
          cVar2S18S30P034P008P062nsss(0) <='1';
          else
          cVar2S18S30P034P008P062nsss(0) <='0';
          end if;
        if(cVar1S19S30P017P044P034P014(0)='1' AND  D(13)='0' AND A(12)='1' )then
          cVar2S19S30P046P015nsss(0) <='1';
          else
          cVar2S19S30P046P015nsss(0) <='0';
          end if;
        if(cVar1S0S31P033P054P061P032(0)='1' AND  A(22)='0' AND D(18)='1' )then
          cVar2S0S31P014P059nsss(0) <='1';
          else
          cVar2S0S31P014P059nsss(0) <='0';
          end if;
        if(cVar1S1S31P033P054N061P063(0)='1' AND  B(21)='0' AND A(27)='0' )then
          cVar2S1S31P034P004nsss(0) <='1';
          else
          cVar2S1S31P034P004nsss(0) <='0';
          end if;
        if(cVar1S2S31P033P054N061P063(0)='1' AND  D(16)='1' AND A(12)='1' )then
          cVar2S2S31P067P015nsss(0) <='1';
          else
          cVar2S2S31P067P015nsss(0) <='0';
          end if;
        if(cVar1S3S31N033P061P029P011(0)='1' AND  A(15)='0' )then
          cVar2S3S31P009nsss(0) <='1';
          else
          cVar2S3S31P009nsss(0) <='0';
          end if;
        if(cVar1S4S31N033P061P029N011(0)='1' AND  E(12)='1' )then
          cVar2S4S31P052nsss(0) <='1';
          else
          cVar2S4S31P052nsss(0) <='0';
          end if;
        if(cVar1S5S31N033P061P029N011(0)='1' AND  E(12)='0' AND A(25)='1' )then
          cVar2S5S31N052P008nsss(0) <='1';
          else
          cVar2S5S31N052P008nsss(0) <='0';
          end if;
        if(cVar1S6S31N033P061P029N011(0)='1' AND  E(12)='0' AND A(25)='0' AND A(24)='1' )then
          cVar2S6S31N052N008P010nsss(0) <='1';
          else
          cVar2S6S31N052N008P010nsss(0) <='0';
          end if;
        if(cVar1S7S31N033P061N029P040(0)='1' AND  B(18)='1' )then
          cVar2S7S31P021nsss(0) <='1';
          else
          cVar2S7S31P021nsss(0) <='0';
          end if;
        if(cVar1S8S31N033P061N029P040(0)='1' AND  B(18)='0' AND A(28)='1' )then
          cVar2S8S31N021P002nsss(0) <='1';
          else
          cVar2S8S31N021P002nsss(0) <='0';
          end if;
        if(cVar1S9S31N033P061N029P040(0)='1' AND  B(18)='0' AND A(28)='0' AND A(27)='1' )then
          cVar2S9S31N021N002P004nsss(0) <='1';
          else
          cVar2S9S31N021N002P004nsss(0) <='0';
          end if;
        if(cVar1S10S31N033P061N029N040(0)='1' AND  D(15)='0' AND E(14)='1' AND D(14)='1' )then
          cVar2S10S31P038P044P042nsss(0) <='1';
          else
          cVar2S10S31P038P044P042nsss(0) <='0';
          end if;
        if(cVar1S11S31N033P061N029N040(0)='1' AND  D(15)='1' AND A(24)='1' )then
          cVar2S11S31P038P010nsss(0) <='1';
          else
          cVar2S11S31P038P010nsss(0) <='0';
          end if;
        if(cVar1S12S31N033P061P059P032(0)='1' AND  E( 9)='0' )then
          cVar2S12S31P064nsss(0) <='1';
          else
          cVar2S12S31P064nsss(0) <='0';
          end if;
        if(cVar1S13S31N033P061P059P032(0)='1' AND  E( 9)='1' AND D(17)='1' )then
          cVar2S13S31P064P063nsss(0) <='1';
          else
          cVar2S13S31P064P063nsss(0) <='0';
          end if;
        if(cVar1S14S31N033P061P059P032(0)='1' AND  E(16)='1' )then
          cVar2S14S31P069nsss(0) <='1';
          else
          cVar2S14S31P069nsss(0) <='0';
          end if;
        if(cVar1S15S31N033P061P059P032(0)='1' AND  E(16)='0' AND E( 9)='1' AND A(11)='0' )then
          cVar2S15S31N069P064P017nsss(0) <='1';
          else
          cVar2S15S31N069P064P017nsss(0) <='0';
          end if;
        if(cVar1S16S31N033P061N059P018(0)='1' AND  B(21)='0' AND A(25)='0' AND A(12)='1' )then
          cVar2S16S31P034P008P015nsss(0) <='1';
          else
          cVar2S16S31P034P008P015nsss(0) <='0';
          end if;
        if(cVar1S17S31N033P061N059N018(0)='1' AND  D(17)='1' AND A(22)='0' AND E(16)='0' )then
          cVar2S17S31P063P014P069nsss(0) <='1';
          else
          cVar2S17S31P063P014P069nsss(0) <='0';
          end if;
        if(cVar1S0S32P061P033P060P064(0)='1' AND  E( 8)='1' AND A(17)='0' )then
          cVar2S0S32P068P005nsss(0) <='1';
          else
          cVar2S0S32P068P005nsss(0) <='0';
          end if;
        if(cVar1S1S32P061P033P060P064(0)='1' AND  E( 8)='0' AND D(19)='1' )then
          cVar2S1S32N068P055nsss(0) <='1';
          else
          cVar2S1S32N068P055nsss(0) <='0';
          end if;
        if(cVar1S2S32P061P033P060P064(0)='1' AND  E( 8)='0' AND D(19)='0' AND D(11)='1' )then
          cVar2S2S32N068N055P054nsss(0) <='1';
          else
          cVar2S2S32N068N055P054nsss(0) <='0';
          end if;
        if(cVar1S3S32P061P033P060N064(0)='1' AND  D( 9)='0' AND E(23)='1' AND D(23)='1' )then
          cVar2S3S32P062P041P039nsss(0) <='1';
          else
          cVar2S3S32P062P041P039nsss(0) <='0';
          end if;
        if(cVar1S4S32P061P033P060N064(0)='1' AND  D( 9)='0' AND E(23)='0' )then
          cVar2S4S32P062N041psss(0) <='1';
          else
          cVar2S4S32P062N041psss(0) <='0';
          end if;
        if(cVar1S6S32P061P033P060N032(0)='1' AND  B(11)='1' AND B(21)='0' AND A(13)='0' )then
          cVar2S6S32P035P034P013nsss(0) <='1';
          else
          cVar2S6S32P035P034P013nsss(0) <='0';
          end if;
        if(cVar1S7S32P061P033P060N032(0)='1' AND  B(11)='0' AND E(17)='0' AND D( 8)='1' )then
          cVar2S7S32N035P065P066nsss(0) <='1';
          else
          cVar2S7S32N035P065P066nsss(0) <='0';
          end if;
        if(cVar1S8S32P061P033P065P060(0)='1' AND  A(13)='1' AND A(11)='0' )then
          cVar2S8S32P013P017nsss(0) <='1';
          else
          cVar2S8S32P013P017nsss(0) <='0';
          end if;
        if(cVar1S9S32P061P033P065P060(0)='1' AND  A(13)='0' AND D(16)='0' AND A(22)='1' )then
          cVar2S9S32N013P067P014nsss(0) <='1';
          else
          cVar2S9S32N013P067P014nsss(0) <='0';
          end if;
        if(cVar1S10S32P061P033P065N060(0)='1' AND  B(21)='0' AND D(23)='1' )then
          cVar2S10S32P034P039nsss(0) <='1';
          else
          cVar2S10S32P034P039nsss(0) <='0';
          end if;
        if(cVar1S11S32P061P033P065P019(0)='1' AND  A(21)='1' AND B(21)='1' )then
          cVar2S11S32P016P034nsss(0) <='1';
          else
          cVar2S11S32P016P034nsss(0) <='0';
          end if;
        if(cVar1S12S32P061P059P032P064(0)='1' AND  B(12)='1' AND D(10)='0' )then
          cVar2S12S32P033P058nsss(0) <='1';
          else
          cVar2S12S32P033P058nsss(0) <='0';
          end if;
        if(cVar1S13S32P061P059P032P064(0)='1' AND  B(12)='0' AND B(21)='1' )then
          cVar2S13S32N033P034nsss(0) <='1';
          else
          cVar2S13S32N033P034nsss(0) <='0';
          end if;
        if(cVar1S14S32P061P059P032P064(0)='1' AND  B(12)='0' AND B(21)='0' AND B(11)='1' )then
          cVar2S14S32N033N034P035nsss(0) <='1';
          else
          cVar2S14S32N033N034P035nsss(0) <='0';
          end if;
        if(cVar1S15S32P061P059P032P064(0)='1' AND  A(13)='0' AND D(17)='1' )then
          cVar2S15S32P013P063nsss(0) <='1';
          else
          cVar2S15S32P013P063nsss(0) <='0';
          end if;
        if(cVar1S16S32P061P059P032P067(0)='1' AND  B(21)='0' )then
          cVar2S16S32P034nsss(0) <='1';
          else
          cVar2S16S32P034nsss(0) <='0';
          end if;
        if(cVar1S17S32P061P059P032N067(0)='1' AND  E( 9)='1' )then
          cVar2S17S32P064nsss(0) <='1';
          else
          cVar2S17S32P064nsss(0) <='0';
          end if;
        if(cVar1S18S32P061P059P032N067(0)='1' AND  E( 9)='0' AND E( 8)='1' AND A(10)='1' )then
          cVar2S18S32N064P068P019nsss(0) <='1';
          else
          cVar2S18S32N064P068P019nsss(0) <='0';
          end if;
        if(cVar1S19S32P061N059P018P034(0)='1' AND  A(25)='0' AND A(12)='1' AND A(22)='0' )then
          cVar2S19S32P008P015P014nsss(0) <='1';
          else
          cVar2S19S32P008P015P014nsss(0) <='0';
          end if;
        if(cVar1S20S32P061N059P018P034(0)='1' AND  A(25)='0' AND A(12)='0' AND A(22)='1' )then
          cVar2S20S32P008N015P014nsss(0) <='1';
          else
          cVar2S20S32P008N015P014nsss(0) <='0';
          end if;
        if(cVar1S21S32P061N059N018P063(0)='1' AND  A(14)='0' AND A(22)='0' AND A(21)='1' )then
          cVar2S21S32P011P014P016nsss(0) <='1';
          else
          cVar2S21S32P011P014P016nsss(0) <='0';
          end if;
        if(cVar1S0S33P062P013P054P037(0)='1' AND  A(17)='0' AND D(12)='0' )then
          cVar2S0S33P005P050nsss(0) <='1';
          else
          cVar2S0S33P005P050nsss(0) <='0';
          end if;
        if(cVar1S1S33P062P013P054N037(0)='1' AND  B(11)='1' AND A(15)='0' )then
          cVar2S1S33P035P009nsss(0) <='1';
          else
          cVar2S1S33P035P009nsss(0) <='0';
          end if;
        if(cVar1S2S33P062P013P054N037(0)='1' AND  B(11)='0' AND A(19)='0' AND E(20)='1' )then
          cVar2S2S33N035P001P053nsss(0) <='1';
          else
          cVar2S2S33N035P001P053nsss(0) <='0';
          end if;
        if(cVar1S3S33P062P013P054P068(0)='1' AND  A(12)='0' AND A(11)='0' )then
          cVar2S3S33P015P017nsss(0) <='1';
          else
          cVar2S3S33P015P017nsss(0) <='0';
          end if;
        if(cVar1S4S33P062P013P067P059(0)='1' AND  B(23)='0' AND A(10)='0' AND E( 8)='0' )then
          cVar2S4S33P030P019P068nsss(0) <='1';
          else
          cVar2S4S33P030P019P068nsss(0) <='0';
          end if;
        if(cVar1S5S33P062P013P067P059(0)='1' AND  B(23)='0' AND A(10)='1' AND E( 9)='1' )then
          cVar2S5S33P030P019P064nsss(0) <='1';
          else
          cVar2S5S33P030P019P064nsss(0) <='0';
          end if;
        if(cVar1S6S33P062P013P067P011(0)='1' AND  A(26)='0' AND A(24)='0' AND A(10)='0' )then
          cVar2S6S33P006P010P019nsss(0) <='1';
          else
          cVar2S6S33P006P010P019nsss(0) <='0';
          end if;
        if(cVar1S8S33N062P041N020P035(0)='1' AND  D(20)='0' AND B(18)='1' )then
          cVar2S8S33P051P021nsss(0) <='1';
          else
          cVar2S8S33P051P021nsss(0) <='0';
          end if;
        if(cVar1S9S33N062P041N020P035(0)='1' AND  D(20)='0' AND B(18)='0' AND A(25)='0' )then
          cVar2S9S33P051N021P008nsss(0) <='1';
          else
          cVar2S9S33P051N021P008nsss(0) <='0';
          end if;
        if(cVar1S10S33N062N041P033P061(0)='1' AND  B(22)='0' AND A(12)='1' )then
          cVar2S10S33P032P015nsss(0) <='1';
          else
          cVar2S10S33P032P015nsss(0) <='0';
          end if;
        if(cVar1S11S33N062N041P033P061(0)='1' AND  B(22)='0' AND A(12)='0' AND A(13)='1' )then
          cVar2S11S33P032N015P013nsss(0) <='1';
          else
          cVar2S11S33P032N015P013nsss(0) <='0';
          end if;
        if(cVar1S12S33N062N041P033N061(0)='1' AND  D(17)='0' AND B(21)='0' AND E(11)='0' )then
          cVar2S12S33P063P034P056nsss(0) <='1';
          else
          cVar2S12S33P063P034P056nsss(0) <='0';
          end if;
        if(cVar1S13S33N062N041P033N061(0)='1' AND  D(17)='0' AND B(21)='1' AND A(13)='1' )then
          cVar2S13S33P063P034P013nsss(0) <='1';
          else
          cVar2S13S33P063P034P013nsss(0) <='0';
          end if;
        if(cVar1S14S33N062N041P033N061(0)='1' AND  D(17)='1' AND D(16)='1' )then
          cVar2S14S33P063P067nsss(0) <='1';
          else
          cVar2S14S33P063P067nsss(0) <='0';
          end if;
        if(cVar1S15S33N062N041N033P039(0)='1' AND  A(14)='1' AND B(14)='1' )then
          cVar2S15S33P011P029nsss(0) <='1';
          else
          cVar2S15S33P011P029nsss(0) <='0';
          end if;
        if(cVar1S16S33N062N041N033P039(0)='1' AND  A(14)='1' AND B(14)='0' AND E(16)='0' )then
          cVar2S16S33P011N029P069nsss(0) <='1';
          else
          cVar2S16S33P011N029P069nsss(0) <='0';
          end if;
        if(cVar1S17S33N062N041N033P039(0)='1' AND  A(14)='0' AND E(14)='1' )then
          cVar2S17S33N011P044nsss(0) <='1';
          else
          cVar2S17S33N011P044nsss(0) <='0';
          end if;
        if(cVar1S18S33N062N041N033P039(0)='1' AND  A(25)='0' AND A(23)='0' AND A(22)='1' )then
          cVar2S18S33P008P012P014nsss(0) <='1';
          else
          cVar2S18S33P008P012P014nsss(0) <='0';
          end if;
        if(cVar1S0S34P011P029P062P003(0)='1' AND  A(17)='0' )then
          cVar2S0S34P005nsss(0) <='1';
          else
          cVar2S0S34P005nsss(0) <='0';
          end if;
        if(cVar1S1S34P011P029P062P003(0)='1' AND  A(17)='1' AND A(11)='0' )then
          cVar2S1S34P005P017nsss(0) <='1';
          else
          cVar2S1S34P005P017nsss(0) <='0';
          end if;
        if(cVar1S2S34P011P029P062P003(0)='1' AND  A(21)='1' AND A(20)='0' )then
          cVar2S2S34P016P018nsss(0) <='1';
          else
          cVar2S2S34P016P018nsss(0) <='0';
          end if;
        if(cVar1S3S34P011P029N062P059(0)='1' AND  E(16)='1' AND D(20)='0' )then
          cVar2S3S34P069P051nsss(0) <='1';
          else
          cVar2S3S34P069P051nsss(0) <='0';
          end if;
        if(cVar1S4S34P011P029N062P059(0)='1' AND  E(16)='0' AND B(22)='0' AND E(18)='1' )then
          cVar2S4S34N069P032P061nsss(0) <='1';
          else
          cVar2S4S34N069P032P061nsss(0) <='0';
          end if;
        if(cVar1S5S34P011P029N062P059(0)='1' AND  E(16)='0' AND B(22)='1' AND E(18)='0' )then
          cVar2S5S34N069P032P061nsss(0) <='1';
          else
          cVar2S5S34N069P032P061nsss(0) <='0';
          end if;
        if(cVar1S6S34P011P029N062N059(0)='1' AND  E(18)='0' AND A(27)='1' )then
          cVar2S6S34P061P004nsss(0) <='1';
          else
          cVar2S6S34P061P004nsss(0) <='0';
          end if;
        if(cVar1S7S34P011P029N062N059(0)='1' AND  E(18)='0' AND A(27)='0' AND A(12)='0' )then
          cVar2S7S34P061N004P015nsss(0) <='1';
          else
          cVar2S7S34P061N004P015nsss(0) <='0';
          end if;
        if(cVar1S8S34P011P029N062N059(0)='1' AND  E(18)='1' AND A(20)='1' AND D(17)='0' )then
          cVar2S8S34P061P018P063nsss(0) <='1';
          else
          cVar2S8S34P061P018P063nsss(0) <='0';
          end if;
        if(cVar1S10S34P011P029N052P004(0)='1' AND  B(12)='0' AND A(24)='1' AND A(10)='0' )then
          cVar2S10S34P033P010P019nsss(0) <='1';
          else
          cVar2S10S34P033P010P019nsss(0) <='0';
          end if;
        if(cVar1S11S34P011P029N052P004(0)='1' AND  B(12)='0' AND A(24)='0' AND A(25)='1' )then
          cVar2S11S34P033N010P008nsss(0) <='1';
          else
          cVar2S11S34P033N010P008nsss(0) <='0';
          end if;
        if(cVar1S12S34P011P013P032P029(0)='1' AND  A(10)='0' )then
          cVar2S12S34P019nsss(0) <='1';
          else
          cVar2S12S34P019nsss(0) <='0';
          end if;
        if(cVar1S13S34P011P013P032N029(0)='1' AND  A(18)='0' AND A(12)='1' AND A(26)='0' )then
          cVar2S13S34P003P015P006nsss(0) <='1';
          else
          cVar2S13S34P003P015P006nsss(0) <='0';
          end if;
        if(cVar1S14S34P011P013P032N029(0)='1' AND  A(18)='0' AND A(12)='0' AND B(13)='1' )then
          cVar2S14S34P003N015P031nsss(0) <='1';
          else
          cVar2S14S34P003N015P031nsss(0) <='0';
          end if;
        if(cVar1S15S34P011P013P032N029(0)='1' AND  A(18)='1' AND A(12)='1' AND A(20)='0' )then
          cVar2S15S34P003P015P018nsss(0) <='1';
          else
          cVar2S15S34P003P015P018nsss(0) <='0';
          end if;
        if(cVar1S16S34P011P013P004P008(0)='1' AND  B(18)='0' AND A(16)='1' AND A(21)='1' )then
          cVar2S16S34P021P007P016nsss(0) <='1';
          else
          cVar2S16S34P021P007P016nsss(0) <='0';
          end if;
        if(cVar1S17S34P011P013P004P008(0)='1' AND  E(16)='0' AND A(26)='0' AND E(17)='1' )then
          cVar2S17S34P069P006P065nsss(0) <='1';
          else
          cVar2S17S34P069P006P065nsss(0) <='0';
          end if;
        if(cVar1S0S35P015P022P034P054(0)='1' AND  D(17)='0' AND D( 8)='1' )then
          cVar2S0S35P063P066nsss(0) <='1';
          else
          cVar2S0S35P063P066nsss(0) <='0';
          end if;
        if(cVar1S1S35P015P022P034P054(0)='1' AND  D(17)='0' AND D( 8)='0' AND E(17)='0' )then
          cVar2S1S35P063N066P065nsss(0) <='1';
          else
          cVar2S1S35P063N066P065nsss(0) <='0';
          end if;
        if(cVar1S2S35P015P022P034P054(0)='1' AND  D(17)='1' AND B(11)='1' AND D(16)='0' )then
          cVar2S2S35P063P035P067nsss(0) <='1';
          else
          cVar2S2S35P063P035P067nsss(0) <='0';
          end if;
        if(cVar1S3S35P015P022P034P054(0)='1' AND  A(28)='0' AND E(11)='1' AND B(20)='1' )then
          cVar2S3S35P002P056P036nsss(0) <='1';
          else
          cVar2S3S35P002P056P036nsss(0) <='0';
          end if;
        if(cVar1S4S35P015P022P034P044(0)='1' AND  D(22)='0' AND D(17)='1' AND A(10)='0' )then
          cVar2S4S35P043P063P019nsss(0) <='1';
          else
          cVar2S4S35P043P063P019nsss(0) <='0';
          end if;
        if(cVar1S6S35N015P064P043P033(0)='1' AND  E( 8)='1' AND B(26)='0' )then
          cVar2S6S35P068P024nsss(0) <='1';
          else
          cVar2S6S35P068P024nsss(0) <='0';
          end if;
        if(cVar1S7S35N015P064P043P033(0)='1' AND  E( 8)='0' AND D(19)='1' )then
          cVar2S7S35N068P055nsss(0) <='1';
          else
          cVar2S7S35N068P055nsss(0) <='0';
          end if;
        if(cVar1S8S35N015P064P043P033(0)='1' AND  E( 8)='0' AND D(19)='0' AND A(22)='1' )then
          cVar2S8S35N068N055P014nsss(0) <='1';
          else
          cVar2S8S35N068N055P014nsss(0) <='0';
          end if;
        if(cVar1S9S35N015P064P043P033(0)='1' AND  E(10)='1' )then
          cVar2S9S35P060nsss(0) <='1';
          else
          cVar2S9S35P060nsss(0) <='0';
          end if;
        if(cVar1S10S35N015N064P068P034(0)='1' AND  D(17)='1' AND A(23)='0' )then
          cVar2S10S35P063P012nsss(0) <='1';
          else
          cVar2S10S35P063P012nsss(0) <='0';
          end if;
        if(cVar1S11S35N015N064P068P034(0)='1' AND  D(17)='1' AND A(23)='1' AND A(22)='0' )then
          cVar2S11S35P063P012P014nsss(0) <='1';
          else
          cVar2S11S35P063P012P014nsss(0) <='0';
          end if;
        if(cVar1S12S35N015N064P068P034(0)='1' AND  D(17)='0' AND E(17)='0' AND B(11)='0' )then
          cVar2S12S35N063P065P035nsss(0) <='1';
          else
          cVar2S12S35N063P065P035nsss(0) <='0';
          end if;
        if(cVar1S13S35N015N064P068N034(0)='1' AND  B(28)='1' AND D(23)='1' )then
          cVar2S13S35P020P039nsss(0) <='1';
          else
          cVar2S13S35P020P039nsss(0) <='0';
          end if;
        if(cVar1S14S35N015N064P068N034(0)='1' AND  B(28)='1' AND D(23)='0' AND B(11)='0' )then
          cVar2S14S35P020N039P035nsss(0) <='1';
          else
          cVar2S14S35P020N039P035nsss(0) <='0';
          end if;
        if(cVar1S15S35N015N064P068N034(0)='1' AND  B(28)='0' AND A(14)='1' )then
          cVar2S15S35N020P011nsss(0) <='1';
          else
          cVar2S15S35N020P011nsss(0) <='0';
          end if;
        if(cVar1S16S35N015N064P068N034(0)='1' AND  B(28)='0' AND A(14)='0' AND A(26)='1' )then
          cVar2S16S35N020N011P006nsss(0) <='1';
          else
          cVar2S16S35N020N011P006nsss(0) <='0';
          end if;
        if(cVar1S17S35N015N064P068P011(0)='1' AND  A(25)='1' AND A(23)='0' )then
          cVar2S17S35P008P012nsss(0) <='1';
          else
          cVar2S17S35P008P012nsss(0) <='0';
          end if;
        if(cVar1S18S35N015N064P068P011(0)='1' AND  A(25)='0' AND D( 9)='0' AND D(22)='1' )then
          cVar2S18S35N008P062P043nsss(0) <='1';
          else
          cVar2S18S35N008P062P043nsss(0) <='0';
          end if;
        if(cVar1S19S35N015N064P068P011(0)='1' AND  A(25)='0' AND D( 9)='1' AND E(10)='1' )then
          cVar2S19S35N008P062P060nsss(0) <='1';
          else
          cVar2S19S35N008P062P060nsss(0) <='0';
          end if;
        if(cVar1S20S35N015N064P068P011(0)='1' AND  E(17)='0' AND B(11)='1' )then
          cVar2S20S35P065P035nsss(0) <='1';
          else
          cVar2S20S35P065P035nsss(0) <='0';
          end if;
        if(cVar1S0S36P011P015P065P063(0)='1' AND  E(10)='0' AND D( 8)='0' )then
          cVar2S0S36P060P066nsss(0) <='1';
          else
          cVar2S0S36P060P066nsss(0) <='0';
          end if;
        if(cVar1S1S36P011P015P065P063(0)='1' AND  E(10)='0' AND D( 8)='1' AND A(23)='1' )then
          cVar2S1S36P060P066P012nsss(0) <='1';
          else
          cVar2S1S36P060P066P012nsss(0) <='0';
          end if;
        if(cVar1S2S36P011P015P065P063(0)='1' AND  E(10)='1' AND A(22)='1' )then
          cVar2S2S36P060P014nsss(0) <='1';
          else
          cVar2S2S36P060P014nsss(0) <='0';
          end if;
        if(cVar1S3S36P011P015P065N063(0)='1' AND  A(21)='0' AND D(16)='1' )then
          cVar2S3S36P016P067nsss(0) <='1';
          else
          cVar2S3S36P016P067nsss(0) <='0';
          end if;
        if(cVar1S4S36P011P015P065N063(0)='1' AND  A(21)='0' AND D(16)='0' AND E( 8)='1' )then
          cVar2S4S36P016N067P068nsss(0) <='1';
          else
          cVar2S4S36P016N067P068nsss(0) <='0';
          end if;
        if(cVar1S5S36P011P015P065N063(0)='1' AND  A(21)='1' AND D( 8)='1' )then
          cVar2S5S36P016P066nsss(0) <='1';
          else
          cVar2S5S36P016P066nsss(0) <='0';
          end if;
        if(cVar1S6S36P011P015N065P063(0)='1' AND  B(21)='0' AND B(14)='0' )then
          cVar2S6S36P034P029nsss(0) <='1';
          else
          cVar2S6S36P034P029nsss(0) <='0';
          end if;
        if(cVar1S7S36P011P015N065P063(0)='1' AND  B(21)='0' AND B(14)='1' AND E(12)='1' )then
          cVar2S7S36P034P029P052nsss(0) <='1';
          else
          cVar2S7S36P034P029P052nsss(0) <='0';
          end if;
        if(cVar1S8S36P011P015N065P063(0)='1' AND  B(21)='1' AND B(14)='1' )then
          cVar2S8S36P034P029nsss(0) <='1';
          else
          cVar2S8S36P034P029nsss(0) <='0';
          end if;
        if(cVar1S9S36P011P015N065P063(0)='1' AND  B(21)='1' AND B(14)='0' AND E(18)='1' )then
          cVar2S9S36P034N029P061nsss(0) <='1';
          else
          cVar2S9S36P034N029P061nsss(0) <='0';
          end if;
        if(cVar1S10S36P011P015N065P063(0)='1' AND  E( 9)='1' AND D( 8)='0' )then
          cVar2S10S36P064P066nsss(0) <='1';
          else
          cVar2S10S36P064P066nsss(0) <='0';
          end if;
        if(cVar1S11S36P011P015N065P063(0)='1' AND  E( 9)='0' AND A(13)='1' AND A(10)='0' )then
          cVar2S11S36N064P013P019nsss(0) <='1';
          else
          cVar2S11S36N064P013P019nsss(0) <='0';
          end if;
        if(cVar1S12S36P011P015P022P059(0)='1' AND  A(27)='0' AND B(26)='0' AND A(23)='0' )then
          cVar2S12S36P004P024P012nsss(0) <='1';
          else
          cVar2S12S36P004P024P012nsss(0) <='0';
          end if;
        if(cVar1S13S36P011P015P022N059(0)='1' AND  A(13)='1' AND E(23)='0' AND D( 9)='0' )then
          cVar2S13S36P013P041P062nsss(0) <='1';
          else
          cVar2S13S36P013P041P062nsss(0) <='0';
          end if;
        if(cVar1S14S36P011P015P022N059(0)='1' AND  A(13)='0' AND B(13)='0' AND E(23)='1' )then
          cVar2S14S36N013P031P041nsss(0) <='1';
          else
          cVar2S14S36N013P031P041nsss(0) <='0';
          end if;
        if(cVar1S15S36P011P015P022N059(0)='1' AND  A(13)='0' AND B(13)='1' AND D( 8)='1' )then
          cVar2S15S36N013P031P066nsss(0) <='1';
          else
          cVar2S15S36N013P031P066nsss(0) <='0';
          end if;
        if(cVar1S17S36P011P004P029N054(0)='1' AND  D(20)='1' )then
          cVar2S17S36P051nsss(0) <='1';
          else
          cVar2S17S36P051nsss(0) <='0';
          end if;
        if(cVar1S18S36P011P004P029N054(0)='1' AND  D(20)='0' AND E(12)='1' )then
          cVar2S18S36N051P052nsss(0) <='1';
          else
          cVar2S18S36N051P052nsss(0) <='0';
          end if;
        if(cVar1S19S36P011P004N029P002(0)='1' AND  B(18)='0' AND D(23)='0' AND B(24)='1' )then
          cVar2S19S36P021P039P028nsss(0) <='1';
          else
          cVar2S19S36P021P039P028nsss(0) <='0';
          end if;
        if(cVar1S20S36P011P004N029P002(0)='1' AND  A(29)='0' AND E(17)='0' AND A(12)='1' )then
          cVar2S20S36P000P065P015nsss(0) <='1';
          else
          cVar2S20S36P000P065P015nsss(0) <='0';
          end if;
        if(cVar1S21S36P011P004P000P056(0)='1' AND  A(18)='0' AND A(25)='0' AND E( 9)='1' )then
          cVar2S21S36P003P008P064nsss(0) <='1';
          else
          cVar2S21S36P003P008P064nsss(0) <='0';
          end if;
        if(cVar1S0S37P015P031P022P006(0)='1' AND  E(22)='0' AND E(20)='1' AND A(29)='0' )then
          cVar2S0S37P045P053P000nsss(0) <='1';
          else
          cVar2S0S37P045P053P000nsss(0) <='0';
          end if;
        if(cVar1S1S37P015P031P022P006(0)='1' AND  E(22)='0' AND E(20)='0' AND D(20)='0' )then
          cVar2S1S37P045N053P051nsss(0) <='1';
          else
          cVar2S1S37P045N053P051nsss(0) <='0';
          end if;
        if(cVar1S2S37P015P031P022P006(0)='1' AND  E(22)='1' AND E( 8)='1' )then
          cVar2S2S37P045P068nsss(0) <='1';
          else
          cVar2S2S37P045P068nsss(0) <='0';
          end if;
        if(cVar1S3S37P015P031P022P006(0)='1' AND  B(20)='0' AND D(11)='0' AND A(21)='0' )then
          cVar2S3S37P036P054P016nsss(0) <='1';
          else
          cVar2S3S37P036P054P016nsss(0) <='0';
          end if;
        if(cVar1S5S37P015P031P004P030(0)='1' AND  A(24)='1' )then
          cVar2S5S37P010nsss(0) <='1';
          else
          cVar2S5S37P010nsss(0) <='0';
          end if;
        if(cVar1S6S37P015P031P004P030(0)='1' AND  A(24)='0' AND D(18)='1' )then
          cVar2S6S37N010P059nsss(0) <='1';
          else
          cVar2S6S37N010P059nsss(0) <='0';
          end if;
        if(cVar1S8S37N015P065P007N052(0)='1' AND  D(12)='0' AND E(10)='0' AND D(17)='1' )then
          cVar2S8S37P050P060P063nsss(0) <='1';
          else
          cVar2S8S37P050P060P063nsss(0) <='0';
          end if;
        if(cVar1S9S37N015P065P007N052(0)='1' AND  D(12)='0' AND E(10)='1' AND D( 9)='1' )then
          cVar2S9S37P050P060P062nsss(0) <='1';
          else
          cVar2S9S37P050P060P062nsss(0) <='0';
          end if;
        if(cVar1S10S37N015P065P007P009(0)='1' AND  A(24)='0' AND A(20)='1' )then
          cVar2S10S37P010P018nsss(0) <='1';
          else
          cVar2S10S37P010P018nsss(0) <='0';
          end if;
        if(cVar1S12S37N015N065P022N043(0)='1' AND  B(26)='0' AND E(16)='0' AND A(27)='1' )then
          cVar2S12S37P024P069P004nsss(0) <='1';
          else
          cVar2S12S37P024P069P004nsss(0) <='0';
          end if;
        if(cVar1S13S37N015N065N022P043(0)='1' AND  D( 9)='1' AND E(12)='1' )then
          cVar2S13S37P062P052nsss(0) <='1';
          else
          cVar2S13S37P062P052nsss(0) <='0';
          end if;
        if(cVar1S14S37N015N065N022P043(0)='1' AND  D( 9)='1' AND E(12)='0' AND E(18)='0' )then
          cVar2S14S37P062N052P061nsss(0) <='1';
          else
          cVar2S14S37P062N052P061nsss(0) <='0';
          end if;
        if(cVar1S15S37N015N065N022P043(0)='1' AND  D( 9)='0' AND D(17)='1' AND A(24)='1' )then
          cVar2S15S37N062P063P010nsss(0) <='1';
          else
          cVar2S15S37N062P063P010nsss(0) <='0';
          end if;
        if(cVar1S16S37N015N065N022P043(0)='1' AND  E(22)='1' AND A(17)='1' )then
          cVar2S16S37P045P005nsss(0) <='1';
          else
          cVar2S16S37P045P005nsss(0) <='0';
          end if;
        if(cVar1S17S37N015N065N022P043(0)='1' AND  E(22)='1' AND A(17)='0' AND A(22)='0' )then
          cVar2S17S37P045N005P014nsss(0) <='1';
          else
          cVar2S17S37P045N005P014nsss(0) <='0';
          end if;
        if(cVar1S18S37N015N065N022P043(0)='1' AND  E(22)='0' AND A(15)='1' )then
          cVar2S18S37N045P009nsss(0) <='1';
          else
          cVar2S18S37N045P009nsss(0) <='0';
          end if;
        if(cVar1S0S38P006P024P015P014(0)='1' AND  E(16)='0' AND E(10)='1' AND A(21)='0' )then
          cVar2S0S38P069P060P016nsss(0) <='1';
          else
          cVar2S0S38P069P060P016nsss(0) <='0';
          end if;
        if(cVar1S1S38P006P024P015P014(0)='1' AND  E(16)='0' AND E(10)='0' )then
          cVar2S1S38P069N060psss(0) <='1';
          else
          cVar2S1S38P069N060psss(0) <='0';
          end if;
        if(cVar1S2S38P006P024P015P014(0)='1' AND  E(16)='1' AND D(16)='1' AND B(22)='1' )then
          cVar2S2S38P069P067P032nsss(0) <='1';
          else
          cVar2S2S38P069P067P032nsss(0) <='0';
          end if;
        if(cVar1S3S38P006P024P015N014(0)='1' AND  D(16)='1' AND B(11)='0' )then
          cVar2S3S38P067P035nsss(0) <='1';
          else
          cVar2S3S38P067P035nsss(0) <='0';
          end if;
        if(cVar1S4S38P006P024P015N014(0)='1' AND  D(16)='1' AND B(11)='1' AND D(17)='1' )then
          cVar2S4S38P067P035P063nsss(0) <='1';
          else
          cVar2S4S38P067P035P063nsss(0) <='0';
          end if;
        if(cVar1S5S38P006P024P015N014(0)='1' AND  D(16)='0' AND B(22)='0' )then
          cVar2S5S38N067P032nsss(0) <='1';
          else
          cVar2S5S38N067P032nsss(0) <='0';
          end if;
        if(cVar1S6S38P006P024P015N014(0)='1' AND  D(16)='0' AND B(22)='1' AND A(23)='1' )then
          cVar2S6S38N067P032P012nsss(0) <='1';
          else
          cVar2S6S38N067P032P012nsss(0) <='0';
          end if;
        if(cVar1S7S38P006P024P015P053(0)='1' AND  A(29)='0' AND B(21)='0' )then
          cVar2S7S38P000P034nsss(0) <='1';
          else
          cVar2S7S38P000P034nsss(0) <='0';
          end if;
        if(cVar1S8S38P006P024P015N053(0)='1' AND  D(20)='0' AND D( 8)='1' )then
          cVar2S8S38P051P066nsss(0) <='1';
          else
          cVar2S8S38P051P066nsss(0) <='0';
          end if;
        if(cVar1S9S38P006P024P015N053(0)='1' AND  D(20)='1' AND A(22)='0' AND E(21)='1' )then
          cVar2S9S38P051P014P049nsss(0) <='1';
          else
          cVar2S9S38P051P014P049nsss(0) <='0';
          end if;
        if(cVar1S11S38P006P024P014N047(0)='1' AND  E(21)='0' AND A(29)='1' )then
          cVar2S11S38P049P000nsss(0) <='1';
          else
          cVar2S11S38P049P000nsss(0) <='0';
          end if;
        if(cVar1S12S38P006P024P014N047(0)='1' AND  E(21)='0' AND A(29)='0' AND A(11)='1' )then
          cVar2S12S38P049N000P017nsss(0) <='1';
          else
          cVar2S12S38P049N000P017nsss(0) <='0';
          end if;
        if(cVar1S13S38P006P024P014P067(0)='1' AND  B(25)='0' AND A(12)='0' AND D( 8)='0' )then
          cVar2S13S38P026P015P066nsss(0) <='1';
          else
          cVar2S13S38P026P015P066nsss(0) <='0';
          end if;
        if(cVar1S14S38P006P034P024P051(0)='1' AND  A(14)='0' AND A(13)='0' )then
          cVar2S14S38P011P013nsss(0) <='1';
          else
          cVar2S14S38P011P013nsss(0) <='0';
          end if;
        if(cVar1S15S38P006P034N024P065(0)='1' AND  A(17)='0' AND A(29)='0' AND D(16)='0' )then
          cVar2S15S38P005P000P067nsss(0) <='1';
          else
          cVar2S15S38P005P000P067nsss(0) <='0';
          end if;
        if(cVar1S16S38P006P034N024P065(0)='1' AND  A(17)='1' AND A(24)='1' )then
          cVar2S16S38P005P010nsss(0) <='1';
          else
          cVar2S16S38P005P010nsss(0) <='0';
          end if;
        if(cVar1S17S38P006P034N024P065(0)='1' AND  A(11)='0' AND A(24)='0' AND D(17)='0' )then
          cVar2S17S38P017P010P063nsss(0) <='1';
          else
          cVar2S17S38P017P010P063nsss(0) <='0';
          end if;
        if(cVar1S18S38P006P034P036P011(0)='1' AND  E( 8)='0' AND E(17)='1' )then
          cVar2S18S38P068P065nsss(0) <='1';
          else
          cVar2S18S38P068P065nsss(0) <='0';
          end if;
        if(cVar1S0S39P006P067P024P043(0)='1' AND  E(17)='1' AND E( 8)='0' AND D( 9)='0' )then
          cVar2S0S39P065P068P062nsss(0) <='1';
          else
          cVar2S0S39P065P068P062nsss(0) <='0';
          end if;
        if(cVar1S1S39P006P067P024P043(0)='1' AND  E(17)='1' AND E( 8)='1' AND A(23)='1' )then
          cVar2S1S39P065P068P012nsss(0) <='1';
          else
          cVar2S1S39P065P068P012nsss(0) <='0';
          end if;
        if(cVar1S2S39P006P067P024P043(0)='1' AND  E(17)='0' AND D(17)='0' )then
          cVar2S2S39N065P063nsss(0) <='1';
          else
          cVar2S2S39N065P063nsss(0) <='0';
          end if;
        if(cVar1S3S39P006P067P024P043(0)='1' AND  E(17)='0' AND D(17)='1' AND E( 9)='1' )then
          cVar2S3S39N065P063P064nsss(0) <='1';
          else
          cVar2S3S39N065P063P064nsss(0) <='0';
          end if;
        if(cVar1S4S39P006P067P024P043(0)='1' AND  E(22)='1' )then
          cVar2S4S39P045nsss(0) <='1';
          else
          cVar2S4S39P045nsss(0) <='0';
          end if;
        if(cVar1S5S39P006P067P024P014(0)='1' AND  B(11)='0' AND A(25)='0' AND A(12)='0' )then
          cVar2S5S39P035P008P015nsss(0) <='1';
          else
          cVar2S5S39P035P008P015nsss(0) <='0';
          end if;
        if(cVar1S6S39P006N067P015P045(0)='1' AND  B(27)='0' AND E( 8)='0' AND B(13)='0' )then
          cVar2S6S39P022P068P031nsss(0) <='1';
          else
          cVar2S6S39P022P068P031nsss(0) <='0';
          end if;
        if(cVar1S7S39P006N067P015P045(0)='1' AND  B(27)='0' AND E( 8)='1' AND E(18)='1' )then
          cVar2S7S39P022P068P061nsss(0) <='1';
          else
          cVar2S7S39P022P068P061nsss(0) <='0';
          end if;
        if(cVar1S8S39P006N067P015P045(0)='1' AND  B(27)='1' AND A(22)='0' AND A(20)='1' )then
          cVar2S8S39P022P014P018nsss(0) <='1';
          else
          cVar2S8S39P022P014P018nsss(0) <='0';
          end if;
        if(cVar1S9S39P006N067P015P045(0)='1' AND  B(20)='1' )then
          cVar2S9S39P036nsss(0) <='1';
          else
          cVar2S9S39P036nsss(0) <='0';
          end if;
        if(cVar1S10S39P006N067N015P014(0)='1' AND  E(16)='0' AND E(10)='1' AND B(20)='0' )then
          cVar2S10S39P069P060P036nsss(0) <='1';
          else
          cVar2S10S39P069P060P036nsss(0) <='0';
          end if;
        if(cVar1S11S39P006N067N015P014(0)='1' AND  E(16)='0' AND E(10)='0' )then
          cVar2S11S39P069N060psss(0) <='1';
          else
          cVar2S11S39P069N060psss(0) <='0';
          end if;
        if(cVar1S12S39P006N067N015N014(0)='1' AND  B(22)='0' AND B(10)='1' AND E(23)='1' )then
          cVar2S12S39P032P037P041nsss(0) <='1';
          else
          cVar2S12S39P032P037P041nsss(0) <='0';
          end if;
        if(cVar1S13S39P006N067N015N014(0)='1' AND  B(22)='1' AND A(23)='1' AND A(20)='0' )then
          cVar2S13S39P032P012P018nsss(0) <='1';
          else
          cVar2S13S39P032P012P018nsss(0) <='0';
          end if;
        if(cVar1S14S39P006P051P024P011(0)='1' AND  D(21)='1' )then
          cVar2S14S39P047nsss(0) <='1';
          else
          cVar2S14S39P047nsss(0) <='0';
          end if;
        if(cVar1S15S39P006P051P024P011(0)='1' AND  D(21)='0' AND A(13)='0' AND A(12)='0' )then
          cVar2S15S39N047P013P015nsss(0) <='1';
          else
          cVar2S15S39N047P013P015nsss(0) <='0';
          end if;
        if(cVar1S16S39P006P051N024P065(0)='1' AND  B(18)='1' )then
          cVar2S16S39P021nsss(0) <='1';
          else
          cVar2S16S39P021nsss(0) <='0';
          end if;
        if(cVar1S17S39P006P051N024P065(0)='1' AND  A(22)='0' AND A(13)='0' AND A(20)='0' )then
          cVar2S17S39P014P013P018nsss(0) <='1';
          else
          cVar2S17S39P014P013P018nsss(0) <='0';
          end if;
        if(cVar1S18S39P006P051P067P014(0)='1' AND  E(20)='0' )then
          cVar2S18S39P053nsss(0) <='1';
          else
          cVar2S18S39P053nsss(0) <='0';
          end if;
        if(cVar1S0S40P014P032P030P012(0)='1' AND  E(11)='1' )then
          cVar2S0S40P056nsss(0) <='1';
          else
          cVar2S0S40P056nsss(0) <='0';
          end if;
        if(cVar1S1S40P014P032P030P012(0)='1' AND  E(11)='0' AND A(20)='0' )then
          cVar2S1S40N056P018nsss(0) <='1';
          else
          cVar2S1S40N056P018nsss(0) <='0';
          end if;
        if(cVar1S2S40P014P032P030P012(0)='1' AND  E(11)='0' AND A(20)='1' AND A(12)='1' )then
          cVar2S2S40N056P018P015nsss(0) <='1';
          else
          cVar2S2S40N056P018P015nsss(0) <='0';
          end if;
        if(cVar1S3S40P014P032P030N012(0)='1' AND  A(24)='1' )then
          cVar2S3S40P010nsss(0) <='1';
          else
          cVar2S3S40P010nsss(0) <='0';
          end if;
        if(cVar1S4S40P014P032P030N012(0)='1' AND  A(24)='0' AND E(19)='1' )then
          cVar2S4S40N010P057nsss(0) <='1';
          else
          cVar2S4S40N010P057nsss(0) <='0';
          end if;
        if(cVar1S5S40P014P032P030N012(0)='1' AND  A(24)='0' AND E(19)='0' AND A(21)='1' )then
          cVar2S5S40N010N057P016nsss(0) <='1';
          else
          cVar2S5S40N010N057P016nsss(0) <='0';
          end if;
        if(cVar1S6S40P014P032N030P057(0)='1' AND  D(19)='0' AND B(15)='1' AND A(15)='1' )then
          cVar2S6S40P055P027P009nsss(0) <='1';
          else
          cVar2S6S40P055P027P009nsss(0) <='0';
          end if;
        if(cVar1S7S40P014P032N030P057(0)='1' AND  D(19)='0' AND B(15)='0' )then
          cVar2S7S40P055N027psss(0) <='1';
          else
          cVar2S7S40P055N027psss(0) <='0';
          end if;
        if(cVar1S8S40P014P032N030P057(0)='1' AND  D(19)='1' AND A(13)='0' AND A(21)='1' )then
          cVar2S8S40P055P013P016nsss(0) <='1';
          else
          cVar2S8S40P055P013P016nsss(0) <='0';
          end if;
        if(cVar1S9S40P014P032N030P057(0)='1' AND  B(13)='1' AND A(13)='1' )then
          cVar2S9S40P031P013nsss(0) <='1';
          else
          cVar2S9S40P031P013nsss(0) <='0';
          end if;
        if(cVar1S10S40P014P032N030P057(0)='1' AND  B(13)='0' AND A(29)='0' AND A(24)='1' )then
          cVar2S10S40N031P000P010nsss(0) <='1';
          else
          cVar2S10S40N031P000P010nsss(0) <='0';
          end if;
        if(cVar1S11S40P014P032P010P012(0)='1' AND  B(20)='0' AND B(10)='1' )then
          cVar2S11S40P036P037nsss(0) <='1';
          else
          cVar2S11S40P036P037nsss(0) <='0';
          end if;
        if(cVar1S12S40P014P032P010P012(0)='1' AND  B(20)='0' AND B(10)='0' AND E(18)='0' )then
          cVar2S12S40P036N037P061nsss(0) <='1';
          else
          cVar2S12S40P036N037P061nsss(0) <='0';
          end if;
        if(cVar1S13S40P014P032P010N012(0)='1' AND  A(20)='1' AND A(13)='1' )then
          cVar2S13S40P018P013nsss(0) <='1';
          else
          cVar2S13S40P018P013nsss(0) <='0';
          end if;
        if(cVar1S14S40P014P032P010N012(0)='1' AND  A(20)='1' AND A(13)='0' AND A(10)='0' )then
          cVar2S14S40P018N013P019nsss(0) <='1';
          else
          cVar2S14S40P018N013P019nsss(0) <='0';
          end if;
        if(cVar1S15S40P014P032P010P017(0)='1' AND  A(13)='1' )then
          cVar2S15S40P013nsss(0) <='1';
          else
          cVar2S15S40P013nsss(0) <='0';
          end if;
        if(cVar1S16S40P014P024P044P032(0)='1' AND  A(25)='0' AND E(10)='1' )then
          cVar2S16S40P008P060nsss(0) <='1';
          else
          cVar2S16S40P008P060nsss(0) <='0';
          end if;
        if(cVar1S17S40P014P024P044P032(0)='1' AND  A(25)='0' AND E(10)='0' AND B(21)='0' )then
          cVar2S17S40P008N060P034nsss(0) <='1';
          else
          cVar2S17S40P008N060P034nsss(0) <='0';
          end if;
        if(cVar1S18S40P014P024P044N032(0)='1' AND  E(16)='0' AND B(11)='1' AND A(23)='1' )then
          cVar2S18S40P069P035P012nsss(0) <='1';
          else
          cVar2S18S40P069P035P012nsss(0) <='0';
          end if;
        if(cVar1S19S40P014P024P044N032(0)='1' AND  E(16)='1' AND B(10)='1' AND D(16)='1' )then
          cVar2S19S40P069P037P067nsss(0) <='1';
          else
          cVar2S19S40P069P037P067nsss(0) <='0';
          end if;
        if(cVar1S20S40P014P024P044N032(0)='1' AND  E(16)='1' AND B(10)='0' AND B(11)='1' )then
          cVar2S20S40P069N037P035nsss(0) <='1';
          else
          cVar2S20S40P069N037P035nsss(0) <='0';
          end if;
        if(cVar1S21S40P014P024P044P062(0)='1' AND  A(11)='0' AND A(20)='1' )then
          cVar2S21S40P017P018nsss(0) <='1';
          else
          cVar2S21S40P017P018nsss(0) <='0';
          end if;
        if(cVar1S22S40P014P024P054P036(0)='1' AND  A(18)='0' AND D(22)='1' )then
          cVar2S22S40P003P043nsss(0) <='1';
          else
          cVar2S22S40P003P043nsss(0) <='0';
          end if;
        if(cVar1S1S41P035P015P027N050(0)='1' AND  A(22)='0' AND E(13)='1' )then
          cVar2S1S41P014P048nsss(0) <='1';
          else
          cVar2S1S41P014P048nsss(0) <='0';
          end if;
        if(cVar1S2S41P035P015N027P022(0)='1' AND  D(22)='1' )then
          cVar2S2S41P043nsss(0) <='1';
          else
          cVar2S2S41P043nsss(0) <='0';
          end if;
        if(cVar1S3S41P035P015N027P022(0)='1' AND  D(22)='0' AND A(11)='0' AND A(24)='0' )then
          cVar2S3S41N043P017P010nsss(0) <='1';
          else
          cVar2S3S41N043P017P010nsss(0) <='0';
          end if;
        if(cVar1S4S41P035P015N027N022(0)='1' AND  D(22)='0' AND E(11)='1' AND A(27)='0' )then
          cVar2S4S41P043P056P004nsss(0) <='1';
          else
          cVar2S4S41P043P056P004nsss(0) <='0';
          end if;
        if(cVar1S5S41P035P015N027N022(0)='1' AND  D(22)='0' AND E(11)='0' AND D(21)='1' )then
          cVar2S5S41P043N056P047nsss(0) <='1';
          else
          cVar2S5S41P043N056P047nsss(0) <='0';
          end if;
        if(cVar1S6S41P035P015N027N022(0)='1' AND  D(22)='1' AND A(17)='1' )then
          cVar2S6S41P043P005nsss(0) <='1';
          else
          cVar2S6S41P043P005nsss(0) <='0';
          end if;
        if(cVar1S7S41P035P015N027N022(0)='1' AND  D(22)='1' AND A(17)='0' AND B(26)='1' )then
          cVar2S7S41P043N005P024nsss(0) <='1';
          else
          cVar2S7S41P043N005P024nsss(0) <='0';
          end if;
        if(cVar1S8S41P035P015P026P061(0)='1' AND  A(27)='0' AND A(23)='0' )then
          cVar2S8S41P004P012nsss(0) <='1';
          else
          cVar2S8S41P004P012nsss(0) <='0';
          end if;
        if(cVar1S9S41P035P015P026P061(0)='1' AND  A(27)='0' AND A(23)='1' AND B(10)='1' )then
          cVar2S9S41P004P012P037nsss(0) <='1';
          else
          cVar2S9S41P004P012P037nsss(0) <='0';
          end if;
        if(cVar1S10S41P035P015N026P062(0)='1' AND  D(18)='1' AND E(11)='1' )then
          cVar2S10S41P059P056nsss(0) <='1';
          else
          cVar2S10S41P059P056nsss(0) <='0';
          end if;
        if(cVar1S11S41P035P015N026P062(0)='1' AND  D(18)='1' AND E(11)='0' AND A(27)='0' )then
          cVar2S11S41P059N056P004nsss(0) <='1';
          else
          cVar2S11S41P059N056P004nsss(0) <='0';
          end if;
        if(cVar1S12S41P035P015N026P062(0)='1' AND  D(18)='0' AND A(23)='1' AND A(13)='0' )then
          cVar2S12S41N059P012P013nsss(0) <='1';
          else
          cVar2S12S41N059P012P013nsss(0) <='0';
          end if;
        if(cVar1S13S41P035P015N026P062(0)='1' AND  D(18)='0' AND A(23)='0' AND A(18)='1' )then
          cVar2S13S41N059N012P003nsss(0) <='1';
          else
          cVar2S13S41N059N012P003nsss(0) <='0';
          end if;
        if(cVar1S14S41P035P015N026P062(0)='1' AND  A(15)='0' AND A(25)='1' AND A(21)='0' )then
          cVar2S14S41P009P008P016nsss(0) <='1';
          else
          cVar2S14S41P009P008P016nsss(0) <='0';
          end if;
        if(cVar1S15S41P035P045P006P063(0)='1' AND  A(23)='1' AND D(16)='0' )then
          cVar2S15S41P012P067nsss(0) <='1';
          else
          cVar2S15S41P012P067nsss(0) <='0';
          end if;
        if(cVar1S16S41P035P045P006P063(0)='1' AND  A(23)='0' AND A(15)='0' AND A(14)='0' )then
          cVar2S16S41N012P009P011nsss(0) <='1';
          else
          cVar2S16S41N012P009P011nsss(0) <='0';
          end if;
        if(cVar1S17S41P035P045P006N063(0)='1' AND  B(21)='0' AND B(27)='0' AND D(18)='1' )then
          cVar2S17S41P034P022P059nsss(0) <='1';
          else
          cVar2S17S41P034P022P059nsss(0) <='0';
          end if;
        if(cVar1S18S41P035P045P006N063(0)='1' AND  B(21)='1' AND B(10)='1' AND A(20)='1' )then
          cVar2S18S41P034P037P018nsss(0) <='1';
          else
          cVar2S18S41P034P037P018nsss(0) <='0';
          end if;
        if(cVar1S19S41P035P045P006P034(0)='1' AND  E(17)='0' AND A(23)='1' AND A(12)='0' )then
          cVar2S19S41P065P012P015nsss(0) <='1';
          else
          cVar2S19S41P065P012P015nsss(0) <='0';
          end if;
        if(cVar1S0S42P015P035P001P002(0)='1' AND  B(15)='1' AND D(12)='1' )then
          cVar2S0S42P027P050nsss(0) <='1';
          else
          cVar2S0S42P027P050nsss(0) <='0';
          end if;
        if(cVar1S1S42P015P035P001P002(0)='1' AND  B(15)='1' AND D(12)='0' AND E(21)='1' )then
          cVar2S1S42P027N050P049nsss(0) <='1';
          else
          cVar2S1S42P027N050P049nsss(0) <='0';
          end if;
        if(cVar1S2S42P015P035P001P002(0)='1' AND  B(15)='0' AND E(21)='0' AND A(16)='0' )then
          cVar2S2S42N027P049P007nsss(0) <='1';
          else
          cVar2S2S42N027P049P007nsss(0) <='0';
          end if;
        if(cVar1S3S42P015P035P001P002(0)='1' AND  B(15)='0' AND E(21)='1' AND D(21)='1' )then
          cVar2S3S42N027P049P047nsss(0) <='1';
          else
          cVar2S3S42N027P049P047nsss(0) <='0';
          end if;
        if(cVar1S4S42P015P035P001P002(0)='1' AND  E(15)='1' )then
          cVar2S4S42P040nsss(0) <='1';
          else
          cVar2S4S42P040nsss(0) <='0';
          end if;
        if(cVar1S5S42P015P035P001P002(0)='1' AND  E(15)='0' AND A(24)='0' AND A(16)='1' )then
          cVar2S5S42N040P010P007nsss(0) <='1';
          else
          cVar2S5S42N040P010P007nsss(0) <='0';
          end if;
        if(cVar1S6S42P015P035P001P013(0)='1' AND  B(12)='0' AND A(16)='0' AND A(18)='1' )then
          cVar2S6S42P033P007P003nsss(0) <='1';
          else
          cVar2S6S42P033P007P003nsss(0) <='0';
          end if;
        if(cVar1S7S42P015P035P020P045(0)='1' AND  D(16)='0' AND D(10)='1' AND B(10)='0' )then
          cVar2S7S42P067P058P037nsss(0) <='1';
          else
          cVar2S7S42P067P058P037nsss(0) <='0';
          end if;
        if(cVar1S8S42P015P035P020P045(0)='1' AND  D(16)='1' AND D( 8)='0' AND E(16)='1' )then
          cVar2S8S42P067P066P069nsss(0) <='1';
          else
          cVar2S8S42P067P066P069nsss(0) <='0';
          end if;
        if(cVar1S9S42P015P035P020P045(0)='1' AND  D(16)='1' AND D( 8)='1' AND A(25)='1' )then
          cVar2S9S42P067P066P008nsss(0) <='1';
          else
          cVar2S9S42P067P066P008nsss(0) <='0';
          end if;
        if(cVar1S10S42P015P009P034P055(0)='1' AND  D( 8)='0' AND B(11)='1' )then
          cVar2S10S42P066P035nsss(0) <='1';
          else
          cVar2S10S42P066P035nsss(0) <='0';
          end if;
        if(cVar1S11S42P015P009P034P055(0)='1' AND  D( 8)='0' AND B(11)='0' AND A(25)='0' )then
          cVar2S11S42P066N035P008nsss(0) <='1';
          else
          cVar2S11S42P066N035P008nsss(0) <='0';
          end if;
        if(cVar1S12S42P015P009P034P055(0)='1' AND  D( 8)='1' AND B(10)='1' )then
          cVar2S12S42P066P037nsss(0) <='1';
          else
          cVar2S12S42P066P037nsss(0) <='0';
          end if;
        if(cVar1S13S42P015P009P034N055(0)='1' AND  E(17)='0' AND B(20)='0' AND D( 8)='1' )then
          cVar2S13S42P065P036P066nsss(0) <='1';
          else
          cVar2S13S42P065P036P066nsss(0) <='0';
          end if;
        if(cVar1S14S42P015P009P034N055(0)='1' AND  E(17)='1' AND A(20)='1' AND E( 8)='1' )then
          cVar2S14S42P065P018P068nsss(0) <='1';
          else
          cVar2S14S42P065P018P068nsss(0) <='0';
          end if;
        if(cVar1S15S42P015P009P034N055(0)='1' AND  E(17)='1' AND A(20)='0' AND B(11)='1' )then
          cVar2S15S42P065N018P035nsss(0) <='1';
          else
          cVar2S15S42P065N018P035nsss(0) <='0';
          end if;
        if(cVar1S16S42P015P009P034P063(0)='1' AND  A(13)='0' AND A(10)='0' AND A(23)='0' )then
          cVar2S16S42P013P019P012nsss(0) <='1';
          else
          cVar2S16S42P013P019P012nsss(0) <='0';
          end if;
        if(cVar1S17S42P015P009P034P063(0)='1' AND  A(13)='0' AND A(10)='1' AND A(20)='0' )then
          cVar2S17S42P013P019P018nsss(0) <='1';
          else
          cVar2S17S42P013P019P018nsss(0) <='0';
          end if;
        if(cVar1S18S42P015P009P034P063(0)='1' AND  A(13)='1' AND A(21)='1' AND A(22)='0' )then
          cVar2S18S42P013P016P014nsss(0) <='1';
          else
          cVar2S18S42P013P016P014nsss(0) <='0';
          end if;
        if(cVar1S19S42P015P009P034N063(0)='1' AND  E(17)='0' AND A(20)='1' AND A(24)='0' )then
          cVar2S19S42P065P018P010nsss(0) <='1';
          else
          cVar2S19S42P065P018P010nsss(0) <='0';
          end if;
        if(cVar1S20S42P015P009P041P004(0)='1' AND  B(15)='1' )then
          cVar2S20S42P027nsss(0) <='1';
          else
          cVar2S20S42P027nsss(0) <='0';
          end if;
        if(cVar1S0S43P015P034P022P016(0)='1' AND  A(15)='0' AND B(22)='1' AND B(12)='0' )then
          cVar2S0S43P009P032P033nsss(0) <='1';
          else
          cVar2S0S43P009P032P033nsss(0) <='0';
          end if;
        if(cVar1S1S43P015P034P022P016(0)='1' AND  A(15)='0' AND B(22)='0' )then
          cVar2S1S43P009N032psss(0) <='1';
          else
          cVar2S1S43P009N032psss(0) <='0';
          end if;
        if(cVar1S2S43P015P034P022P016(0)='1' AND  A(15)='1' AND A(27)='0' AND D(16)='1' )then
          cVar2S2S43P009P004P067nsss(0) <='1';
          else
          cVar2S2S43P009P004P067nsss(0) <='0';
          end if;
        if(cVar1S3S43P015P034P022P016(0)='1' AND  A(25)='0' AND A(28)='0' AND D(12)='0' )then
          cVar2S3S43P008P002P050nsss(0) <='1';
          else
          cVar2S3S43P008P002P050nsss(0) <='0';
          end if;
        if(cVar1S4S43P015P034P022P016(0)='1' AND  A(25)='1' AND A(20)='0' AND D(18)='0' )then
          cVar2S4S43P008P018P059nsss(0) <='1';
          else
          cVar2S4S43P008P018P059nsss(0) <='0';
          end if;
        if(cVar1S5S43P015P034P022P009(0)='1' AND  A(21)='0' AND A(10)='1' )then
          cVar2S5S43P016P019nsss(0) <='1';
          else
          cVar2S5S43P016P019nsss(0) <='0';
          end if;
        if(cVar1S6S43P015P034P043P044(0)='1' AND  E(19)='0' AND D(17)='1' AND A(26)='0' )then
          cVar2S6S43P057P063P006nsss(0) <='1';
          else
          cVar2S6S43P057P063P006nsss(0) <='0';
          end if;
        if(cVar1S8S43N015P027N048P005(0)='1' AND  E(21)='1' )then
          cVar2S8S43P049nsss(0) <='1';
          else
          cVar2S8S43P049nsss(0) <='0';
          end if;
        if(cVar1S9S43N015P027N048P005(0)='1' AND  E(21)='0' AND B(11)='0' AND A(18)='1' )then
          cVar2S9S43N049P035P003nsss(0) <='1';
          else
          cVar2S9S43N049P035P003nsss(0) <='0';
          end if;
        if(cVar1S10S43N015N027P030P012(0)='1' AND  A(20)='0' AND A(14)='0' AND A(24)='0' )then
          cVar2S10S43P018P011P010nsss(0) <='1';
          else
          cVar2S10S43P018P011P010nsss(0) <='0';
          end if;
        if(cVar1S11S43N015N027P030N012(0)='1' AND  A(24)='1' )then
          cVar2S11S43P010nsss(0) <='1';
          else
          cVar2S11S43P010nsss(0) <='0';
          end if;
        if(cVar1S12S43N015N027P030N012(0)='1' AND  A(24)='0' AND E(19)='1' )then
          cVar2S12S43N010P057nsss(0) <='1';
          else
          cVar2S12S43N010P057nsss(0) <='0';
          end if;
        if(cVar1S13S43N015N027P030N012(0)='1' AND  A(24)='0' AND E(19)='0' AND A(21)='1' )then
          cVar2S13S43N010N057P016nsss(0) <='1';
          else
          cVar2S13S43N010N057P016nsss(0) <='0';
          end if;
        if(cVar1S14S43N015N027N030P040(0)='1' AND  B(18)='1' )then
          cVar2S14S43P021nsss(0) <='1';
          else
          cVar2S14S43P021nsss(0) <='0';
          end if;
        if(cVar1S15S43N015N027N030P040(0)='1' AND  B(18)='0' AND B(28)='1' )then
          cVar2S15S43N021P020nsss(0) <='1';
          else
          cVar2S15S43N021P020nsss(0) <='0';
          end if;
        if(cVar1S16S43N015N027N030P040(0)='1' AND  B(18)='0' AND B(28)='0' AND A(20)='1' )then
          cVar2S16S43N021N020P018nsss(0) <='1';
          else
          cVar2S16S43N021N020P018nsss(0) <='0';
          end if;
        if(cVar1S17S43N015N027N030N040(0)='1' AND  D(15)='0' AND A(28)='0' AND B(14)='1' )then
          cVar2S17S43P038P002P029nsss(0) <='1';
          else
          cVar2S17S43P038P002P029nsss(0) <='0';
          end if;
        if(cVar1S1S44P015P027P000N048(0)='1' AND  A(17)='0' AND B(11)='0' )then
          cVar2S1S44P005P035nsss(0) <='1';
          else
          cVar2S1S44P005P035nsss(0) <='0';
          end if;
        if(cVar1S2S44P015N027P018P068(0)='1' AND  A(22)='1' AND D( 8)='0' )then
          cVar2S2S44P014P066nsss(0) <='1';
          else
          cVar2S2S44P014P066nsss(0) <='0';
          end if;
        if(cVar1S3S44P015N027P018P068(0)='1' AND  A(22)='0' AND B(22)='0' )then
          cVar2S3S44N014P032nsss(0) <='1';
          else
          cVar2S3S44N014P032nsss(0) <='0';
          end if;
        if(cVar1S4S44P015N027P018P068(0)='1' AND  A(22)='0' AND B(22)='1' AND A(23)='1' )then
          cVar2S4S44N014P032P012nsss(0) <='1';
          else
          cVar2S4S44N014P032P012nsss(0) <='0';
          end if;
        if(cVar1S5S44P015N027P018P068(0)='1' AND  D(16)='0' AND B(22)='1' AND B(10)='0' )then
          cVar2S5S44P067P032P037nsss(0) <='1';
          else
          cVar2S5S44P067P032P037nsss(0) <='0';
          end if;
        if(cVar1S6S44P015N027P018P068(0)='1' AND  D(16)='0' AND B(22)='0' AND D(20)='1' )then
          cVar2S6S44P067N032P051nsss(0) <='1';
          else
          cVar2S6S44P067N032P051nsss(0) <='0';
          end if;
        if(cVar1S7S44P015N027P018P068(0)='1' AND  D(16)='1' AND A(23)='1' AND A(10)='1' )then
          cVar2S7S44P067P012P019nsss(0) <='1';
          else
          cVar2S7S44P067P012P019nsss(0) <='0';
          end if;
        if(cVar1S8S44P015N027P018P013(0)='1' AND  B(13)='1' )then
          cVar2S8S44P031nsss(0) <='1';
          else
          cVar2S8S44P031nsss(0) <='0';
          end if;
        if(cVar1S9S44P015N027P018P013(0)='1' AND  B(13)='0' AND E(18)='1' AND D(17)='0' )then
          cVar2S9S44N031P061P063nsss(0) <='1';
          else
          cVar2S9S44N031P061P063nsss(0) <='0';
          end if;
        if(cVar1S10S44P015N027P018P013(0)='1' AND  B(13)='0' AND E(18)='0' AND A(14)='0' )then
          cVar2S10S44N031N061P011nsss(0) <='1';
          else
          cVar2S10S44N031N061P011nsss(0) <='0';
          end if;
        if(cVar1S11S44P015N027P018N013(0)='1' AND  A(29)='1' AND B(20)='0' AND E(16)='0' )then
          cVar2S11S44P000P036P069nsss(0) <='1';
          else
          cVar2S11S44P000P036P069nsss(0) <='0';
          end if;
        if(cVar1S12S44P015N027P018N013(0)='1' AND  A(29)='0' AND E( 8)='1' AND D(19)='0' )then
          cVar2S12S44N000P068P055nsss(0) <='1';
          else
          cVar2S12S44N000P068P055nsss(0) <='0';
          end if;
        if(cVar1S13S44P015N027P018N013(0)='1' AND  A(29)='0' AND E( 8)='0' AND A(14)='1' )then
          cVar2S13S44N000N068P011nsss(0) <='1';
          else
          cVar2S13S44N000N068P011nsss(0) <='0';
          end if;
        if(cVar1S14S44P015P051P068P036(0)='1' AND  B(13)='0' AND E(17)='0' AND D(21)='0' )then
          cVar2S14S44P031P065P047nsss(0) <='1';
          else
          cVar2S14S44P031P065P047nsss(0) <='0';
          end if;
        if(cVar1S15S44P015P051P068P036(0)='1' AND  B(13)='0' AND E(17)='1' AND A(10)='0' )then
          cVar2S15S44P031P065P019nsss(0) <='1';
          else
          cVar2S15S44P031P065P019nsss(0) <='0';
          end if;
        if(cVar1S16S44P015P051P068P036(0)='1' AND  B(13)='1' AND B(21)='1' )then
          cVar2S16S44P031P034nsss(0) <='1';
          else
          cVar2S16S44P031P034nsss(0) <='0';
          end if;
        if(cVar1S17S44P015P051P068P036(0)='1' AND  A(25)='0' AND A(27)='0' AND B(10)='1' )then
          cVar2S17S44P008P004P037nsss(0) <='1';
          else
          cVar2S17S44P008P004P037nsss(0) <='0';
          end if;
        if(cVar1S18S44P015P051P068P018(0)='1' AND  E(19)='0' AND A(29)='0' )then
          cVar2S18S44P057P000nsss(0) <='1';
          else
          cVar2S18S44P057P000nsss(0) <='0';
          end if;
        if(cVar1S19S44P015P051P068N018(0)='1' AND  D(17)='0' AND A(21)='1' AND A(15)='0' )then
          cVar2S19S44P063P016P009nsss(0) <='1';
          else
          cVar2S19S44P063P016P009nsss(0) <='0';
          end if;
        if(cVar1S20S44P015P051P068N018(0)='1' AND  D(17)='0' AND A(21)='0' AND A(22)='1' )then
          cVar2S20S44P063N016P014nsss(0) <='1';
          else
          cVar2S20S44P063N016P014nsss(0) <='0';
          end if;
        if(cVar1S21S44P015P051P053P000(0)='1' AND  A(26)='0' AND B(11)='0' )then
          cVar2S21S44P006P035nsss(0) <='1';
          else
          cVar2S21S44P006P035nsss(0) <='0';
          end if;
        if(cVar1S22S44P015P051N053P049(0)='1' AND  A(23)='0' )then
          cVar2S22S44P012nsss(0) <='1';
          else
          cVar2S22S44P012nsss(0) <='0';
          end if;
        if(cVar1S0S45P015P018P030P056(0)='1' AND  A(29)='1' AND A(21)='1' )then
          cVar2S0S45P000P016nsss(0) <='1';
          else
          cVar2S0S45P000P016nsss(0) <='0';
          end if;
        if(cVar1S1S45P015P018P030P056(0)='1' AND  A(29)='1' AND A(21)='0' AND D(16)='0' )then
          cVar2S1S45P000N016P067nsss(0) <='1';
          else
          cVar2S1S45P000N016P067nsss(0) <='0';
          end if;
        if(cVar1S2S45P015P018P030P056(0)='1' AND  A(29)='0' AND E(16)='0' AND B(22)='0' )then
          cVar2S2S45N000P069P032nsss(0) <='1';
          else
          cVar2S2S45N000P069P032nsss(0) <='0';
          end if;
        if(cVar1S3S45P015P018P030P056(0)='1' AND  A(29)='0' AND E(16)='1' AND D(16)='1' )then
          cVar2S3S45N000P069P067nsss(0) <='1';
          else
          cVar2S3S45N000P069P067nsss(0) <='0';
          end if;
        if(cVar1S4S45P015P018P030P056(0)='1' AND  E( 9)='1' )then
          cVar2S4S45P064nsss(0) <='1';
          else
          cVar2S4S45P064nsss(0) <='0';
          end if;
        if(cVar1S5S45P015P018P030P056(0)='1' AND  E( 9)='0' AND E(16)='1' AND A(13)='1' )then
          cVar2S5S45N064P069P013nsss(0) <='1';
          else
          cVar2S5S45N064P069P013nsss(0) <='0';
          end if;
        if(cVar1S7S45P015P018P030N069(0)='1' AND  E(19)='0' AND A(21)='1' AND A(22)='1' )then
          cVar2S7S45N057P016P014nsss(0) <='1';
          else
          cVar2S7S45N057P016P014nsss(0) <='0';
          end if;
        if(cVar1S8S45P015N018P019P017(0)='1' AND  B(21)='1' AND E( 9)='1' )then
          cVar2S8S45P034P064nsss(0) <='1';
          else
          cVar2S8S45P034P064nsss(0) <='0';
          end if;
        if(cVar1S9S45P015N018P019P017(0)='1' AND  B(21)='1' AND E( 9)='0' AND D( 8)='0' )then
          cVar2S9S45P034N064P066nsss(0) <='1';
          else
          cVar2S9S45P034N064P066nsss(0) <='0';
          end if;
        if(cVar1S10S45P015N018P019P017(0)='1' AND  B(21)='0' )then
          cVar2S10S45N034psss(0) <='1';
          else
          cVar2S10S45N034psss(0) <='0';
          end if;
        if(cVar1S11S45P015N018P019P017(0)='1' AND  E( 9)='0' AND B(14)='0' AND E(16)='1' )then
          cVar2S11S45P064P029P069nsss(0) <='1';
          else
          cVar2S11S45P064P029P069nsss(0) <='0';
          end if;
        if(cVar1S12S45P015N018P019P017(0)='1' AND  E( 9)='1' AND A(24)='1' )then
          cVar2S12S45P064P010nsss(0) <='1';
          else
          cVar2S12S45P064P010nsss(0) <='0';
          end if;
        if(cVar1S13S45P015N018N019P067(0)='1' AND  A(22)='1' AND A(11)='1' AND D( 8)='0' )then
          cVar2S13S45P014P017P066nsss(0) <='1';
          else
          cVar2S13S45P014P017P066nsss(0) <='0';
          end if;
        if(cVar1S14S45P015N018N019P067(0)='1' AND  A(22)='1' AND A(11)='0' AND D(21)='0' )then
          cVar2S14S45P014N017P047nsss(0) <='1';
          else
          cVar2S14S45P014N017P047nsss(0) <='0';
          end if;
        if(cVar1S15S45P015N018N019P067(0)='1' AND  A(22)='0' AND B(15)='1' )then
          cVar2S15S45N014P027nsss(0) <='1';
          else
          cVar2S15S45N014P027nsss(0) <='0';
          end if;
        if(cVar1S16S45P015N018N019P067(0)='1' AND  A(22)='0' AND B(15)='0' AND D( 8)='1' )then
          cVar2S16S45N014N027P066nsss(0) <='1';
          else
          cVar2S16S45N014N027P066nsss(0) <='0';
          end if;
        if(cVar1S17S45P015P051P068P022(0)='1' AND  B(16)='1' AND A(20)='0' )then
          cVar2S17S45P025P018nsss(0) <='1';
          else
          cVar2S17S45P025P018nsss(0) <='0';
          end if;
        if(cVar1S18S45P015P051P068P022(0)='1' AND  A(13)='0' AND A(10)='1' )then
          cVar2S18S45P013P019nsss(0) <='1';
          else
          cVar2S18S45P013P019nsss(0) <='0';
          end if;
        if(cVar1S19S45P015P051P068P018(0)='1' AND  E(19)='0' AND A(26)='0' )then
          cVar2S19S45P057P006nsss(0) <='1';
          else
          cVar2S19S45P057P006nsss(0) <='0';
          end if;
        if(cVar1S20S45P015P051P068N018(0)='1' AND  E(20)='0' AND D(17)='0' AND A(21)='1' )then
          cVar2S20S45P053P063P016nsss(0) <='1';
          else
          cVar2S20S45P053P063P016nsss(0) <='0';
          end if;
        if(cVar1S21S45P015P051P053P000(0)='1' AND  A(26)='0' AND A(23)='0' AND A(21)='0' )then
          cVar2S21S45P006P012P016nsss(0) <='1';
          else
          cVar2S21S45P006P012P016nsss(0) <='0';
          end if;
        if(cVar1S22S45P015P051N053P049(0)='1' AND  A(22)='0' )then
          cVar2S22S45P014nsss(0) <='1';
          else
          cVar2S22S45P014nsss(0) <='0';
          end if;
        if(cVar1S0S46P068P019P057P030(0)='1' AND  A(22)='0' )then
          cVar2S0S46P014nsss(0) <='1';
          else
          cVar2S0S46P014nsss(0) <='0';
          end if;
        if(cVar1S1S46P068P019P057N030(0)='1' AND  B(13)='1' AND A(13)='1' )then
          cVar2S1S46P031P013nsss(0) <='1';
          else
          cVar2S1S46P031P013nsss(0) <='0';
          end if;
        if(cVar1S2S46P068P019P057N030(0)='1' AND  B(13)='0' AND A(21)='1' AND A(22)='0' )then
          cVar2S2S46N031P016P014nsss(0) <='1';
          else
          cVar2S2S46N031P016P014nsss(0) <='0';
          end if;
        if(cVar1S3S46P068P019N057P005(0)='1' AND  B(17)='1' )then
          cVar2S3S46P023nsss(0) <='1';
          else
          cVar2S3S46P023nsss(0) <='0';
          end if;
        if(cVar1S4S46P068P019N057P005(0)='1' AND  B(17)='0' AND B(13)='0' )then
          cVar2S4S46N023P031nsss(0) <='1';
          else
          cVar2S4S46N023P031nsss(0) <='0';
          end if;
        if(cVar1S5S46P068P019N057N005(0)='1' AND  E(10)='1' AND D( 9)='1' )then
          cVar2S5S46P060P062nsss(0) <='1';
          else
          cVar2S5S46P060P062nsss(0) <='0';
          end if;
        if(cVar1S6S46P068P019N057N005(0)='1' AND  E(10)='1' AND D( 9)='0' AND A(23)='0' )then
          cVar2S6S46P060N062P012nsss(0) <='1';
          else
          cVar2S6S46P060N062P012nsss(0) <='0';
          end if;
        if(cVar1S7S46P068P019N057N005(0)='1' AND  E(10)='0' AND A(16)='1' AND D(18)='0' )then
          cVar2S7S46N060P007P059nsss(0) <='1';
          else
          cVar2S7S46N060P007P059nsss(0) <='0';
          end if;
        if(cVar1S8S46P068P019N057N005(0)='1' AND  E(10)='0' AND A(16)='0' AND B(17)='0' )then
          cVar2S8S46N060N007P023nsss(0) <='1';
          else
          cVar2S8S46N060N007P023nsss(0) <='0';
          end if;
        if(cVar1S9S46P068P019P006P043(0)='1' AND  E(21)='0' AND B(12)='0' AND A(19)='1' )then
          cVar2S9S46P049P033P001nsss(0) <='1';
          else
          cVar2S9S46P049P033P001nsss(0) <='0';
          end if;
        if(cVar1S10S46P068P019P006P043(0)='1' AND  E(21)='1' AND D(20)='0' AND E(16)='0' )then
          cVar2S10S46P049P051P069nsss(0) <='1';
          else
          cVar2S10S46P049P051P069nsss(0) <='0';
          end if;
        if(cVar1S11S46P068P019P006P043(0)='1' AND  A(22)='0' AND E(22)='1' )then
          cVar2S11S46P014P045nsss(0) <='1';
          else
          cVar2S11S46P014P045nsss(0) <='0';
          end if;
        if(cVar1S12S46P068P019P006P060(0)='1' AND  D(23)='0' AND A(24)='0' AND A(21)='0' )then
          cVar2S12S46P039P010P016nsss(0) <='1';
          else
          cVar2S12S46P039P010P016nsss(0) <='0';
          end if;
        if(cVar1S13S46P068P009P064P053(0)='1' AND  E(16)='0' AND B(21)='1' )then
          cVar2S13S46P069P034nsss(0) <='1';
          else
          cVar2S13S46P069P034nsss(0) <='0';
          end if;
        if(cVar1S14S46P068P009P064P053(0)='1' AND  E(16)='0' AND B(21)='0' AND D( 8)='1' )then
          cVar2S14S46P069N034P066nsss(0) <='1';
          else
          cVar2S14S46P069N034P066nsss(0) <='0';
          end if;
        if(cVar1S15S46P068P009P064P053(0)='1' AND  E(16)='1' AND B(20)='1' )then
          cVar2S15S46P069P036nsss(0) <='1';
          else
          cVar2S15S46P069P036nsss(0) <='0';
          end if;
        if(cVar1S16S46P068P009N064P056(0)='1' AND  B(13)='1' )then
          cVar2S16S46P031nsss(0) <='1';
          else
          cVar2S16S46P031nsss(0) <='0';
          end if;
        if(cVar1S17S46P068P009N064P056(0)='1' AND  B(13)='0' AND B(23)='1' )then
          cVar2S17S46N031P030nsss(0) <='1';
          else
          cVar2S17S46N031P030nsss(0) <='0';
          end if;
        if(cVar1S18S46P068P009N064N056(0)='1' AND  E(19)='0' AND A(25)='1' AND A(27)='0' )then
          cVar2S18S46P057P008P004nsss(0) <='1';
          else
          cVar2S18S46P057P008P004nsss(0) <='0';
          end if;
        if(cVar1S19S46P068P009N064N056(0)='1' AND  E(19)='1' AND E(16)='1' )then
          cVar2S19S46P057P069nsss(0) <='1';
          else
          cVar2S19S46P057P069nsss(0) <='0';
          end if;
        if(cVar1S20S46P068P009P002P066(0)='1' AND  B(10)='1' AND E(10)='0' AND D( 9)='1' )then
          cVar2S20S46P037P060P062nsss(0) <='1';
          else
          cVar2S20S46P037P060P062nsss(0) <='0';
          end if;
        if(cVar1S21S46P068P009P002P066(0)='1' AND  B(10)='0' AND E(16)='0' AND B(20)='1' )then
          cVar2S21S46N037P069P036nsss(0) <='1';
          else
          cVar2S21S46N037P069P036nsss(0) <='0';
          end if;
        if(cVar1S0S47P019P033P006P043(0)='1' AND  D(18)='1' AND A(29)='0' AND E(19)='0' )then
          cVar2S0S47P059P000P057nsss(0) <='1';
          else
          cVar2S0S47P059P000P057nsss(0) <='0';
          end if;
        if(cVar1S1S47P019P033P006P043(0)='1' AND  D(18)='0' AND E(18)='0' )then
          cVar2S1S47N059P061nsss(0) <='1';
          else
          cVar2S1S47N059P061nsss(0) <='0';
          end if;
        if(cVar1S2S47P019P033P006P043(0)='1' AND  E(22)='1' AND A(22)='0' )then
          cVar2S2S47P045P014nsss(0) <='1';
          else
          cVar2S2S47P045P014nsss(0) <='0';
          end if;
        if(cVar1S3S47P019P033P006P010(0)='1' AND  E(10)='0' AND B(26)='1' )then
          cVar2S3S47P060P024nsss(0) <='1';
          else
          cVar2S3S47P060P024nsss(0) <='0';
          end if;
        if(cVar1S4S47P019P033P006P010(0)='1' AND  E( 8)='1' AND A(13)='0' )then
          cVar2S4S47P068P013nsss(0) <='1';
          else
          cVar2S4S47P068P013nsss(0) <='0';
          end if;
        if(cVar1S5S47P019P033P016P065(0)='1' AND  D(18)='1' )then
          cVar2S5S47P059nsss(0) <='1';
          else
          cVar2S5S47P059nsss(0) <='0';
          end if;
        if(cVar1S6S47P019P033P016P065(0)='1' AND  D(18)='0' AND E(16)='0' AND D( 8)='1' )then
          cVar2S6S47N059P069P066nsss(0) <='1';
          else
          cVar2S6S47N059P069P066nsss(0) <='0';
          end if;
        if(cVar1S7S47P019P033P016P067(0)='1' AND  A(14)='0' )then
          cVar2S7S47P011nsss(0) <='1';
          else
          cVar2S7S47P011nsss(0) <='0';
          end if;
        if(cVar1S8S47P019P033P016N067(0)='1' AND  A(13)='1' AND A(22)='0' )then
          cVar2S8S47P013P014nsss(0) <='1';
          else
          cVar2S8S47P013P014nsss(0) <='0';
          end if;
        if(cVar1S9S47N019P057P041P000(0)='1' AND  A(24)='1' AND B(24)='1' )then
          cVar2S9S47P010P028nsss(0) <='1';
          else
          cVar2S9S47P010P028nsss(0) <='0';
          end if;
        if(cVar1S10S47N019P057P041P000(0)='1' AND  A(24)='1' AND B(24)='0' AND B(23)='1' )then
          cVar2S10S47P010N028P030nsss(0) <='1';
          else
          cVar2S10S47P010N028P030nsss(0) <='0';
          end if;
        if(cVar1S11S47N019P057P041P000(0)='1' AND  A(24)='0' AND B(20)='1' AND A(22)='0' )then
          cVar2S11S47N010P036P014nsss(0) <='1';
          else
          cVar2S11S47N010P036P014nsss(0) <='0';
          end if;
        if(cVar1S12S47N019P057P041P000(0)='1' AND  A(24)='0' AND B(20)='0' AND A(25)='0' )then
          cVar2S12S47N010N036P008nsss(0) <='1';
          else
          cVar2S12S47N010N036P008nsss(0) <='0';
          end if;
        if(cVar1S13S47N019N057P069P030(0)='1' AND  D(18)='0' AND E(18)='0' AND E(15)='1' )then
          cVar2S13S47P059P061P040nsss(0) <='1';
          else
          cVar2S13S47P059P061P040nsss(0) <='0';
          end if;
        if(cVar1S14S47N019N057P069P030(0)='1' AND  D(18)='0' AND E(18)='1' AND A(20)='1' )then
          cVar2S14S47P059P061P018nsss(0) <='1';
          else
          cVar2S14S47P059P061P018nsss(0) <='0';
          end if;
        if(cVar1S15S47N019N057P069P030(0)='1' AND  D(18)='1' AND B(12)='1' AND D(10)='0' )then
          cVar2S15S47P059P033P058nsss(0) <='1';
          else
          cVar2S15S47P059P033P058nsss(0) <='0';
          end if;
        if(cVar1S16S47N019N057P069P030(0)='1' AND  A(28)='1' )then
          cVar2S16S47P002nsss(0) <='1';
          else
          cVar2S16S47P002nsss(0) <='0';
          end if;
        if(cVar1S17S47N019N057P069P030(0)='1' AND  A(28)='0' AND D(11)='1' )then
          cVar2S17S47N002P054nsss(0) <='1';
          else
          cVar2S17S47N002P054nsss(0) <='0';
          end if;
        if(cVar1S18S47N019N057P069P030(0)='1' AND  A(28)='0' AND D(11)='0' AND A(16)='1' )then
          cVar2S18S47N002N054P007nsss(0) <='1';
          else
          cVar2S18S47N002N054P007nsss(0) <='0';
          end if;
        if(cVar1S19S47N019N057P069P029(0)='1' AND  D( 8)='0' )then
          cVar2S19S47P066nsss(0) <='1';
          else
          cVar2S19S47P066nsss(0) <='0';
          end if;
        if(cVar1S20S47N019N057P069N029(0)='1' AND  D(20)='0' AND E(18)='1' AND B(22)='1' )then
          cVar2S20S47P051P061P032nsss(0) <='1';
          else
          cVar2S20S47P051P061P032nsss(0) <='0';
          end if;
        if(cVar1S21S47N019N057P069N029(0)='1' AND  D(20)='1' AND E(20)='1' AND A(20)='1' )then
          cVar2S21S47P051P053P018nsss(0) <='1';
          else
          cVar2S21S47P051P053P018nsss(0) <='0';
          end if;
        if(cVar1S0S48P019P069P061P007(0)='1' AND  B(16)='1' )then
          cVar2S0S48P025nsss(0) <='1';
          else
          cVar2S0S48P025nsss(0) <='0';
          end if;
        if(cVar1S1S48P019P069P061P007(0)='1' AND  B(16)='0' AND A(15)='1' AND A(14)='0' )then
          cVar2S1S48N025P009P011nsss(0) <='1';
          else
          cVar2S1S48N025P009P011nsss(0) <='0';
          end if;
        if(cVar1S2S48P019P069P061P007(0)='1' AND  B(16)='0' AND A(15)='0' AND A(26)='0' )then
          cVar2S2S48N025N009P006nsss(0) <='1';
          else
          cVar2S2S48N025N009P006nsss(0) <='0';
          end if;
        if(cVar1S3S48P019P069P061N007(0)='1' AND  E(21)='0' AND D(21)='0' )then
          cVar2S3S48P049P047nsss(0) <='1';
          else
          cVar2S3S48P049P047nsss(0) <='0';
          end if;
        if(cVar1S4S48P019P069P061N007(0)='1' AND  E(21)='1' AND A(15)='1' )then
          cVar2S4S48P049P009nsss(0) <='1';
          else
          cVar2S4S48P049P009nsss(0) <='0';
          end if;
        if(cVar1S5S48P019P069P061N007(0)='1' AND  E(21)='1' AND A(15)='0' AND B(25)='1' )then
          cVar2S5S48P049N009P026nsss(0) <='1';
          else
          cVar2S5S48P049N009P026nsss(0) <='0';
          end if;
        if(cVar1S6S48P019P069P061P033(0)='1' AND  B(22)='0' )then
          cVar2S6S48P032nsss(0) <='1';
          else
          cVar2S6S48P032nsss(0) <='0';
          end if;
        if(cVar1S7S48P019P069P061N033(0)='1' AND  B(23)='1' )then
          cVar2S7S48P030nsss(0) <='1';
          else
          cVar2S7S48P030nsss(0) <='0';
          end if;
        if(cVar1S8S48P019P069P061N033(0)='1' AND  B(23)='0' AND B(13)='1' )then
          cVar2S8S48N030P031nsss(0) <='1';
          else
          cVar2S8S48N030P031nsss(0) <='0';
          end if;
        if(cVar1S9S48P019P069P045P043(0)='1' AND  B(14)='1' AND E( 8)='0' )then
          cVar2S9S48P029P068nsss(0) <='1';
          else
          cVar2S9S48P029P068nsss(0) <='0';
          end if;
        if(cVar1S10S48P019P069P045P043(0)='1' AND  B(14)='0' AND A(18)='0' AND B(22)='1' )then
          cVar2S10S48N029P003P032nsss(0) <='1';
          else
          cVar2S10S48N029P003P032nsss(0) <='0';
          end if;
        if(cVar1S11S48P019P059P041P003(0)='1' AND  E(20)='0' AND B(28)='0' )then
          cVar2S11S48P053P020nsss(0) <='1';
          else
          cVar2S11S48P053P020nsss(0) <='0';
          end if;
        if(cVar1S12S48P019N059P061P033(0)='1' AND  A(18)='1' AND E( 9)='0' AND E(19)='0' )then
          cVar2S12S48P003P064P057nsss(0) <='1';
          else
          cVar2S12S48P003P064P057nsss(0) <='0';
          end if;
        if(cVar1S13S48P019N059P061P033(0)='1' AND  A(18)='0' AND B(25)='1' AND A(25)='1' )then
          cVar2S13S48N003P026P008nsss(0) <='1';
          else
          cVar2S13S48N003P026P008nsss(0) <='0';
          end if;
        if(cVar1S14S48P019N059P061P033(0)='1' AND  A(21)='0' AND E(17)='0' AND A(20)='0' )then
          cVar2S14S48P016P065P018nsss(0) <='1';
          else
          cVar2S14S48P016P065P018nsss(0) <='0';
          end if;
        if(cVar1S15S48P019N059P061P033(0)='1' AND  A(21)='1' AND D(16)='1' AND A(23)='0' )then
          cVar2S15S48P016P067P012nsss(0) <='1';
          else
          cVar2S15S48P016P067P012nsss(0) <='0';
          end if;
        if(cVar1S16S48P019N059P061P018(0)='1' AND  B(21)='0' AND A(13)='1' )then
          cVar2S16S48P034P013nsss(0) <='1';
          else
          cVar2S16S48P034P013nsss(0) <='0';
          end if;
        if(cVar1S17S48P019N059P061P018(0)='1' AND  B(21)='0' AND A(13)='0' AND D(16)='0' )then
          cVar2S17S48P034N013P067nsss(0) <='1';
          else
          cVar2S17S48P034N013P067nsss(0) <='0';
          end if;
        if(cVar1S0S49P019P033P057P013(0)='1' AND  B(21)='1' AND B(22)='0' AND A(12)='0' )then
          cVar2S0S49P034P032P015nsss(0) <='1';
          else
          cVar2S0S49P034P032P015nsss(0) <='0';
          end if;
        if(cVar1S1S49P019P033P057P013(0)='1' AND  B(21)='0' AND B(24)='1' AND A(24)='1' )then
          cVar2S1S49N034P028P010nsss(0) <='1';
          else
          cVar2S1S49N034P028P010nsss(0) <='0';
          end if;
        if(cVar1S2S49P019P033P057P013(0)='1' AND  B(21)='0' AND B(24)='0' )then
          cVar2S2S49N034N028psss(0) <='1';
          else
          cVar2S2S49N034N028psss(0) <='0';
          end if;
        if(cVar1S3S49P019P033P057P013(0)='1' AND  D(23)='0' AND D( 9)='0' AND E(18)='1' )then
          cVar2S3S49P039P062P061nsss(0) <='1';
          else
          cVar2S3S49P039P062P061nsss(0) <='0';
          end if;
        if(cVar1S4S49P019P033P057P030(0)='1' AND  E( 8)='0' )then
          cVar2S4S49P068nsss(0) <='1';
          else
          cVar2S4S49P068nsss(0) <='0';
          end if;
        if(cVar1S5S49P019P033P057N030(0)='1' AND  B(21)='0' AND E(20)='0' AND A(20)='0' )then
          cVar2S5S49P034P053P018nsss(0) <='1';
          else
          cVar2S5S49P034P053P018nsss(0) <='0';
          end if;
        if(cVar1S6S49P019P033P016P065(0)='1' AND  A(11)='1' AND B(10)='0' AND B(11)='0' )then
          cVar2S6S49P017P037P035nsss(0) <='1';
          else
          cVar2S6S49P017P037P035nsss(0) <='0';
          end if;
        if(cVar1S7S49P019P033P016P065(0)='1' AND  A(11)='0' AND D( 8)='1' )then
          cVar2S7S49N017P066nsss(0) <='1';
          else
          cVar2S7S49N017P066nsss(0) <='0';
          end if;
        if(cVar1S8S49P019P033P016P067(0)='1' AND  D( 8)='0' AND A(22)='0' )then
          cVar2S8S49P066P014nsss(0) <='1';
          else
          cVar2S8S49P066P014nsss(0) <='0';
          end if;
        if(cVar1S9S49P019P033P016N067(0)='1' AND  A(13)='1' AND A(22)='0' )then
          cVar2S9S49P013P014nsss(0) <='1';
          else
          cVar2S9S49P013P014nsss(0) <='0';
          end if;
        if(cVar1S11S49N019P007N025P059(0)='1' AND  D(11)='0' AND E(17)='0' )then
          cVar2S11S49P054P065nsss(0) <='1';
          else
          cVar2S11S49P054P065nsss(0) <='0';
          end if;
        if(cVar1S12S49N019P007N025P059(0)='1' AND  D(11)='0' AND E(17)='1' AND B(21)='1' )then
          cVar2S12S49P054P065P034nsss(0) <='1';
          else
          cVar2S12S49P054P065P034nsss(0) <='0';
          end if;
        if(cVar1S13S49N019N007P060P004(0)='1' AND  A(19)='0' AND B(12)='1' AND B(10)='0' )then
          cVar2S13S49P001P033P037nsss(0) <='1';
          else
          cVar2S13S49P001P033P037nsss(0) <='0';
          end if;
        if(cVar1S14S49N019N007P060P004(0)='1' AND  A(19)='0' AND B(12)='0' AND B(22)='1' )then
          cVar2S14S49P001N033P032nsss(0) <='1';
          else
          cVar2S14S49P001N033P032nsss(0) <='0';
          end if;
        if(cVar1S15S49N019N007N060P057(0)='1' AND  A(24)='1' AND B(24)='1' )then
          cVar2S15S49P010P028nsss(0) <='1';
          else
          cVar2S15S49P010P028nsss(0) <='0';
          end if;
        if(cVar1S16S49N019N007N060P057(0)='1' AND  A(24)='1' AND B(24)='0' AND B(23)='1' )then
          cVar2S16S49P010N028P030nsss(0) <='1';
          else
          cVar2S16S49P010N028P030nsss(0) <='0';
          end if;
        if(cVar1S17S49N019N007N060P057(0)='1' AND  A(24)='0' AND B(20)='1' )then
          cVar2S17S49N010P036nsss(0) <='1';
          else
          cVar2S17S49N010P036nsss(0) <='0';
          end if;
        if(cVar1S18S49N019N007N060P057(0)='1' AND  A(24)='0' AND B(20)='0' AND B(22)='1' )then
          cVar2S18S49N010N036P032nsss(0) <='1';
          else
          cVar2S18S49N010N036P032nsss(0) <='0';
          end if;
        if(cVar1S19S49N019N007N060N057(0)='1' AND  B(23)='0' AND A(13)='1' AND B(13)='1' )then
          cVar2S19S49P030P013P031nsss(0) <='1';
          else
          cVar2S19S49P030P013P031nsss(0) <='0';
          end if;
        if(cVar1S20S49N019N007N060N057(0)='1' AND  B(23)='1' AND A(23)='1' AND A(22)='0' )then
          cVar2S20S49P030P012P014nsss(0) <='1';
          else
          cVar2S20S49P030P012P014nsss(0) <='0';
          end if;
        if(cVar1S1S50P019P014P027N009(0)='1' AND  B(10)='0' AND B(25)='0' )then
          cVar2S1S50P037P026nsss(0) <='1';
          else
          cVar2S1S50P037P026nsss(0) <='0';
          end if;
        if(cVar1S2S50P019P014N027P050(0)='1' AND  B(20)='1' )then
          cVar2S2S50P036nsss(0) <='1';
          else
          cVar2S2S50P036nsss(0) <='0';
          end if;
        if(cVar1S3S50P019P014N027P050(0)='1' AND  B(20)='0' AND A(13)='0' AND B(13)='0' )then
          cVar2S3S50N036P013P031nsss(0) <='1';
          else
          cVar2S3S50N036P013P031nsss(0) <='0';
          end if;
        if(cVar1S4S50P019P014N027P050(0)='1' AND  B(20)='0' AND A(13)='1' AND A(24)='1' )then
          cVar2S4S50N036P013P010nsss(0) <='1';
          else
          cVar2S4S50N036P013P010nsss(0) <='0';
          end if;
        if(cVar1S5S50P019P014N027P050(0)='1' AND  A(27)='0' AND B(14)='1' )then
          cVar2S5S50P004P029nsss(0) <='1';
          else
          cVar2S5S50P004P029nsss(0) <='0';
          end if;
        if(cVar1S6S50P019P014P030P063(0)='1' AND  A(14)='1' AND A(26)='0' AND A(28)='0' )then
          cVar2S6S50P011P006P002nsss(0) <='1';
          else
          cVar2S6S50P011P006P002nsss(0) <='0';
          end if;
        if(cVar1S7S50P019P014P030P063(0)='1' AND  A(14)='0' AND D(11)='0' AND B(20)='0' )then
          cVar2S7S50N011P054P036nsss(0) <='1';
          else
          cVar2S7S50N011P054P036nsss(0) <='0';
          end if;
        if(cVar1S8S50P019P014P030P063(0)='1' AND  A(14)='0' AND D(11)='1' AND A(20)='1' )then
          cVar2S8S50N011P054P018nsss(0) <='1';
          else
          cVar2S8S50N011P054P018nsss(0) <='0';
          end if;
        if(cVar1S9S50P019P014P030P063(0)='1' AND  E(17)='1' AND A(26)='0' AND B(10)='1' )then
          cVar2S9S50P065P006P037nsss(0) <='1';
          else
          cVar2S9S50P065P006P037nsss(0) <='0';
          end if;
        if(cVar1S11S50P019P002P020P013(0)='1' AND  D( 9)='0' AND D(23)='0' AND D(22)='0' )then
          cVar2S11S50P062P039P043nsss(0) <='1';
          else
          cVar2S11S50P062P039P043nsss(0) <='0';
          end if;
        if(cVar1S12S50P019P002P020P013(0)='1' AND  D( 9)='1' AND E( 9)='1' AND A(25)='1' )then
          cVar2S12S50P062P064P008nsss(0) <='1';
          else
          cVar2S12S50P062P064P008nsss(0) <='0';
          end if;
        if(cVar1S13S50P019P002P020N013(0)='1' AND  B(21)='1' AND B(22)='0' )then
          cVar2S13S50P034P032nsss(0) <='1';
          else
          cVar2S13S50P034P032nsss(0) <='0';
          end if;
        if(cVar1S14S50P019P002P020N013(0)='1' AND  B(21)='0' AND E(16)='1' AND A(23)='1' )then
          cVar2S14S50N034P069P012nsss(0) <='1';
          else
          cVar2S14S50N034P069P012nsss(0) <='0';
          end if;
        if(cVar1S15S50P019P002P020P013(0)='1' AND  A(23)='0' AND E( 8)='1' )then
          cVar2S15S50P012P068nsss(0) <='1';
          else
          cVar2S15S50P012P068nsss(0) <='0';
          end if;
        if(cVar1S16S50P019P002P054P009(0)='1' AND  B(20)='1' AND A(24)='0' )then
          cVar2S16S50P036P010nsss(0) <='1';
          else
          cVar2S16S50P036P010nsss(0) <='0';
          end if;
        if(cVar1S17S50P019P002P054P009(0)='1' AND  B(20)='0' AND A(25)='1' AND A(12)='1' )then
          cVar2S17S50N036P008P015nsss(0) <='1';
          else
          cVar2S17S50N036P008P015nsss(0) <='0';
          end if;
        if(cVar1S0S51P019P002P020P039(0)='1' AND  E(15)='0' AND D(15)='0' AND B(18)='0' )then
          cVar2S0S51P040P038P021nsss(0) <='1';
          else
          cVar2S0S51P040P038P021nsss(0) <='0';
          end if;
        if(cVar1S1S51P019P002P020P039(0)='1' AND  E(15)='1' AND D( 8)='1' )then
          cVar2S1S51P040P066nsss(0) <='1';
          else
          cVar2S1S51P040P066nsss(0) <='0';
          end if;
        if(cVar1S2S51P019P002P020P039(0)='1' AND  A(23)='0' AND A(13)='0' AND A(21)='0' )then
          cVar2S2S51P012P013P016nsss(0) <='1';
          else
          cVar2S2S51P012P013P016nsss(0) <='0';
          end if;
        if(cVar1S3S51P019P002P020P013(0)='1' AND  A(23)='0' AND E( 8)='1' )then
          cVar2S3S51P012P068nsss(0) <='1';
          else
          cVar2S3S51P012P068nsss(0) <='0';
          end if;
        if(cVar1S4S51P019P002P054P000(0)='1' AND  B(20)='1' AND A(24)='0' )then
          cVar2S4S51P036P010nsss(0) <='1';
          else
          cVar2S4S51P036P010nsss(0) <='0';
          end if;
        if(cVar1S5S51P019P002P054P000(0)='1' AND  B(20)='0' AND A(25)='1' AND A(21)='0' )then
          cVar2S5S51N036P008P016nsss(0) <='1';
          else
          cVar2S5S51N036P008P016nsss(0) <='0';
          end if;
        if(cVar1S6S51P019P002P054P000(0)='1' AND  B(20)='0' AND A(25)='0' AND D( 8)='1' )then
          cVar2S6S51N036N008P066nsss(0) <='1';
          else
          cVar2S6S51N036N008P066nsss(0) <='0';
          end if;
        if(cVar1S7S51N019P017P042P015(0)='1' AND  A(23)='1' AND D(12)='0' AND A(27)='0' )then
          cVar2S7S51P012P050P004nsss(0) <='1';
          else
          cVar2S7S51P012P050P004nsss(0) <='0';
          end if;
        if(cVar1S8S51N019P017P042P015(0)='1' AND  A(23)='0' AND D(12)='1' AND A(22)='0' )then
          cVar2S8S51N012P050P014nsss(0) <='1';
          else
          cVar2S8S51N012P050P014nsss(0) <='0';
          end if;
        if(cVar1S9S51N019P017P042P015(0)='1' AND  A(23)='0' AND D(12)='0' AND E(18)='1' )then
          cVar2S9S51N012N050P061nsss(0) <='1';
          else
          cVar2S9S51N012N050P061nsss(0) <='0';
          end if;
        if(cVar1S10S51N019P017P042P015(0)='1' AND  E(18)='0' AND B(12)='0' AND A(28)='0' )then
          cVar2S10S51P061P033P002nsss(0) <='1';
          else
          cVar2S10S51P061P033P002nsss(0) <='0';
          end if;
        if(cVar1S12S51N019N017P005N023(0)='1' AND  B(18)='1' )then
          cVar2S12S51P021nsss(0) <='1';
          else
          cVar2S12S51P021nsss(0) <='0';
          end if;
        if(cVar1S13S51N019N017P005N023(0)='1' AND  B(18)='0' AND A(26)='0' AND D(11)='0' )then
          cVar2S13S51N021P006P054nsss(0) <='1';
          else
          cVar2S13S51N021P006P054nsss(0) <='0';
          end if;
        if(cVar1S14S51N019N017N005P012(0)='1' AND  B(23)='0' AND D(13)='1' )then
          cVar2S14S51P030P046nsss(0) <='1';
          else
          cVar2S14S51P030P046nsss(0) <='0';
          end if;
        if(cVar1S15S51N019N017N005P012(0)='1' AND  B(23)='0' AND D(13)='0' AND B(13)='1' )then
          cVar2S15S51P030N046P031nsss(0) <='1';
          else
          cVar2S15S51P030N046P031nsss(0) <='0';
          end if;
        if(cVar1S16S51N019N017N005P012(0)='1' AND  B(23)='1' AND E(19)='1' )then
          cVar2S16S51P030P057nsss(0) <='1';
          else
          cVar2S16S51P030P057nsss(0) <='0';
          end if;
        if(cVar1S17S51N019N017N005P012(0)='1' AND  B(23)='1' AND E(19)='0' AND A(12)='1' )then
          cVar2S17S51P030N057P015nsss(0) <='1';
          else
          cVar2S17S51P030N057P015nsss(0) <='0';
          end if;
        if(cVar1S18S51N019N017N005P012(0)='1' AND  E(19)='1' AND A(24)='0' )then
          cVar2S18S51P057P010nsss(0) <='1';
          else
          cVar2S18S51P057P010nsss(0) <='0';
          end if;
        if(cVar1S19S51N019N017N005P012(0)='1' AND  E(19)='0' AND A(29)='1' AND B(10)='0' )then
          cVar2S19S51N057P000P037nsss(0) <='1';
          else
          cVar2S19S51N057P000P037nsss(0) <='0';
          end if;
        if(cVar1S20S51N019N017N005P012(0)='1' AND  E(19)='0' AND A(29)='0' AND A(13)='1' )then
          cVar2S20S51N057N000P013nsss(0) <='1';
          else
          cVar2S20S51N057N000P013nsss(0) <='0';
          end if;
        if(cVar1S0S52P019P012P030P050(0)='1' AND  A(27)='0' AND E(13)='1' )then
          cVar2S0S52P004P048nsss(0) <='1';
          else
          cVar2S0S52P004P048nsss(0) <='0';
          end if;
        if(cVar1S1S52P019P012P030P050(0)='1' AND  A(27)='0' AND E(13)='0' AND E(12)='1' )then
          cVar2S1S52P004N048P052nsss(0) <='1';
          else
          cVar2S1S52P004N048P052nsss(0) <='0';
          end if;
        if(cVar1S2S52P019P012P030N050(0)='1' AND  E(13)='0' AND B(15)='0' )then
          cVar2S2S52P048P027nsss(0) <='1';
          else
          cVar2S2S52P048P027nsss(0) <='0';
          end if;
        if(cVar1S3S52P019P012P030N050(0)='1' AND  E(13)='0' AND B(15)='1' AND A(15)='1' )then
          cVar2S3S52P048P027P009nsss(0) <='1';
          else
          cVar2S3S52P048P027P009nsss(0) <='0';
          end if;
        if(cVar1S4S52P019P012P030N050(0)='1' AND  E(13)='1' AND B(16)='1' )then
          cVar2S4S52P048P025nsss(0) <='1';
          else
          cVar2S4S52P048P025nsss(0) <='0';
          end if;
        if(cVar1S5S52P019P012P030N050(0)='1' AND  E(13)='1' AND B(16)='0' AND D(13)='1' )then
          cVar2S5S52P048N025P046nsss(0) <='1';
          else
          cVar2S5S52P048N025P046nsss(0) <='0';
          end if;
        if(cVar1S6S52P019P012P030P010(0)='1' AND  A(22)='0' )then
          cVar2S6S52P014nsss(0) <='1';
          else
          cVar2S6S52P014nsss(0) <='0';
          end if;
        if(cVar1S7S52P019P012P030N010(0)='1' AND  A(21)='1' AND A(11)='1' )then
          cVar2S7S52P016P017nsss(0) <='1';
          else
          cVar2S7S52P016P017nsss(0) <='0';
          end if;
        if(cVar1S8S52P019P012P030N010(0)='1' AND  A(21)='0' AND E(19)='1' )then
          cVar2S8S52N016P057nsss(0) <='1';
          else
          cVar2S8S52N016P057nsss(0) <='0';
          end if;
        if(cVar1S9S52P019P012P008P031(0)='1' AND  D(10)='1' )then
          cVar2S9S52P058nsss(0) <='1';
          else
          cVar2S9S52P058nsss(0) <='0';
          end if;
        if(cVar1S10S52P019P012P008P031(0)='1' AND  D(10)='0' AND A(22)='0' )then
          cVar2S10S52N058P014nsss(0) <='1';
          else
          cVar2S10S52N058P014nsss(0) <='0';
          end if;
        if(cVar1S11S52P019P012P008N031(0)='1' AND  B(23)='1' AND A(22)='0' )then
          cVar2S11S52P030P014nsss(0) <='1';
          else
          cVar2S11S52P030P014nsss(0) <='0';
          end if;
        if(cVar1S12S52P019P012P008N031(0)='1' AND  B(23)='0' AND A(29)='1' AND B(20)='0' )then
          cVar2S12S52N030P000P036nsss(0) <='1';
          else
          cVar2S12S52N030P000P036nsss(0) <='0';
          end if;
        if(cVar1S13S52P019P012P008N031(0)='1' AND  B(23)='0' AND A(29)='0' AND A(28)='1' )then
          cVar2S13S52N030N000P002nsss(0) <='1';
          else
          cVar2S13S52N030N000P002nsss(0) <='0';
          end if;
        if(cVar1S14S52P019P012P008P011(0)='1' AND  D(12)='0' AND D(18)='1' )then
          cVar2S14S52P050P059nsss(0) <='1';
          else
          cVar2S14S52P050P059nsss(0) <='0';
          end if;
        if(cVar1S15S52P019P033P049P028(0)='1' AND  A(24)='1' AND A(23)='0' )then
          cVar2S15S52P010P012nsss(0) <='1';
          else
          cVar2S15S52P010P012nsss(0) <='0';
          end if;
        if(cVar1S16S52P019P033P049P028(0)='1' AND  A(24)='0' AND A(15)='0' AND A(14)='1' )then
          cVar2S16S52N010P009P011nsss(0) <='1';
          else
          cVar2S16S52N010P009P011nsss(0) <='0';
          end if;
        if(cVar1S17S52P019P033P049P068(0)='1' AND  A(21)='0' )then
          cVar2S17S52P016nsss(0) <='1';
          else
          cVar2S17S52P016nsss(0) <='0';
          end if;
        if(cVar1S18S52P019P033P016P065(0)='1' AND  A(11)='1' AND B(10)='0' )then
          cVar2S18S52P017P037nsss(0) <='1';
          else
          cVar2S18S52P017P037nsss(0) <='0';
          end if;
        if(cVar1S19S52P019P033P016P065(0)='1' AND  A(11)='0' AND A(23)='0' AND D( 8)='1' )then
          cVar2S19S52N017P012P066nsss(0) <='1';
          else
          cVar2S19S52N017P012P066nsss(0) <='0';
          end if;
        if(cVar1S20S52P019P033P016P067(0)='1' AND  A(11)='1' )then
          cVar2S20S52P017nsss(0) <='1';
          else
          cVar2S20S52P017nsss(0) <='0';
          end if;
        if(cVar1S0S53P019P033P049P048(0)='1' AND  A(24)='0' AND D(13)='0' )then
          cVar2S0S53P010P046nsss(0) <='1';
          else
          cVar2S0S53P010P046nsss(0) <='0';
          end if;
        if(cVar1S1S53P019P033P049P048(0)='1' AND  A(24)='1' AND A(23)='0' AND B(24)='1' )then
          cVar2S1S53P010P012P028nsss(0) <='1';
          else
          cVar2S1S53P010P012P028nsss(0) <='0';
          end if;
        if(cVar1S2S53P019P033P049P048(0)='1' AND  B(25)='1' )then
          cVar2S2S53P026nsss(0) <='1';
          else
          cVar2S2S53P026nsss(0) <='0';
          end if;
        if(cVar1S3S53P019P033P049P048(0)='1' AND  B(25)='0' AND B(10)='0' AND A(22)='1' )then
          cVar2S3S53N026P037P014nsss(0) <='1';
          else
          cVar2S3S53N026P037P014nsss(0) <='0';
          end if;
        if(cVar1S4S53P019P033P049P068(0)='1' AND  A(25)='1' )then
          cVar2S4S53P008nsss(0) <='1';
          else
          cVar2S4S53P008nsss(0) <='0';
          end if;
        if(cVar1S5S53P019P033P049P068(0)='1' AND  A(25)='0' AND D(21)='1' )then
          cVar2S5S53N008P047nsss(0) <='1';
          else
          cVar2S5S53N008P047nsss(0) <='0';
          end if;
        if(cVar1S6S53P019P033P016P065(0)='1' AND  E(10)='1' AND A(12)='1' )then
          cVar2S6S53P060P015nsss(0) <='1';
          else
          cVar2S6S53P060P015nsss(0) <='0';
          end if;
        if(cVar1S7S53P019P033P016P065(0)='1' AND  E(10)='0' AND E( 9)='0' AND A(11)='1' )then
          cVar2S7S53N060P064P017nsss(0) <='1';
          else
          cVar2S7S53N060P064P017nsss(0) <='0';
          end if;
        if(cVar1S8S53P019P033P016P067(0)='1' AND  D( 8)='0' AND A(22)='0' )then
          cVar2S8S53P066P014nsss(0) <='1';
          else
          cVar2S8S53P066P014nsss(0) <='0';
          end if;
        if(cVar1S10S53N019P050P021N027(0)='1' AND  D(23)='0' AND A(16)='0' AND B(22)='0' )then
          cVar2S10S53P039P007P032nsss(0) <='1';
          else
          cVar2S10S53P039P007P032nsss(0) <='0';
          end if;
        if(cVar1S11S53N019N050P032P008(0)='1' AND  E(10)='1' )then
          cVar2S11S53P060nsss(0) <='1';
          else
          cVar2S11S53P060nsss(0) <='0';
          end if;
        if(cVar1S12S53N019N050P032P008(0)='1' AND  E(10)='0' AND E(16)='1' )then
          cVar2S12S53N060P069nsss(0) <='1';
          else
          cVar2S12S53N060P069nsss(0) <='0';
          end if;
        if(cVar1S13S53N019N050P032P008(0)='1' AND  E(10)='0' AND E(16)='0' AND A(21)='1' )then
          cVar2S13S53N060N069P016nsss(0) <='1';
          else
          cVar2S13S53N060N069P016nsss(0) <='0';
          end if;
        if(cVar1S14S53N019N050N032P023(0)='1' AND  D(14)='1' )then
          cVar2S14S53P042nsss(0) <='1';
          else
          cVar2S14S53P042nsss(0) <='0';
          end if;
        if(cVar1S15S53N019N050N032P023(0)='1' AND  D(14)='0' AND E(22)='1' )then
          cVar2S15S53N042P045nsss(0) <='1';
          else
          cVar2S15S53N042P045nsss(0) <='0';
          end if;
        if(cVar1S16S53N019N050N032N023(0)='1' AND  D(14)='0' AND E(14)='0' AND D(13)='1' )then
          cVar2S16S53P042P044P046nsss(0) <='1';
          else
          cVar2S16S53P042P044P046nsss(0) <='0';
          end if;
        if(cVar1S17S53N019N050N032N023(0)='1' AND  D(14)='1' AND E(17)='1' )then
          cVar2S17S53P042P065nsss(0) <='1';
          else
          cVar2S17S53P042P065nsss(0) <='0';
          end if;
        if(cVar1S0S54P019P015P017P012(0)='1' AND  D(12)='0' AND A(27)='0' )then
          cVar2S0S54P050P004nsss(0) <='1';
          else
          cVar2S0S54P050P004nsss(0) <='0';
          end if;
        if(cVar1S1S54P019P015P017N012(0)='1' AND  D(14)='0' AND E(17)='1' AND E( 9)='0' )then
          cVar2S1S54P042P065P064nsss(0) <='1';
          else
          cVar2S1S54P042P065P064nsss(0) <='0';
          end if;
        if(cVar1S2S54P019P015P017N012(0)='1' AND  D(14)='0' AND E(17)='0' )then
          cVar2S2S54P042N065psss(0) <='1';
          else
          cVar2S2S54P042N065psss(0) <='0';
          end if;
        if(cVar1S3S54P019P015N017P063(0)='1' AND  B(21)='0' AND B(10)='0' )then
          cVar2S3S54P034P037nsss(0) <='1';
          else
          cVar2S3S54P034P037nsss(0) <='0';
          end if;
        if(cVar1S4S54P019P015N017P063(0)='1' AND  B(21)='1' AND B(10)='1' AND E( 8)='0' )then
          cVar2S4S54P034P037P068nsss(0) <='1';
          else
          cVar2S4S54P034P037P068nsss(0) <='0';
          end if;
        if(cVar1S5S54P019P015N017P063(0)='1' AND  B(11)='0' AND E(12)='1' )then
          cVar2S5S54P035P052nsss(0) <='1';
          else
          cVar2S5S54P035P052nsss(0) <='0';
          end if;
        if(cVar1S6S54P019P015P017P061(0)='1' AND  B(12)='1' )then
          cVar2S6S54P033nsss(0) <='1';
          else
          cVar2S6S54P033nsss(0) <='0';
          end if;
        if(cVar1S7S54P019P015P017P061(0)='1' AND  B(12)='0' AND A(14)='0' AND D(17)='1' )then
          cVar2S7S54N033P011P063nsss(0) <='1';
          else
          cVar2S7S54N033P011P063nsss(0) <='0';
          end if;
        if(cVar1S8S54P019P015P017N061(0)='1' AND  D(19)='1' )then
          cVar2S8S54P055nsss(0) <='1';
          else
          cVar2S8S54P055nsss(0) <='0';
          end if;
        if(cVar1S9S54P019P015P017N061(0)='1' AND  D(19)='0' AND D( 9)='1' AND B(11)='1' )then
          cVar2S9S54N055P062P035nsss(0) <='1';
          else
          cVar2S9S54N055P062P035nsss(0) <='0';
          end if;
        if(cVar1S10S54P019P015P017N061(0)='1' AND  D(19)='0' AND D( 9)='0' AND A(14)='1' )then
          cVar2S10S54N055N062P011nsss(0) <='1';
          else
          cVar2S10S54N055N062P011nsss(0) <='0';
          end if;
        if(cVar1S11S54P019P015P017P061(0)='1' AND  A(28)='0' AND A(21)='1' AND A(13)='1' )then
          cVar2S11S54P002P016P013nsss(0) <='1';
          else
          cVar2S11S54P002P016P013nsss(0) <='0';
          end if;
        if(cVar1S12S54P019P015P017P061(0)='1' AND  B(12)='1' )then
          cVar2S12S54P033nsss(0) <='1';
          else
          cVar2S12S54P033nsss(0) <='0';
          end if;
        if(cVar1S13S54P019P033P060P017(0)='1' AND  E( 9)='0' AND A(14)='0' )then
          cVar2S13S54P064P011nsss(0) <='1';
          else
          cVar2S13S54P064P011nsss(0) <='0';
          end if;
        if(cVar1S14S54P019P033P060P017(0)='1' AND  E( 9)='0' AND A(14)='1' AND A(12)='0' )then
          cVar2S14S54P064P011P015nsss(0) <='1';
          else
          cVar2S14S54P064P011P015nsss(0) <='0';
          end if;
        if(cVar1S15S54P019P033P060P017(0)='1' AND  E( 9)='1' AND A(14)='1' AND E(16)='1' )then
          cVar2S15S54P064P011P069nsss(0) <='1';
          else
          cVar2S15S54P064P011P069nsss(0) <='0';
          end if;
        if(cVar1S16S54P019P033P060N017(0)='1' AND  E( 9)='1' AND D(10)='0' AND A(18)='0' )then
          cVar2S16S54P064P058P003nsss(0) <='1';
          else
          cVar2S16S54P064P058P003nsss(0) <='0';
          end if;
        if(cVar1S17S54P019P033P060N017(0)='1' AND  E( 9)='0' AND B(24)='1' )then
          cVar2S17S54N064P028nsss(0) <='1';
          else
          cVar2S17S54N064P028nsss(0) <='0';
          end if;
        if(cVar1S18S54P019P033P060N017(0)='1' AND  E( 9)='0' AND B(24)='0' AND E(14)='1' )then
          cVar2S18S54N064N028P044nsss(0) <='1';
          else
          cVar2S18S54N064N028P044nsss(0) <='0';
          end if;
        if(cVar1S19S54P019P033P060P009(0)='1' AND  B(13)='1' )then
          cVar2S19S54P031nsss(0) <='1';
          else
          cVar2S19S54P031nsss(0) <='0';
          end if;
        if(cVar1S20S54P019P033P060P009(0)='1' AND  B(13)='0' AND B(22)='1' )then
          cVar2S20S54N031P032nsss(0) <='1';
          else
          cVar2S20S54N031P032nsss(0) <='0';
          end if;
        if(cVar1S21S54P019P033P016P065(0)='1' AND  E(10)='1' )then
          cVar2S21S54P060nsss(0) <='1';
          else
          cVar2S21S54P060nsss(0) <='0';
          end if;
        if(cVar1S22S54P019P033P016P065(0)='1' AND  E(10)='0' AND E( 9)='0' AND A(23)='0' )then
          cVar2S22S54N060P064P012nsss(0) <='1';
          else
          cVar2S22S54N060P064P012nsss(0) <='0';
          end if;
        if(cVar1S23S54P019P033P016P067(0)='1' AND  D( 8)='0' AND A(22)='0' )then
          cVar2S23S54P066P014nsss(0) <='1';
          else
          cVar2S23S54P066P014nsss(0) <='0';
          end if;
        if(cVar1S24S54P019P033P016N067(0)='1' AND  A(13)='1' AND A(22)='0' )then
          cVar2S24S54P013P014nsss(0) <='1';
          else
          cVar2S24S54P013P014nsss(0) <='0';
          end if;
        if(cVar1S0S55P015P068P051P022(0)='1' AND  A(29)='1' AND B(10)='1' )then
          cVar2S0S55P000P037nsss(0) <='1';
          else
          cVar2S0S55P000P037nsss(0) <='0';
          end if;
        if(cVar1S1S55P015P068P051P022(0)='1' AND  A(29)='1' AND B(10)='0' AND A(28)='0' )then
          cVar2S1S55P000N037P002nsss(0) <='1';
          else
          cVar2S1S55P000N037P002nsss(0) <='0';
          end if;
        if(cVar1S2S55P015P068P051P022(0)='1' AND  A(29)='0' AND A(27)='0' AND D(22)='0' )then
          cVar2S2S55N000P004P043nsss(0) <='1';
          else
          cVar2S2S55N000P004P043nsss(0) <='0';
          end if;
        if(cVar1S3S55P015P068P051P022(0)='1' AND  A(29)='0' AND A(27)='1' AND B(20)='0' )then
          cVar2S3S55N000P004P036nsss(0) <='1';
          else
          cVar2S3S55N000P004P036nsss(0) <='0';
          end if;
        if(cVar1S4S55P015P068P051P022(0)='1' AND  A(10)='1' AND A(21)='0' )then
          cVar2S4S55P019P016nsss(0) <='1';
          else
          cVar2S4S55P019P016nsss(0) <='0';
          end if;
        if(cVar1S5S55P015P068P051P053(0)='1' AND  A(26)='0' AND B(20)='1' )then
          cVar2S5S55P006P036nsss(0) <='1';
          else
          cVar2S5S55P006P036nsss(0) <='0';
          end if;
        if(cVar1S6S55P015P068P051P053(0)='1' AND  A(26)='0' AND B(20)='0' AND A(20)='0' )then
          cVar2S6S55P006N036P018nsss(0) <='1';
          else
          cVar2S6S55P006N036P018nsss(0) <='0';
          end if;
        if(cVar1S7S55P015P068P051N053(0)='1' AND  E(21)='1' AND A(22)='0' )then
          cVar2S7S55P049P014nsss(0) <='1';
          else
          cVar2S7S55P049P014nsss(0) <='0';
          end if;
        if(cVar1S8S55P015P068P009P010(0)='1' AND  A(29)='0' AND B(20)='0' AND A(25)='0' )then
          cVar2S8S55P000P036P008nsss(0) <='1';
          else
          cVar2S8S55P000P036P008nsss(0) <='0';
          end if;
        if(cVar1S9S55P015P068P009N010(0)='1' AND  A(26)='0' AND D(19)='0' AND A(25)='1' )then
          cVar2S9S55P006P055P008nsss(0) <='1';
          else
          cVar2S9S55P006P055P008nsss(0) <='0';
          end if;
        if(cVar1S10S55P015P068P009P066(0)='1' AND  D(11)='0' AND E(17)='1' )then
          cVar2S10S55P054P065nsss(0) <='1';
          else
          cVar2S10S55P054P065nsss(0) <='0';
          end if;
        if(cVar1S11S55N015P068P003P033(0)='1' AND  E(23)='0' AND B(28)='0' )then
          cVar2S11S55P041P020nsss(0) <='1';
          else
          cVar2S11S55P041P020nsss(0) <='0';
          end if;
        if(cVar1S12S55N015P068P003P033(0)='1' AND  E(23)='0' AND B(28)='1' AND A(10)='1' )then
          cVar2S12S55P041P020P019nsss(0) <='1';
          else
          cVar2S12S55P041P020P019nsss(0) <='0';
          end if;
        if(cVar1S13S55N015P068P003P033(0)='1' AND  A(25)='1' )then
          cVar2S13S55P008nsss(0) <='1';
          else
          cVar2S13S55P008nsss(0) <='0';
          end if;
        if(cVar1S14S55N015P068P003P033(0)='1' AND  A(25)='0' AND E(16)='0' AND E(10)='1' )then
          cVar2S14S55N008P069P060nsss(0) <='1';
          else
          cVar2S14S55N008P069P060nsss(0) <='0';
          end if;
        if(cVar1S15S55N015P068P003P065(0)='1' AND  A(15)='0' AND A(14)='0' AND D( 8)='0' )then
          cVar2S15S55P009P011P066nsss(0) <='1';
          else
          cVar2S15S55P009P011P066nsss(0) <='0';
          end if;
        if(cVar1S16S55N015N068P069P008(0)='1' AND  E(17)='1' AND A(24)='0' AND D(16)='1' )then
          cVar2S16S55P065P010P067nsss(0) <='1';
          else
          cVar2S16S55P065P010P067nsss(0) <='0';
          end if;
        if(cVar1S17S55N015N068P069P008(0)='1' AND  E(17)='0' AND A(21)='0' )then
          cVar2S17S55N065P016nsss(0) <='1';
          else
          cVar2S17S55N065P016nsss(0) <='0';
          end if;
        if(cVar1S18S55N015N068P069P008(0)='1' AND  E(17)='0' AND A(21)='1' AND B(20)='1' )then
          cVar2S18S55N065P016P036nsss(0) <='1';
          else
          cVar2S18S55N065P016P036nsss(0) <='0';
          end if;
        if(cVar1S19S55N015N068P069P008(0)='1' AND  D( 8)='0' AND B(26)='0' AND A(10)='1' )then
          cVar2S19S55P066P024P019nsss(0) <='1';
          else
          cVar2S19S55P066P024P019nsss(0) <='0';
          end if;
        if(cVar1S20S55N015N068N069P004(0)='1' AND  B(27)='1' )then
          cVar2S20S55P022nsss(0) <='1';
          else
          cVar2S20S55P022nsss(0) <='0';
          end if;
        if(cVar1S21S55N015N068N069P004(0)='1' AND  B(27)='0' AND A(21)='1' AND B(20)='0' )then
          cVar2S21S55N022P016P036nsss(0) <='1';
          else
          cVar2S21S55N022P016P036nsss(0) <='0';
          end if;
        if(cVar1S22S55N015N068N069N004(0)='1' AND  D(14)='0' AND E(14)='0' AND B(12)='1' )then
          cVar2S22S55P042P044P033nsss(0) <='1';
          else
          cVar2S22S55P042P044P033nsss(0) <='0';
          end if;
        if(cVar1S23S55N015N068N069N004(0)='1' AND  D(14)='1' AND A(17)='1' )then
          cVar2S23S55P042P005nsss(0) <='1';
          else
          cVar2S23S55P042P005nsss(0) <='0';
          end if;
        if(cVar1S24S55N015N068N069N004(0)='1' AND  D(14)='1' AND A(17)='0' AND A(23)='1' )then
          cVar2S24S55P042N005P012nsss(0) <='1';
          else
          cVar2S24S55P042N005P012nsss(0) <='0';
          end if;
        if(cVar1S0S56P068P015P066P034(0)='1' AND  D(17)='1' AND A(25)='0' )then
          cVar2S0S56P063P008nsss(0) <='1';
          else
          cVar2S0S56P063P008nsss(0) <='0';
          end if;
        if(cVar1S1S56P068P015P066P034(0)='1' AND  D(17)='0' AND D(16)='1' AND A(24)='0' )then
          cVar2S1S56N063P067P010nsss(0) <='1';
          else
          cVar2S1S56N063P067P010nsss(0) <='0';
          end if;
        if(cVar1S2S56P068P015P066P034(0)='1' AND  D(17)='0' AND D(16)='0' AND A(24)='1' )then
          cVar2S2S56N063N067P010nsss(0) <='1';
          else
          cVar2S2S56N063N067P010nsss(0) <='0';
          end if;
        if(cVar1S3S56P068P015P066N034(0)='1' AND  B(15)='1' AND A(15)='1' )then
          cVar2S3S56P027P009nsss(0) <='1';
          else
          cVar2S3S56P027P009nsss(0) <='0';
          end if;
        if(cVar1S4S56P068P015P066N034(0)='1' AND  B(15)='1' AND A(15)='0' AND A(13)='0' )then
          cVar2S4S56P027N009P013nsss(0) <='1';
          else
          cVar2S4S56P027N009P013nsss(0) <='0';
          end if;
        if(cVar1S5S56P068P015P066N034(0)='1' AND  B(15)='0' AND D(16)='0' )then
          cVar2S5S56N027P067nsss(0) <='1';
          else
          cVar2S5S56N027P067nsss(0) <='0';
          end if;
        if(cVar1S6S56P068P015P066N034(0)='1' AND  B(15)='0' AND D(16)='1' AND E(17)='1' )then
          cVar2S6S56N027P067P065nsss(0) <='1';
          else
          cVar2S6S56N027P067P065nsss(0) <='0';
          end if;
        if(cVar1S7S56P068P015P066P008(0)='1' AND  D(12)='0' AND E(10)='1' )then
          cVar2S7S56P050P060nsss(0) <='1';
          else
          cVar2S7S56P050P060nsss(0) <='0';
          end if;
        if(cVar1S8S56P068P015P051P022(0)='1' AND  A(29)='1' AND B(10)='1' )then
          cVar2S8S56P000P037nsss(0) <='1';
          else
          cVar2S8S56P000P037nsss(0) <='0';
          end if;
        if(cVar1S9S56P068P015P051P022(0)='1' AND  A(29)='1' AND B(10)='0' AND A(28)='0' )then
          cVar2S9S56P000N037P002nsss(0) <='1';
          else
          cVar2S9S56P000N037P002nsss(0) <='0';
          end if;
        if(cVar1S10S56P068P015P051P022(0)='1' AND  A(29)='0' AND A(21)='0' AND E(16)='1' )then
          cVar2S10S56N000P016P069nsss(0) <='1';
          else
          cVar2S10S56N000P016P069nsss(0) <='0';
          end if;
        if(cVar1S11S56P068P015P051P022(0)='1' AND  A(13)='0' AND A(10)='1' )then
          cVar2S11S56P013P019nsss(0) <='1';
          else
          cVar2S11S56P013P019nsss(0) <='0';
          end if;
        if(cVar1S12S56P068P015P051P053(0)='1' AND  A(26)='0' AND D(16)='0' )then
          cVar2S12S56P006P067nsss(0) <='1';
          else
          cVar2S12S56P006P067nsss(0) <='0';
          end if;
        if(cVar1S13S56P068P015P051N053(0)='1' AND  E(21)='1' AND A(22)='0' )then
          cVar2S13S56P049P014nsss(0) <='1';
          else
          cVar2S13S56P049P014nsss(0) <='0';
          end if;
        if(cVar1S14S56P068P009P024P052(0)='1' AND  A(21)='0' AND A(20)='0' )then
          cVar2S14S56P016P018nsss(0) <='1';
          else
          cVar2S14S56P016P018nsss(0) <='0';
          end if;
        if(cVar1S15S56P068P009P024P052(0)='1' AND  A(21)='1' )then
          cVar2S15S56P016psss(0) <='1';
          else
          cVar2S15S56P016psss(0) <='0';
          end if;
        if(cVar1S16S56P068P009P024N052(0)='1' AND  E( 9)='1' AND D(20)='0' )then
          cVar2S16S56P064P051nsss(0) <='1';
          else
          cVar2S16S56P064P051nsss(0) <='0';
          end if;
        if(cVar1S17S56P068P009P024N052(0)='1' AND  E( 9)='0' AND B(21)='0' AND E(11)='1' )then
          cVar2S17S56N064P034P056nsss(0) <='1';
          else
          cVar2S17S56N064P034P056nsss(0) <='0';
          end if;
        if(cVar1S19S56P068P009P024N006(0)='1' AND  A(21)='0' AND A(22)='0' AND A(20)='1' )then
          cVar2S19S56P016P014P018nsss(0) <='1';
          else
          cVar2S19S56P016P014P018nsss(0) <='0';
          end if;
        if(cVar1S20S56P068P009P002P066(0)='1' AND  D(12)='1' )then
          cVar2S20S56P050nsss(0) <='1';
          else
          cVar2S20S56P050nsss(0) <='0';
          end if;
        if(cVar1S21S56P068P009P002P066(0)='1' AND  D(12)='0' AND A(29)='0' AND A(14)='1' )then
          cVar2S21S56N050P000P011nsss(0) <='1';
          else
          cVar2S21S56N050P000P011nsss(0) <='0';
          end if;
        if(cVar1S0S57P015P051P009P037(0)='1' AND  D(16)='0' AND A(13)='1' AND D(17)='0' )then
          cVar2S0S57P067P013P063nsss(0) <='1';
          else
          cVar2S0S57P067P013P063nsss(0) <='0';
          end if;
        if(cVar1S1S57P015P051P009P037(0)='1' AND  D(16)='0' AND A(13)='0' )then
          cVar2S1S57P067N013psss(0) <='1';
          else
          cVar2S1S57P067N013psss(0) <='0';
          end if;
        if(cVar1S2S57P015P051P009P037(0)='1' AND  D(16)='1' AND B(12)='1' AND A(22)='0' )then
          cVar2S2S57P067P033P014nsss(0) <='1';
          else
          cVar2S2S57P067P033P014nsss(0) <='0';
          end if;
        if(cVar1S3S57P015P051P009P037(0)='1' AND  A(13)='0' AND A(20)='1' AND D(10)='0' )then
          cVar2S3S57P013P018P058nsss(0) <='1';
          else
          cVar2S3S57P013P018P058nsss(0) <='0';
          end if;
        if(cVar1S4S57P015P051P009P037(0)='1' AND  A(13)='0' AND A(20)='0' AND E(10)='1' )then
          cVar2S4S57P013N018P060nsss(0) <='1';
          else
          cVar2S4S57P013N018P060nsss(0) <='0';
          end if;
        if(cVar1S5S57P015P051P009P037(0)='1' AND  A(13)='1' AND A(11)='0' AND A(20)='1' )then
          cVar2S5S57P013P017P018nsss(0) <='1';
          else
          cVar2S5S57P013P017P018nsss(0) <='0';
          end if;
        if(cVar1S6S57P015P051P009P037(0)='1' AND  A(13)='1' AND A(11)='1' AND B(26)='1' )then
          cVar2S6S57P013P017P024nsss(0) <='1';
          else
          cVar2S6S57P013P017P024nsss(0) <='0';
          end if;
        if(cVar1S7S57P015P051P009P068(0)='1' AND  A(23)='0' AND A(13)='0' AND A(24)='0' )then
          cVar2S7S57P012P013P010nsss(0) <='1';
          else
          cVar2S7S57P012P013P010nsss(0) <='0';
          end if;
        if(cVar1S8S57P015P051P009P068(0)='1' AND  A(23)='0' AND A(13)='1' AND A(22)='1' )then
          cVar2S8S57P012P013P014nsss(0) <='1';
          else
          cVar2S8S57P012P013P014nsss(0) <='0';
          end if;
        if(cVar1S9S57P015P051P009P068(0)='1' AND  A(23)='1' AND A(21)='0' AND A(24)='1' )then
          cVar2S9S57P012P016P010nsss(0) <='1';
          else
          cVar2S9S57P012P016P010nsss(0) <='0';
          end if;
        if(cVar1S10S57P015P051P009P068(0)='1' AND  D( 8)='1' AND E(17)='1' )then
          cVar2S10S57P066P065nsss(0) <='1';
          else
          cVar2S10S57P066P065nsss(0) <='0';
          end if;
        if(cVar1S11S57P015P051P053P000(0)='1' AND  A(26)='0' AND B(11)='0' )then
          cVar2S11S57P006P035nsss(0) <='1';
          else
          cVar2S11S57P006P035nsss(0) <='0';
          end if;
        if(cVar1S12S57P015P051N053P014(0)='1' AND  E(21)='1' )then
          cVar2S12S57P049nsss(0) <='1';
          else
          cVar2S12S57P049nsss(0) <='0';
          end if;
        if(cVar1S13S57N015P033P034P006(0)='1' AND  A(27)='0' )then
          cVar2S13S57P004nsss(0) <='1';
          else
          cVar2S13S57P004nsss(0) <='0';
          end if;
        if(cVar1S14S57N015P033P034P006(0)='1' AND  A(13)='0' AND A(22)='0' AND D(17)='1' )then
          cVar2S14S57P013P014P063nsss(0) <='1';
          else
          cVar2S14S57P013P014P063nsss(0) <='0';
          end if;
        if(cVar1S15S57N015P033N034P027(0)='1' AND  A(15)='1' )then
          cVar2S15S57P009nsss(0) <='1';
          else
          cVar2S15S57P009nsss(0) <='0';
          end if;
        if(cVar1S16S57N015P033N034P027(0)='1' AND  A(15)='0' AND A(18)='1' )then
          cVar2S16S57N009P003nsss(0) <='1';
          else
          cVar2S16S57N009P003nsss(0) <='0';
          end if;
        if(cVar1S17S57N015P033N034N027(0)='1' AND  D( 8)='1' AND A(18)='0' )then
          cVar2S17S57P066P003nsss(0) <='1';
          else
          cVar2S17S57P066P003nsss(0) <='0';
          end if;
        if(cVar1S18S57N015P033N034N027(0)='1' AND  D( 8)='0' AND B(11)='1' )then
          cVar2S18S57N066P035nsss(0) <='1';
          else
          cVar2S18S57N066P035nsss(0) <='0';
          end if;
        if(cVar1S19S57N015P033N034N027(0)='1' AND  D( 8)='0' AND B(11)='0' AND B(28)='1' )then
          cVar2S19S57N066N035P020nsss(0) <='1';
          else
          cVar2S19S57N066N035P020nsss(0) <='0';
          end if;
        if(cVar1S20S57N015P033P064P056(0)='1' AND  B(26)='0' AND A(28)='0' AND A(13)='1' )then
          cVar2S20S57P024P002P013nsss(0) <='1';
          else
          cVar2S20S57P024P002P013nsss(0) <='0';
          end if;
        if(cVar1S0S58P066P015P033P018(0)='1' AND  A(27)='1' AND B(27)='1' )then
          cVar2S0S58P004P022nsss(0) <='1';
          else
          cVar2S0S58P004P022nsss(0) <='0';
          end if;
        if(cVar1S1S58P066P015P033P018(0)='1' AND  A(27)='1' AND B(27)='0' AND A(21)='1' )then
          cVar2S1S58P004N022P016nsss(0) <='1';
          else
          cVar2S1S58P004N022P016nsss(0) <='0';
          end if;
        if(cVar1S2S58P066P015P033P018(0)='1' AND  A(27)='0' AND D(14)='0' )then
          cVar2S2S58N004P042nsss(0) <='1';
          else
          cVar2S2S58N004P042nsss(0) <='0';
          end if;
        if(cVar1S3S58P066P015P033P018(0)='1' AND  A(27)='0' AND D(14)='1' AND A(17)='1' )then
          cVar2S3S58N004P042P005nsss(0) <='1';
          else
          cVar2S3S58N004P042P005nsss(0) <='0';
          end if;
        if(cVar1S4S58P066P015P033P018(0)='1' AND  D(22)='0' AND A(18)='1' AND A(16)='0' )then
          cVar2S4S58P043P003P007nsss(0) <='1';
          else
          cVar2S4S58P043P003P007nsss(0) <='0';
          end if;
        if(cVar1S5S58P066P015P033P018(0)='1' AND  D(22)='0' AND A(18)='0' AND A(29)='1' )then
          cVar2S5S58P043N003P000nsss(0) <='1';
          else
          cVar2S5S58P043N003P000nsss(0) <='0';
          end if;
        if(cVar1S6S58P066P015P033P018(0)='1' AND  D(22)='1' AND E(22)='1' )then
          cVar2S6S58P043P045nsss(0) <='1';
          else
          cVar2S6S58P043P045nsss(0) <='0';
          end if;
        if(cVar1S7S58P066P015P033P018(0)='1' AND  A(10)='0' AND B(20)='1' )then
          cVar2S7S58P019P036nsss(0) <='1';
          else
          cVar2S7S58P019P036nsss(0) <='0';
          end if;
        if(cVar1S8S58P066P015P033P018(0)='1' AND  A(10)='0' AND B(20)='0' AND A(13)='0' )then
          cVar2S8S58P019N036P013nsss(0) <='1';
          else
          cVar2S8S58P019N036P013nsss(0) <='0';
          end if;
        if(cVar1S9S58P066P015P033P018(0)='1' AND  A(10)='1' AND A(11)='1' AND A(21)='0' )then
          cVar2S9S58P019P017P016nsss(0) <='1';
          else
          cVar2S9S58P019P017P016nsss(0) <='0';
          end if;
        if(cVar1S10S58P066P015P033N018(0)='1' AND  A(13)='1' AND A(23)='0' )then
          cVar2S10S58P013P012nsss(0) <='1';
          else
          cVar2S10S58P013P012nsss(0) <='0';
          end if;
        if(cVar1S11S58P066P015P007P068(0)='1' AND  E(20)='1' AND B(26)='0' AND A(14)='0' )then
          cVar2S11S58P053P024P011nsss(0) <='1';
          else
          cVar2S11S58P053P024P011nsss(0) <='0';
          end if;
        if(cVar1S12S58P066P015P007P068(0)='1' AND  E(20)='0' AND D(20)='0' AND E(16)='1' )then
          cVar2S12S58N053P051P069nsss(0) <='1';
          else
          cVar2S12S58N053P051P069nsss(0) <='0';
          end if;
        if(cVar1S13S58P066P015P007P068(0)='1' AND  E(20)='0' AND D(20)='1' AND A(25)='1' )then
          cVar2S13S58N053P051P008nsss(0) <='1';
          else
          cVar2S13S58N053P051P008nsss(0) <='0';
          end if;
        if(cVar1S14S58P066P015P007P068(0)='1' AND  A(15)='0' AND A(22)='0' AND A(10)='1' )then
          cVar2S14S58P009P014P019nsss(0) <='1';
          else
          cVar2S14S58P009P014P019nsss(0) <='0';
          end if;
        if(cVar1S15S58P066P015P007P059(0)='1' AND  B(23)='1' )then
          cVar2S15S58P030nsss(0) <='1';
          else
          cVar2S15S58P030nsss(0) <='0';
          end if;
        if(cVar1S16S58P066P009P024P045(0)='1' AND  E(18)='1' AND B(12)='1' )then
          cVar2S16S58P061P033nsss(0) <='1';
          else
          cVar2S16S58P061P033nsss(0) <='0';
          end if;
        if(cVar1S17S58P066P009P024P045(0)='1' AND  E(18)='1' AND B(12)='0' AND A(10)='1' )then
          cVar2S17S58P061N033P019nsss(0) <='1';
          else
          cVar2S17S58P061N033P019nsss(0) <='0';
          end if;
        if(cVar1S18S58P066P009P024P045(0)='1' AND  D(22)='1' )then
          cVar2S18S58P043nsss(0) <='1';
          else
          cVar2S18S58P043nsss(0) <='0';
          end if;
        if(cVar1S19S58P066P009P024P053(0)='1' AND  A(26)='1' )then
          cVar2S19S58P006nsss(0) <='1';
          else
          cVar2S19S58P006nsss(0) <='0';
          end if;
        if(cVar1S20S58P066P009P002P037(0)='1' AND  A(22)='1' AND A(11)='0' )then
          cVar2S20S58P014P017nsss(0) <='1';
          else
          cVar2S20S58P014P017nsss(0) <='0';
          end if;
        if(cVar1S21S58P066P009P002P037(0)='1' AND  A(22)='0' AND D( 9)='1' )then
          cVar2S21S58N014P062nsss(0) <='1';
          else
          cVar2S21S58N014P062nsss(0) <='0';
          end if;
        if(cVar1S22S58P066P009P002N037(0)='1' AND  B(22)='1' )then
          cVar2S22S58P032nsss(0) <='1';
          else
          cVar2S22S58P032nsss(0) <='0';
          end if;
        if(cVar1S0S59P018P008P050P067(0)='1' AND  A(21)='0' )then
          cVar2S0S59P016nsss(0) <='1';
          else
          cVar2S0S59P016nsss(0) <='0';
          end if;
        if(cVar1S1S59P018P008P050P067(0)='1' AND  A(21)='1' AND A(29)='1' )then
          cVar2S1S59P016P000nsss(0) <='1';
          else
          cVar2S1S59P016P000nsss(0) <='0';
          end if;
        if(cVar1S2S59P018P008P050P067(0)='1' AND  A(21)='1' AND A(29)='0' AND D(10)='1' )then
          cVar2S2S59P016N000P058nsss(0) <='1';
          else
          cVar2S2S59P016N000P058nsss(0) <='0';
          end if;
        if(cVar1S3S59P018P008P050N067(0)='1' AND  E(12)='0' AND D( 9)='0' AND E( 9)='0' )then
          cVar2S3S59P052P062P064nsss(0) <='1';
          else
          cVar2S3S59P052P062P064nsss(0) <='0';
          end if;
        if(cVar1S4S59P018P008P050N067(0)='1' AND  E(12)='0' AND D( 9)='1' AND B(10)='1' )then
          cVar2S4S59P052P062P037nsss(0) <='1';
          else
          cVar2S4S59P052P062P037nsss(0) <='0';
          end if;
        if(cVar1S5S59P018P008P050P009(0)='1' AND  A(12)='0' )then
          cVar2S5S59P015nsss(0) <='1';
          else
          cVar2S5S59P015nsss(0) <='0';
          end if;
        if(cVar1S6S59P018P008P050N009(0)='1' AND  B(26)='0' AND A(23)='0' AND E(13)='1' )then
          cVar2S6S59P024P012P048nsss(0) <='1';
          else
          cVar2S6S59P024P012P048nsss(0) <='0';
          end if;
        if(cVar1S7S59P018P008P054P015(0)='1' AND  A(28)='0' AND A(22)='0' )then
          cVar2S7S59P002P014nsss(0) <='1';
          else
          cVar2S7S59P002P014nsss(0) <='0';
          end if;
        if(cVar1S8S59P018P008P054P015(0)='1' AND  A(28)='0' AND A(22)='1' AND A(23)='0' )then
          cVar2S8S59P002P014P012nsss(0) <='1';
          else
          cVar2S8S59P002P014P012nsss(0) <='0';
          end if;
        if(cVar1S9S59P018P008P054P015(0)='1' AND  D(17)='1' AND E( 8)='1' )then
          cVar2S9S59P063P068nsss(0) <='1';
          else
          cVar2S9S59P063P068nsss(0) <='0';
          end if;
        if(cVar1S10S59P018P008P054P015(0)='1' AND  D(17)='0' AND A(21)='0' AND A(26)='1' )then
          cVar2S10S59N063P016P006nsss(0) <='1';
          else
          cVar2S10S59N063P016P006nsss(0) <='0';
          end if;
        if(cVar1S11S59N018P061P008P026(0)='1' AND  A(22)='0' )then
          cVar2S11S59P014nsss(0) <='1';
          else
          cVar2S11S59P014nsss(0) <='0';
          end if;
        if(cVar1S12S59N018P061P008N026(0)='1' AND  A(18)='0' AND A(17)='0' AND A(12)='1' )then
          cVar2S12S59P003P005P015nsss(0) <='1';
          else
          cVar2S12S59P003P005P015nsss(0) <='0';
          end if;
        if(cVar1S13S59N018P061P008N026(0)='1' AND  A(18)='1' AND A(23)='1' AND A(22)='1' )then
          cVar2S13S59P003P012P014nsss(0) <='1';
          else
          cVar2S13S59P003P012P014nsss(0) <='0';
          end if;
        if(cVar1S14S59N018P061N008P039(0)='1' AND  B(28)='1' )then
          cVar2S14S59P020nsss(0) <='1';
          else
          cVar2S14S59P020nsss(0) <='0';
          end if;
        if(cVar1S15S59N018P061N008P039(0)='1' AND  B(28)='0' AND A(23)='0' AND E(23)='1' )then
          cVar2S15S59N020P012P041nsss(0) <='1';
          else
          cVar2S15S59N020P012P041nsss(0) <='0';
          end if;
        if(cVar1S16S59N018P061N008N039(0)='1' AND  B(28)='0' AND E(19)='1' AND B(23)='1' )then
          cVar2S16S59P020P057P030nsss(0) <='1';
          else
          cVar2S16S59P020P057P030nsss(0) <='0';
          end if;
        if(cVar1S17S59N018P061N008N039(0)='1' AND  B(28)='1' AND A(28)='1' )then
          cVar2S17S59P020P002nsss(0) <='1';
          else
          cVar2S17S59P020P002nsss(0) <='0';
          end if;
        if(cVar1S18S59N018P061P059P000(0)='1' AND  A(15)='0' AND A(16)='0' )then
          cVar2S18S59P009P007nsss(0) <='1';
          else
          cVar2S18S59P009P007nsss(0) <='0';
          end if;
        if(cVar1S19S59N018P061N059P063(0)='1' AND  A(14)='0' AND A(22)='0' AND E(17)='0' )then
          cVar2S19S59P011P014P065nsss(0) <='1';
          else
          cVar2S19S59P011P014P065nsss(0) <='0';
          end if;
        if(cVar1S20S59N018P061N059N063(0)='1' AND  A(15)='1' )then
          cVar2S20S59P009nsss(0) <='1';
          else
          cVar2S20S59P009nsss(0) <='0';
          end if;
        if(cVar1S0S60P018P061P067P010(0)='1' AND  B(24)='1' )then
          cVar2S0S60P028nsss(0) <='1';
          else
          cVar2S0S60P028nsss(0) <='0';
          end if;
        if(cVar1S1S60P018P061P067P010(0)='1' AND  B(24)='0' AND D(10)='1' )then
          cVar2S1S60N028P058nsss(0) <='1';
          else
          cVar2S1S60N028P058nsss(0) <='0';
          end if;
        if(cVar1S2S60P018P061P067P010(0)='1' AND  B(24)='0' AND D(10)='0' AND D(14)='0' )then
          cVar2S2S60N028N058P042nsss(0) <='1';
          else
          cVar2S2S60N028N058P042nsss(0) <='0';
          end if;
        if(cVar1S3S60P018P061P067N010(0)='1' AND  A(27)='1' )then
          cVar2S3S60P004nsss(0) <='1';
          else
          cVar2S3S60P004nsss(0) <='0';
          end if;
        if(cVar1S4S60P018P061P067N010(0)='1' AND  A(27)='0' AND B(22)='1' )then
          cVar2S4S60N004P032nsss(0) <='1';
          else
          cVar2S4S60N004P032nsss(0) <='0';
          end if;
        if(cVar1S5S60P018P061P067N010(0)='1' AND  A(27)='0' AND B(22)='0' AND B(24)='0' )then
          cVar2S5S60N004N032P028nsss(0) <='1';
          else
          cVar2S5S60N004N032P028nsss(0) <='0';
          end if;
        if(cVar1S6S60P018P061P067P013(0)='1' AND  A(27)='0' AND E(22)='0' )then
          cVar2S6S60P004P045nsss(0) <='1';
          else
          cVar2S6S60P004P045nsss(0) <='0';
          end if;
        if(cVar1S7S60P018P061P067P013(0)='1' AND  B(26)='0' AND B(21)='1' AND A(22)='0' )then
          cVar2S7S60P024P034P014nsss(0) <='1';
          else
          cVar2S7S60P024P034P014nsss(0) <='0';
          end if;
        if(cVar1S8S60P018P061P059P000(0)='1' AND  A(15)='0' AND A(16)='0' AND B(22)='0' )then
          cVar2S8S60P009P007P032nsss(0) <='1';
          else
          cVar2S8S60P009P007P032nsss(0) <='0';
          end if;
        if(cVar1S9S60P018P061N059P063(0)='1' AND  E(10)='1' )then
          cVar2S9S60P060nsss(0) <='1';
          else
          cVar2S9S60P060nsss(0) <='0';
          end if;
        if(cVar1S10S60P018P061N059P063(0)='1' AND  E(10)='0' AND A(22)='0' AND E(17)='0' )then
          cVar2S10S60N060P014P065nsss(0) <='1';
          else
          cVar2S10S60N060P014P065nsss(0) <='0';
          end if;
        if(cVar1S11S60P018P061N059N063(0)='1' AND  A(15)='1' )then
          cVar2S11S60P009nsss(0) <='1';
          else
          cVar2S11S60P009nsss(0) <='0';
          end if;
        if(cVar1S13S60P018P067P019N056(0)='1' AND  A(22)='0' )then
          cVar2S13S60P014nsss(0) <='1';
          else
          cVar2S13S60P014nsss(0) <='0';
          end if;
        if(cVar1S14S60P018P067P019N056(0)='1' AND  A(22)='1' AND A(23)='1' AND E(16)='1' )then
          cVar2S14S60P014P012P069nsss(0) <='1';
          else
          cVar2S14S60P014P012P069nsss(0) <='0';
          end if;
        if(cVar1S15S60P018P067P019N056(0)='1' AND  A(22)='1' AND A(23)='0' AND E( 8)='1' )then
          cVar2S15S60P014N012P068nsss(0) <='1';
          else
          cVar2S15S60P014N012P068nsss(0) <='0';
          end if;
        if(cVar1S16S60P018P067P019P024(0)='1' AND  D(20)='0' AND E(17)='1' AND D( 9)='0' )then
          cVar2S16S60P051P065P062nsss(0) <='1';
          else
          cVar2S16S60P051P065P062nsss(0) <='0';
          end if;
        if(cVar1S17S60P018P067P019P024(0)='1' AND  D(20)='0' AND E(17)='0' AND B(25)='0' )then
          cVar2S17S60P051N065P026nsss(0) <='1';
          else
          cVar2S17S60P051N065P026nsss(0) <='0';
          end if;
        if(cVar1S18S60P018P067P019P024(0)='1' AND  D(20)='1' AND A(12)='1' )then
          cVar2S18S60P051P015nsss(0) <='1';
          else
          cVar2S18S60P051P015nsss(0) <='0';
          end if;
        if(cVar1S19S60P018N067P069P030(0)='1' AND  E(11)='0' AND A(29)='1' AND A(15)='0' )then
          cVar2S19S60P056P000P009nsss(0) <='1';
          else
          cVar2S19S60P056P000P009nsss(0) <='0';
          end if;
        if(cVar1S20S60P018N067P069P030(0)='1' AND  E(11)='1' AND B(21)='0' AND B(20)='1' )then
          cVar2S20S60P056P034P036nsss(0) <='1';
          else
          cVar2S20S60P056P034P036nsss(0) <='0';
          end if;
        if(cVar1S21S60P018N067P069P030(0)='1' AND  E(18)='0' AND A(15)='0' AND E( 8)='1' )then
          cVar2S21S60P061P009P068nsss(0) <='1';
          else
          cVar2S21S60P061P009P068nsss(0) <='0';
          end if;
        if(cVar1S22S60P018N067P069P014(0)='1' AND  D(17)='1' )then
          cVar2S22S60P063nsss(0) <='1';
          else
          cVar2S22S60P063nsss(0) <='0';
          end if;
        if(cVar1S0S61P018P008P024P034(0)='1' AND  E(18)='1' AND A(13)='1' )then
          cVar2S0S61P061P013nsss(0) <='1';
          else
          cVar2S0S61P061P013nsss(0) <='0';
          end if;
        if(cVar1S1S61P018P008P024P034(0)='1' AND  E(18)='1' AND A(13)='0' AND E(10)='0' )then
          cVar2S1S61P061N013P060nsss(0) <='1';
          else
          cVar2S1S61P061N013P060nsss(0) <='0';
          end if;
        if(cVar1S2S61P018P008P024P034(0)='1' AND  E(18)='0' AND B(13)='1' )then
          cVar2S2S61N061P031nsss(0) <='1';
          else
          cVar2S2S61N061P031nsss(0) <='0';
          end if;
        if(cVar1S3S61P018P008P024P034(0)='1' AND  E(18)='0' AND B(13)='0' AND E(16)='0' )then
          cVar2S3S61N061N031P069nsss(0) <='1';
          else
          cVar2S3S61N061N031P069nsss(0) <='0';
          end if;
        if(cVar1S4S61P018P008P024P034(0)='1' AND  E(11)='0' AND A(16)='0' AND D(10)='0' )then
          cVar2S4S61P056P007P058nsss(0) <='1';
          else
          cVar2S4S61P056P007P058nsss(0) <='0';
          end if;
        if(cVar1S6S61P018P008P024N045(0)='1' AND  A(22)='0' AND A(18)='1' )then
          cVar2S6S61P014P003nsss(0) <='1';
          else
          cVar2S6S61P014P003nsss(0) <='0';
          end if;
        if(cVar1S7S61P018P008P024N045(0)='1' AND  A(22)='1' AND A(10)='0' AND A(21)='1' )then
          cVar2S7S61P014P019P016nsss(0) <='1';
          else
          cVar2S7S61P014P019P016nsss(0) <='0';
          end if;
        if(cVar1S8S61P018P008P054P022(0)='1' AND  A(12)='0' AND A(28)='0' )then
          cVar2S8S61P015P002nsss(0) <='1';
          else
          cVar2S8S61P015P002nsss(0) <='0';
          end if;
        if(cVar1S9S61P018P008P054P022(0)='1' AND  A(12)='1' AND D(17)='1' AND E( 8)='1' )then
          cVar2S9S61P015P063P068nsss(0) <='1';
          else
          cVar2S9S61P015P063P068nsss(0) <='0';
          end if;
        if(cVar1S10S61N018P061P050P033(0)='1' AND  B(21)='0' AND A(25)='1' AND A(13)='0' )then
          cVar2S10S61P034P008P013nsss(0) <='1';
          else
          cVar2S10S61P034P008P013nsss(0) <='0';
          end if;
        if(cVar1S11S61N018P061P050P033(0)='1' AND  B(21)='0' AND A(25)='0' )then
          cVar2S11S61P034N008psss(0) <='1';
          else
          cVar2S11S61P034N008psss(0) <='0';
          end if;
        if(cVar1S12S61N018P061N050P004(0)='1' AND  B(27)='1' )then
          cVar2S12S61P022nsss(0) <='1';
          else
          cVar2S12S61P022nsss(0) <='0';
          end if;
        if(cVar1S13S61N018P061N050P004(0)='1' AND  B(27)='0' AND E(15)='1' )then
          cVar2S13S61N022P040nsss(0) <='1';
          else
          cVar2S13S61N022P040nsss(0) <='0';
          end if;
        if(cVar1S14S61N018P061N050P004(0)='1' AND  B(27)='0' AND E(15)='0' AND A(21)='1' )then
          cVar2S14S61N022N040P016nsss(0) <='1';
          else
          cVar2S14S61N022N040P016nsss(0) <='0';
          end if;
        if(cVar1S15S61N018P061N050N004(0)='1' AND  B(27)='0' AND B(24)='1' AND A(24)='1' )then
          cVar2S15S61P022P028P010nsss(0) <='1';
          else
          cVar2S15S61P022P028P010nsss(0) <='0';
          end if;
        if(cVar1S16S61N018P061N050N004(0)='1' AND  B(27)='1' AND D(22)='1' )then
          cVar2S16S61P022P043nsss(0) <='1';
          else
          cVar2S16S61P022P043nsss(0) <='0';
          end if;
        if(cVar1S17S61N018P061P059P000(0)='1' AND  A(16)='0' AND E(16)='1' AND D(17)='0' )then
          cVar2S17S61P007P069P063nsss(0) <='1';
          else
          cVar2S17S61P007P069P063nsss(0) <='0';
          end if;
        if(cVar1S18S61N018P061P059P000(0)='1' AND  A(16)='0' AND E(16)='0' AND B(20)='0' )then
          cVar2S18S61P007N069P036nsss(0) <='1';
          else
          cVar2S18S61P007N069P036nsss(0) <='0';
          end if;
        if(cVar1S19S61N018P061N059P063(0)='1' AND  A(14)='0' AND A(22)='0' AND A(11)='0' )then
          cVar2S19S61P011P014P017nsss(0) <='1';
          else
          cVar2S19S61P011P014P017nsss(0) <='0';
          end if;
        if(cVar1S20S61N018P061N059N063(0)='1' AND  A(15)='1' )then
          cVar2S20S61P009nsss(0) <='1';
          else
          cVar2S20S61P009nsss(0) <='0';
          end if;
        if(cVar1S0S62P000P018P061P028(0)='1' AND  A(24)='1' AND A(22)='0' )then
          cVar2S0S62P010P014nsss(0) <='1';
          else
          cVar2S0S62P010P014nsss(0) <='0';
          end if;
        if(cVar1S1S62P000P018P061P028(0)='1' AND  A(24)='0' AND B(23)='0' AND E(20)='1' )then
          cVar2S1S62N010P030P053nsss(0) <='1';
          else
          cVar2S1S62N010P030P053nsss(0) <='0';
          end if;
        if(cVar1S2S62P000P018P061N028(0)='1' AND  B(25)='1' AND D(11)='0' )then
          cVar2S2S62P026P054nsss(0) <='1';
          else
          cVar2S2S62P026P054nsss(0) <='0';
          end if;
        if(cVar1S3S62P000P018P061N028(0)='1' AND  B(25)='0' AND E(20)='0' AND D(20)='0' )then
          cVar2S3S62N026P053P051nsss(0) <='1';
          else
          cVar2S3S62N026P053P051nsss(0) <='0';
          end if;
        if(cVar1S4S62P000P018P061N028(0)='1' AND  B(25)='0' AND E(20)='1' AND A(14)='1' )then
          cVar2S4S62N026P053P011nsss(0) <='1';
          else
          cVar2S4S62N026P053P011nsss(0) <='0';
          end if;
        if(cVar1S5S62P000P018P061P059(0)='1' AND  E(16)='1' AND D(20)='0' )then
          cVar2S5S62P069P051nsss(0) <='1';
          else
          cVar2S5S62P069P051nsss(0) <='0';
          end if;
        if(cVar1S6S62P000P018P061N059(0)='1' AND  D(17)='1' AND E(10)='1' )then
          cVar2S6S62P063P060nsss(0) <='1';
          else
          cVar2S6S62P063P060nsss(0) <='0';
          end if;
        if(cVar1S7S62P000P018P061N059(0)='1' AND  D(17)='0' AND B(20)='0' AND A(15)='1' )then
          cVar2S7S62N063P036P009nsss(0) <='1';
          else
          cVar2S7S62N063P036P009nsss(0) <='0';
          end if;
        if(cVar1S8S62P000P018P043P024(0)='1' AND  E(22)='0' AND E(18)='1' )then
          cVar2S8S62P045P061nsss(0) <='1';
          else
          cVar2S8S62P045P061nsss(0) <='0';
          end if;
        if(cVar1S9S62P000P018P043P024(0)='1' AND  E(22)='0' AND E(18)='0' AND A(25)='0' )then
          cVar2S9S62P045N061P008nsss(0) <='1';
          else
          cVar2S9S62P045N061P008nsss(0) <='0';
          end if;
        if(cVar1S10S62P000P018P043P024(0)='1' AND  E(22)='1' AND D( 8)='0' AND B(20)='1' )then
          cVar2S10S62P045P066P036nsss(0) <='1';
          else
          cVar2S10S62P045P066P036nsss(0) <='0';
          end if;
        if(cVar1S11S62P000P018P043P045(0)='1' AND  A(12)='1' )then
          cVar2S11S62P015nsss(0) <='1';
          else
          cVar2S11S62P015nsss(0) <='0';
          end if;
        if(cVar1S12S62P000P030P027P056(0)='1' AND  E(19)='0' AND B(13)='0' )then
          cVar2S12S62P057P031nsss(0) <='1';
          else
          cVar2S12S62P057P031nsss(0) <='0';
          end if;
        if(cVar1S0S63P000P018P028P010(0)='1' AND  A(22)='0' )then
          cVar2S0S63P014nsss(0) <='1';
          else
          cVar2S0S63P014nsss(0) <='0';
          end if;
        if(cVar1S1S63P000P018P028N010(0)='1' AND  B(23)='0' AND A(26)='0' AND A(10)='1' )then
          cVar2S1S63P030P006P019nsss(0) <='1';
          else
          cVar2S1S63P030P006P019nsss(0) <='0';
          end if;
        if(cVar1S2S63P000P018N028P030(0)='1' AND  A(23)='1' AND A(22)='0' )then
          cVar2S2S63P012P014nsss(0) <='1';
          else
          cVar2S2S63P012P014nsss(0) <='0';
          end if;
        if(cVar1S3S63P000P018N028P030(0)='1' AND  A(23)='1' AND A(22)='1' AND A(12)='0' )then
          cVar2S3S63P012P014P015nsss(0) <='1';
          else
          cVar2S3S63P012P014P015nsss(0) <='0';
          end if;
        if(cVar1S4S63P000P018N028P030(0)='1' AND  A(23)='0' AND D(10)='1' )then
          cVar2S4S63N012P058nsss(0) <='1';
          else
          cVar2S4S63N012P058nsss(0) <='0';
          end if;
        if(cVar1S5S63P000P018N028P030(0)='1' AND  A(23)='0' AND D(10)='0' AND A(21)='1' )then
          cVar2S5S63N012N058P016nsss(0) <='1';
          else
          cVar2S5S63N012N058P016nsss(0) <='0';
          end if;
        if(cVar1S6S63P000P018N028N030(0)='1' AND  E(19)='0' AND D(11)='0' AND B(25)='1' )then
          cVar2S6S63P057P054P026nsss(0) <='1';
          else
          cVar2S6S63P057P054P026nsss(0) <='0';
          end if;
        if(cVar1S7S63P000P018N028N030(0)='1' AND  E(19)='0' AND D(11)='1' AND A(13)='1' )then
          cVar2S7S63P057P054P013nsss(0) <='1';
          else
          cVar2S7S63P057P054P013nsss(0) <='0';
          end if;
        if(cVar1S8S63P000P018N028N030(0)='1' AND  E(19)='1' AND D( 9)='0' AND D(11)='1' )then
          cVar2S8S63P057P062P054nsss(0) <='1';
          else
          cVar2S8S63P057P062P054nsss(0) <='0';
          end if;
        if(cVar1S9S63P000P018P036P004(0)='1' AND  D( 9)='1' AND E(16)='1' )then
          cVar2S9S63P062P069nsss(0) <='1';
          else
          cVar2S9S63P062P069nsss(0) <='0';
          end if;
        if(cVar1S10S63P000P018P036P004(0)='1' AND  D( 9)='1' AND E(16)='0' AND D( 8)='1' )then
          cVar2S10S63P062N069P066nsss(0) <='1';
          else
          cVar2S10S63P062N069P066nsss(0) <='0';
          end if;
        if(cVar1S11S63P000P018P036P004(0)='1' AND  D( 9)='0' AND A(19)='0' )then
          cVar2S11S63N062P001nsss(0) <='1';
          else
          cVar2S11S63N062P001nsss(0) <='0';
          end if;
        if(cVar1S12S63P000P018P036P004(0)='1' AND  A(21)='0' AND A(22)='1' )then
          cVar2S12S63P016P014nsss(0) <='1';
          else
          cVar2S12S63P016P014nsss(0) <='0';
          end if;
        if(cVar1S13S63P000P018N036P057(0)='1' AND  B(23)='0' AND E(11)='0' AND E(18)='1' )then
          cVar2S13S63P030P056P061nsss(0) <='1';
          else
          cVar2S13S63P030P056P061nsss(0) <='0';
          end if;
        if(cVar1S14S63P000P018N036P057(0)='1' AND  B(23)='1' AND E(16)='1' )then
          cVar2S14S63P030P069nsss(0) <='1';
          else
          cVar2S14S63P030P069nsss(0) <='0';
          end if;
        if(cVar1S15S63P000P018N036P057(0)='1' AND  E( 8)='0' AND A(11)='0' AND D(19)='1' )then
          cVar2S15S63P068P017P055nsss(0) <='1';
          else
          cVar2S15S63P068P017P055nsss(0) <='0';
          end if;
        if(cVar1S16S63P000P018N036P057(0)='1' AND  E( 8)='0' AND A(11)='1' AND D(18)='1' )then
          cVar2S16S63P068P017P059nsss(0) <='1';
          else
          cVar2S16S63P068P017P059nsss(0) <='0';
          end if;
        if(cVar1S17S63P000P030P027P020(0)='1' AND  D(18)='0' AND E(19)='0' AND B(26)='1' )then
          cVar2S17S63P059P057P024nsss(0) <='1';
          else
          cVar2S17S63P059P057P024nsss(0) <='0';
          end if;
        if(cVar1S0S64P018P061P059P028(0)='1' AND  A(24)='1' AND D(16)='0' )then
          cVar2S0S64P010P067nsss(0) <='1';
          else
          cVar2S0S64P010P067nsss(0) <='0';
          end if;
        if(cVar1S1S64P018P061P059P028(0)='1' AND  A(24)='0' AND A(26)='0' AND E(20)='1' )then
          cVar2S1S64N010P006P053nsss(0) <='1';
          else
          cVar2S1S64N010P006P053nsss(0) <='0';
          end if;
        if(cVar1S2S64P018P061P059N028(0)='1' AND  E(23)='1' AND B(28)='1' )then
          cVar2S2S64P041P020nsss(0) <='1';
          else
          cVar2S2S64P041P020nsss(0) <='0';
          end if;
        if(cVar1S3S64P018P061P059N028(0)='1' AND  E(23)='1' AND B(28)='0' AND B(18)='1' )then
          cVar2S3S64P041N020P021nsss(0) <='1';
          else
          cVar2S3S64P041N020P021nsss(0) <='0';
          end if;
        if(cVar1S4S64P018P061P059N028(0)='1' AND  E(23)='0' AND B(28)='0' AND A(28)='0' )then
          cVar2S4S64N041P020P002nsss(0) <='1';
          else
          cVar2S4S64N041P020P002nsss(0) <='0';
          end if;
        if(cVar1S5S64P018P061P059N028(0)='1' AND  E(23)='0' AND B(28)='1' AND E(15)='1' )then
          cVar2S5S64N041P020P040nsss(0) <='1';
          else
          cVar2S5S64N041P020P040nsss(0) <='0';
          end if;
        if(cVar1S6S64P018P061P059P012(0)='1' AND  B(20)='0' AND A(24)='0' )then
          cVar2S6S64P036P010nsss(0) <='1';
          else
          cVar2S6S64P036P010nsss(0) <='0';
          end if;
        if(cVar1S7S64P018P061P059P000(0)='1' AND  A(15)='0' AND A(23)='1' AND A(13)='0' )then
          cVar2S7S64P009P012P013nsss(0) <='1';
          else
          cVar2S7S64P009P012P013nsss(0) <='0';
          end if;
        if(cVar1S8S64P018P061P059P000(0)='1' AND  A(15)='0' AND A(23)='0' AND E( 9)='0' )then
          cVar2S8S64P009N012P064nsss(0) <='1';
          else
          cVar2S8S64P009N012P064nsss(0) <='0';
          end if;
        if(cVar1S9S64P018P061P059P000(0)='1' AND  A(15)='1' AND B(21)='1' )then
          cVar2S9S64P009P034nsss(0) <='1';
          else
          cVar2S9S64P009P034nsss(0) <='0';
          end if;
        if(cVar1S10S64P018P061N059P063(0)='1' AND  A(14)='0' AND A(22)='0' )then
          cVar2S10S64P011P014nsss(0) <='1';
          else
          cVar2S10S64P011P014nsss(0) <='0';
          end if;
        if(cVar1S11S64P018P061N059N063(0)='1' AND  B(20)='0' AND A(15)='1' )then
          cVar2S11S64P036P009nsss(0) <='1';
          else
          cVar2S11S64P036P009nsss(0) <='0';
          end if;
        if(cVar1S12S64P018P034P039P050(0)='1' AND  E( 9)='1' AND A(21)='0' )then
          cVar2S12S64P064P016nsss(0) <='1';
          else
          cVar2S12S64P064P016nsss(0) <='0';
          end if;
        if(cVar1S13S64P018P034P039P050(0)='1' AND  E( 9)='1' AND A(21)='1' AND A(11)='0' )then
          cVar2S13S64P064P016P017nsss(0) <='1';
          else
          cVar2S13S64P064P016P017nsss(0) <='0';
          end if;
        if(cVar1S14S64P018P034P039P050(0)='1' AND  E( 9)='0' AND D( 9)='0' AND A(26)='1' )then
          cVar2S14S64N064P062P006nsss(0) <='1';
          else
          cVar2S14S64N064P062P006nsss(0) <='0';
          end if;
        if(cVar1S15S64P018P034P039P050(0)='1' AND  E( 9)='0' AND D( 9)='1' AND A(13)='1' )then
          cVar2S15S64N064P062P013nsss(0) <='1';
          else
          cVar2S15S64N064P062P013nsss(0) <='0';
          end if;
        if(cVar1S16S64P018P034P039P050(0)='1' AND  E(13)='1' AND A(10)='0' )then
          cVar2S16S64P048P019nsss(0) <='1';
          else
          cVar2S16S64P048P019nsss(0) <='0';
          end if;
        if(cVar1S17S64P018P034P039P050(0)='1' AND  E(13)='0' AND B(14)='1' )then
          cVar2S17S64N048P029nsss(0) <='1';
          else
          cVar2S17S64N048P029nsss(0) <='0';
          end if;
        if(cVar1S18S64P018P034P039P050(0)='1' AND  E(13)='0' AND B(14)='0' AND A(15)='1' )then
          cVar2S18S64N048N029P009nsss(0) <='1';
          else
          cVar2S18S64N048N029P009nsss(0) <='0';
          end if;
        if(cVar1S20S64P018P034P047P069(0)='1' AND  D(19)='0' AND A(15)='1' AND A(13)='0' )then
          cVar2S20S64P055P009P013nsss(0) <='1';
          else
          cVar2S20S64P055P009P013nsss(0) <='0';
          end if;
        if(cVar1S21S64P018P034P047P069(0)='1' AND  D(19)='0' AND A(15)='0' AND B(10)='1' )then
          cVar2S21S64P055N009P037nsss(0) <='1';
          else
          cVar2S21S64P055N009P037nsss(0) <='0';
          end if;
        if(cVar1S22S64P018P034P047P069(0)='1' AND  E(17)='1' AND A(23)='0' AND B(20)='1' )then
          cVar2S22S64P065P012P036nsss(0) <='1';
          else
          cVar2S22S64P065P012P036nsss(0) <='0';
          end if;
        if(cVar1S0S65P018P034P050P039(0)='1' AND  E(17)='1' AND A(26)='0' AND A(21)='0' )then
          cVar2S0S65P065P006P016nsss(0) <='1';
          else
          cVar2S0S65P065P006P016nsss(0) <='0';
          end if;
        if(cVar1S1S65P018P034P050P039(0)='1' AND  E(17)='0' AND B(20)='0' AND D( 9)='0' )then
          cVar2S1S65N065P036P062nsss(0) <='1';
          else
          cVar2S1S65N065P036P062nsss(0) <='0';
          end if;
        if(cVar1S2S65P018P034P050P039(0)='1' AND  E(17)='0' AND B(20)='1' AND E( 9)='1' )then
          cVar2S2S65N065P036P064nsss(0) <='1';
          else
          cVar2S2S65N065P036P064nsss(0) <='0';
          end if;
        if(cVar1S3S65P018P034P050P039(0)='1' AND  A(21)='0' AND E(23)='1' )then
          cVar2S3S65P016P041nsss(0) <='1';
          else
          cVar2S3S65P016P041nsss(0) <='0';
          end if;
        if(cVar1S4S65P018P034P050P039(0)='1' AND  A(21)='0' AND E(23)='0' AND A(22)='1' )then
          cVar2S4S65P016N041P014nsss(0) <='1';
          else
          cVar2S4S65P016N041P014nsss(0) <='0';
          end if;
        if(cVar1S5S65P018P034P050P048(0)='1' AND  A(10)='0' )then
          cVar2S5S65P019nsss(0) <='1';
          else
          cVar2S5S65P019nsss(0) <='0';
          end if;
        if(cVar1S6S65P018P034P050N048(0)='1' AND  B(14)='1' )then
          cVar2S6S65P029nsss(0) <='1';
          else
          cVar2S6S65P029nsss(0) <='0';
          end if;
        if(cVar1S7S65P018P034P050N048(0)='1' AND  B(14)='0' AND A(17)='0' AND A(15)='1' )then
          cVar2S7S65N029P005P009nsss(0) <='1';
          else
          cVar2S7S65N029P005P009nsss(0) <='0';
          end if;
        if(cVar1S8S65P018P034P047P069(0)='1' AND  D(19)='0' AND E(10)='0' AND A(23)='1' )then
          cVar2S8S65P055P060P012nsss(0) <='1';
          else
          cVar2S8S65P055P060P012nsss(0) <='0';
          end if;
        if(cVar1S9S65P018P034P047P069(0)='1' AND  E(17)='1' AND A(23)='0' AND A(12)='1' )then
          cVar2S9S65P065P012P015nsss(0) <='1';
          else
          cVar2S9S65P065P012P015nsss(0) <='0';
          end if;
        if(cVar1S10S65N018P028P030P010(0)='1' AND  E(19)='1' )then
          cVar2S10S65P057nsss(0) <='1';
          else
          cVar2S10S65P057nsss(0) <='0';
          end if;
        if(cVar1S11S65N018P028P030P010(0)='1' AND  E(19)='0' AND E(12)='1' )then
          cVar2S11S65N057P052nsss(0) <='1';
          else
          cVar2S11S65N057P052nsss(0) <='0';
          end if;
        if(cVar1S12S65N018P028P030P010(0)='1' AND  E(19)='0' AND E(12)='0' AND D(20)='1' )then
          cVar2S12S65N057N052P051nsss(0) <='1';
          else
          cVar2S12S65N057N052P051nsss(0) <='0';
          end if;
        if(cVar1S13S65N018P028P030N010(0)='1' AND  A(26)='0' AND D(16)='0' )then
          cVar2S13S65P006P067nsss(0) <='1';
          else
          cVar2S13S65P006P067nsss(0) <='0';
          end if;
        if(cVar1S14S65N018N028P041P039(0)='1' AND  B(28)='1' )then
          cVar2S14S65P020nsss(0) <='1';
          else
          cVar2S14S65P020nsss(0) <='0';
          end if;
        if(cVar1S15S65N018N028P041P039(0)='1' AND  B(28)='0' AND A(23)='0' )then
          cVar2S15S65N020P012nsss(0) <='1';
          else
          cVar2S15S65N020P012nsss(0) <='0';
          end if;
        if(cVar1S16S65N018N028P041N039(0)='1' AND  B(20)='0' AND A(25)='0' AND A(13)='0' )then
          cVar2S16S65P036P008P013nsss(0) <='1';
          else
          cVar2S16S65P036P008P013nsss(0) <='0';
          end if;
        if(cVar1S17S65N018N028N041P039(0)='1' AND  B(28)='0' AND B(12)='0' AND A(21)='1' )then
          cVar2S17S65P020P033P016nsss(0) <='1';
          else
          cVar2S17S65P020P033P016nsss(0) <='0';
          end if;
        if(cVar1S18S65N018N028N041P039(0)='1' AND  B(28)='1' AND E(15)='1' )then
          cVar2S18S65P020P040nsss(0) <='1';
          else
          cVar2S18S65P020P040nsss(0) <='0';
          end if;
        if(cVar1S19S65N018N028N041P039(0)='1' AND  B(28)='1' AND E(15)='0' AND A(16)='1' )then
          cVar2S19S65P020N040P007nsss(0) <='1';
          else
          cVar2S19S65P020N040P007nsss(0) <='0';
          end if;
        if(cVar1S20S65N018N028N041P039(0)='1' AND  A(24)='0' AND A(23)='0' AND A(21)='0' )then
          cVar2S20S65P010P012P016nsss(0) <='1';
          else
          cVar2S20S65P010P012P016nsss(0) <='0';
          end if;
        if(cVar1S1S66P016P000P002N040(0)='1' AND  E(23)='1' )then
          cVar2S1S66P041nsss(0) <='1';
          else
          cVar2S1S66P041nsss(0) <='0';
          end if;
        if(cVar1S2S66P016P000P002N040(0)='1' AND  E(23)='0' AND B(22)='0' )then
          cVar2S2S66N041P032nsss(0) <='1';
          else
          cVar2S2S66N041P032nsss(0) <='0';
          end if;
        if(cVar1S3S66P016P000N002P034(0)='1' AND  B(22)='1' AND A(22)='1' )then
          cVar2S3S66P032P014nsss(0) <='1';
          else
          cVar2S3S66P032P014nsss(0) <='0';
          end if;
        if(cVar1S4S66P016P000N002P034(0)='1' AND  B(22)='1' AND A(22)='0' AND A(13)='1' )then
          cVar2S4S66P032N014P013nsss(0) <='1';
          else
          cVar2S4S66P032N014P013nsss(0) <='0';
          end if;
        if(cVar1S5S66P016P000N002P034(0)='1' AND  B(22)='0' AND A(22)='0' )then
          cVar2S5S66N032P014nsss(0) <='1';
          else
          cVar2S5S66N032P014nsss(0) <='0';
          end if;
        if(cVar1S6S66P016P000N002P034(0)='1' AND  A(22)='1' AND B(22)='0' )then
          cVar2S6S66P014P032nsss(0) <='1';
          else
          cVar2S6S66P014P032nsss(0) <='0';
          end if;
        if(cVar1S7S66P016P000P053P031(0)='1' AND  B(15)='0' AND B(21)='1' AND D( 8)='0' )then
          cVar2S7S66P027P034P066nsss(0) <='1';
          else
          cVar2S7S66P027P034P066nsss(0) <='0';
          end if;
        if(cVar1S8S66P016P039P022P041(0)='1' AND  D(22)='0' AND D(17)='1' AND E(17)='1' )then
          cVar2S8S66P043P063P065nsss(0) <='1';
          else
          cVar2S8S66P043P063P065nsss(0) <='0';
          end if;
        if(cVar1S9S66P016P039P022P041(0)='1' AND  E(16)='0' AND A(24)='0' AND A(12)='1' )then
          cVar2S9S66P069P010P015nsss(0) <='1';
          else
          cVar2S9S66P069P010P015nsss(0) <='0';
          end if;
        if(cVar1S10S66P016P039P022P019(0)='1' AND  A(14)='1' )then
          cVar2S10S66P011nsss(0) <='1';
          else
          cVar2S10S66P011nsss(0) <='0';
          end if;
        if(cVar1S12S66P016P039P007N005(0)='1' AND  E(16)='0' AND D(20)='1' )then
          cVar2S12S66P069P051nsss(0) <='1';
          else
          cVar2S12S66P069P051nsss(0) <='0';
          end if;
        if(cVar1S0S67P014P024P027P044(0)='1' AND  B(10)='1' AND D(23)='0' AND E(19)='0' )then
          cVar2S0S67P037P039P057nsss(0) <='1';
          else
          cVar2S0S67P037P039P057nsss(0) <='0';
          end if;
        if(cVar1S1S67P014P024P027P044(0)='1' AND  B(10)='0' AND E(16)='0' AND B(11)='0' )then
          cVar2S1S67N037P069P035nsss(0) <='1';
          else
          cVar2S1S67N037P069P035nsss(0) <='0';
          end if;
        if(cVar1S2S67P014P024P027P044(0)='1' AND  B(10)='0' AND E(16)='1' AND B(22)='1' )then
          cVar2S2S67N037P069P032nsss(0) <='1';
          else
          cVar2S2S67N037P069P032nsss(0) <='0';
          end if;
        if(cVar1S3S67P014P024P027P044(0)='1' AND  E(17)='0' AND A(11)='0' AND A(20)='1' )then
          cVar2S3S67P065P017P018nsss(0) <='1';
          else
          cVar2S3S67P065P017P018nsss(0) <='0';
          end if;
        if(cVar1S7S67N014P027P009N050(0)='1' AND  A(11)='0' )then
          cVar2S7S67P017nsss(0) <='1';
          else
          cVar2S7S67P017nsss(0) <='0';
          end if;
        if(cVar1S8S67N014P027N009P000(0)='1' AND  E(20)='0' AND A(14)='0' )then
          cVar2S8S67P053P011nsss(0) <='1';
          else
          cVar2S8S67P053P011nsss(0) <='0';
          end if;
        if(cVar1S9S67N014N027P050P024(0)='1' AND  D(21)='1' )then
          cVar2S9S67P047nsss(0) <='1';
          else
          cVar2S9S67P047nsss(0) <='0';
          end if;
        if(cVar1S10S67N014N027P050P024(0)='1' AND  D(21)='0' AND D(22)='1' )then
          cVar2S10S67N047P043nsss(0) <='1';
          else
          cVar2S10S67N047P043nsss(0) <='0';
          end if;
        if(cVar1S11S67N014N027P050N024(0)='1' AND  D(21)='0' AND E(13)='1' AND B(16)='1' )then
          cVar2S11S67P047P048P025nsss(0) <='1';
          else
          cVar2S11S67P047P048P025nsss(0) <='0';
          end if;
        if(cVar1S12S67N014N027P050N024(0)='1' AND  D(21)='1' AND B(25)='1' )then
          cVar2S12S67P047P026nsss(0) <='1';
          else
          cVar2S12S67P047P026nsss(0) <='0';
          end if;
        if(cVar1S13S67N014N027P050P032(0)='1' AND  A(25)='1' AND B(25)='1' )then
          cVar2S13S67P008P026nsss(0) <='1';
          else
          cVar2S13S67P008P026nsss(0) <='0';
          end if;
        if(cVar1S14S67N014N027P050P032(0)='1' AND  A(25)='1' AND B(25)='0' AND A(11)='0' )then
          cVar2S14S67P008N026P017nsss(0) <='1';
          else
          cVar2S14S67P008N026P017nsss(0) <='0';
          end if;
        if(cVar1S15S67N014N027P050P032(0)='1' AND  A(25)='0' AND A(24)='1' AND E(12)='1' )then
          cVar2S15S67N008P010P052nsss(0) <='1';
          else
          cVar2S15S67N008P010P052nsss(0) <='0';
          end if;
        if(cVar1S0S68P006P024P049P026(0)='1' AND  D(19)='1' AND E(17)='1' AND B(21)='0' )then
          cVar2S0S68P055P065P034nsss(0) <='1';
          else
          cVar2S0S68P055P065P034nsss(0) <='0';
          end if;
        if(cVar1S1S68P006P024P049P026(0)='1' AND  D(19)='1' AND E(17)='0' AND E(16)='1' )then
          cVar2S1S68P055N065P069nsss(0) <='1';
          else
          cVar2S1S68P055N065P069nsss(0) <='0';
          end if;
        if(cVar1S2S68P006P024P049P026(0)='1' AND  D(19)='0' AND E(19)='0' AND D(21)='0' )then
          cVar2S2S68N055P057P047nsss(0) <='1';
          else
          cVar2S2S68N055P057P047nsss(0) <='0';
          end if;
        if(cVar1S3S68P006P024P049P026(0)='1' AND  E(13)='1' )then
          cVar2S3S68P048nsss(0) <='1';
          else
          cVar2S3S68P048nsss(0) <='0';
          end if;
        if(cVar1S5S68P006P024P049N026(0)='1' AND  B(15)='1' )then
          cVar2S5S68P027nsss(0) <='1';
          else
          cVar2S5S68P027nsss(0) <='0';
          end if;
        if(cVar1S6S68P006P024P049N026(0)='1' AND  B(15)='0' AND D(13)='1' )then
          cVar2S6S68N027P046nsss(0) <='1';
          else
          cVar2S6S68N027P046nsss(0) <='0';
          end if;
        if(cVar1S8S68P006P024P010N047(0)='1' AND  A(29)='1' )then
          cVar2S8S68P000nsss(0) <='1';
          else
          cVar2S8S68P000nsss(0) <='0';
          end if;
        if(cVar1S9S68P006P024P010N047(0)='1' AND  A(29)='0' AND D(20)='0' AND A(27)='1' )then
          cVar2S9S68N000P051P004nsss(0) <='1';
          else
          cVar2S9S68N000P051P004nsss(0) <='0';
          end if;
        if(cVar1S10S68P006P024P010P019(0)='1' AND  B(20)='0' AND D( 8)='1' )then
          cVar2S10S68P036P066nsss(0) <='1';
          else
          cVar2S10S68P036P066nsss(0) <='0';
          end if;
        if(cVar1S11S68P006P024P002P011(0)='1' AND  D(21)='1' )then
          cVar2S11S68P047nsss(0) <='1';
          else
          cVar2S11S68P047nsss(0) <='0';
          end if;
        if(cVar1S12S68P006P024P002P011(0)='1' AND  D(21)='0' AND A(13)='0' AND A(12)='0' )then
          cVar2S12S68N047P013P015nsss(0) <='1';
          else
          cVar2S12S68N047P013P015nsss(0) <='0';
          end if;
        if(cVar1S13S68P006N024P065P034(0)='1' AND  A(17)='0' AND A(29)='0' AND A(28)='1' )then
          cVar2S13S68P005P000P002nsss(0) <='1';
          else
          cVar2S13S68P005P000P002nsss(0) <='0';
          end if;
        if(cVar1S14S68P006N024P065P034(0)='1' AND  A(17)='1' AND A(24)='1' )then
          cVar2S14S68P005P010nsss(0) <='1';
          else
          cVar2S14S68P005P010nsss(0) <='0';
          end if;
        if(cVar1S15S68P006N024P065P034(0)='1' AND  B(20)='0' AND A(14)='0' AND A(12)='1' )then
          cVar2S15S68P036P011P015nsss(0) <='1';
          else
          cVar2S15S68P036P011P015nsss(0) <='0';
          end if;
        if(cVar1S16S68P006N024P065P013(0)='1' AND  A(22)='0' AND D(16)='1' )then
          cVar2S16S68P014P067nsss(0) <='1';
          else
          cVar2S16S68P014P067nsss(0) <='0';
          end if;
        if(cVar1S0S69P055P026P010P057(0)='1' AND  A(23)='0' )then
          cVar2S0S69P012nsss(0) <='1';
          else
          cVar2S0S69P012nsss(0) <='0';
          end if;
        if(cVar1S1S69P055P026P010P057(0)='1' AND  A(23)='1' AND A(22)='0' )then
          cVar2S1S69P012P014nsss(0) <='1';
          else
          cVar2S1S69P012P014nsss(0) <='0';
          end if;
        if(cVar1S2S69P055P026P010N057(0)='1' AND  A(23)='1' )then
          cVar2S2S69P012nsss(0) <='1';
          else
          cVar2S2S69P012nsss(0) <='0';
          end if;
        if(cVar1S4S69P055P026N010N065(0)='1' AND  A(26)='0' AND E(16)='1' AND E(19)='1' )then
          cVar2S4S69P006P069P057nsss(0) <='1';
          else
          cVar2S4S69P006P069P057nsss(0) <='0';
          end if;
        if(cVar1S5S69P055P026N010N065(0)='1' AND  A(26)='0' AND E(16)='0' AND A(14)='1' )then
          cVar2S5S69P006N069P011nsss(0) <='1';
          else
          cVar2S5S69P006N069P011nsss(0) <='0';
          end if;
        if(cVar1S6S69N055P030P026P004(0)='1' AND  A(25)='1' )then
          cVar2S6S69P008nsss(0) <='1';
          else
          cVar2S6S69P008nsss(0) <='0';
          end if;
        if(cVar1S7S69N055P030P026P004(0)='1' AND  A(25)='0' AND E(11)='0' )then
          cVar2S7S69N008P056nsss(0) <='1';
          else
          cVar2S7S69N008P056nsss(0) <='0';
          end if;
        if(cVar1S8S69N055P030N026P057(0)='1' AND  B(26)='1' AND A(24)='0' )then
          cVar2S8S69P024P010nsss(0) <='1';
          else
          cVar2S8S69P024P010nsss(0) <='0';
          end if;
        if(cVar1S9S69N055P030N026P057(0)='1' AND  B(26)='0' AND D(21)='1' AND B(15)='1' )then
          cVar2S9S69N024P047P027nsss(0) <='1';
          else
          cVar2S9S69N024P047P027nsss(0) <='0';
          end if;
        if(cVar1S11S69N055P030P063N002(0)='1' AND  E(11)='1' AND A(23)='1' )then
          cVar2S11S69P056P012nsss(0) <='1';
          else
          cVar2S11S69P056P012nsss(0) <='0';
          end if;
        if(cVar1S12S69N055P030P063N002(0)='1' AND  E(11)='0' AND D(18)='1' AND A(23)='1' )then
          cVar2S12S69N056P059P012nsss(0) <='1';
          else
          cVar2S12S69N056P059P012nsss(0) <='0';
          end if;
        if(cVar1S13S69N055P030P063N002(0)='1' AND  E(11)='0' AND D(18)='0' AND B(11)='1' )then
          cVar2S13S69N056N059P035nsss(0) <='1';
          else
          cVar2S13S69N056N059P035nsss(0) <='0';
          end if;
        if(cVar1S14S69N055P030P063P014(0)='1' AND  A(20)='1' )then
          cVar2S14S69P018nsss(0) <='1';
          else
          cVar2S14S69P018nsss(0) <='0';
          end if;
        if(cVar1S0S70P050P027P048P025(0)='1' AND  D(13)='0' AND B(18)='1' AND E(15)='1' )then
          cVar2S0S70P046P021P040nsss(0) <='1';
          else
          cVar2S0S70P046P021P040nsss(0) <='0';
          end if;
        if(cVar1S1S70P050P027P048P025(0)='1' AND  D(13)='0' AND B(18)='0' AND E(15)='0' )then
          cVar2S1S70P046N021P040nsss(0) <='1';
          else
          cVar2S1S70P046N021P040nsss(0) <='0';
          end if;
        if(cVar1S2S70P050P027P048P025(0)='1' AND  D(13)='1' AND A(20)='1' AND A(10)='0' )then
          cVar2S2S70P046P018P019nsss(0) <='1';
          else
          cVar2S2S70P046P018P019nsss(0) <='0';
          end if;
        if(cVar1S3S70P050P027P048P025(0)='1' AND  E(22)='1' )then
          cVar2S3S70P045nsss(0) <='1';
          else
          cVar2S3S70P045nsss(0) <='0';
          end if;
        if(cVar1S4S70P050P027P048P025(0)='1' AND  E(22)='0' AND B(26)='1' )then
          cVar2S4S70N045P024nsss(0) <='1';
          else
          cVar2S4S70N045P024nsss(0) <='0';
          end if;
        if(cVar1S5S70P050P027P048P025(0)='1' AND  E(22)='0' AND B(26)='0' AND A(16)='1' )then
          cVar2S5S70N045N024P007nsss(0) <='1';
          else
          cVar2S5S70N045N024P007nsss(0) <='0';
          end if;
        if(cVar1S7S70P050P027P048N025(0)='1' AND  D(21)='1' )then
          cVar2S7S70P047nsss(0) <='1';
          else
          cVar2S7S70P047nsss(0) <='0';
          end if;
        if(cVar1S8S70P050P027P048N025(0)='1' AND  D(21)='0' AND A(23)='1' AND B(20)='0' )then
          cVar2S8S70N047P012P036nsss(0) <='1';
          else
          cVar2S8S70N047P012P036nsss(0) <='0';
          end if;
        if(cVar1S9S70P050P027P048N025(0)='1' AND  D(21)='0' AND A(23)='0' AND E(16)='1' )then
          cVar2S9S70N047N012P069nsss(0) <='1';
          else
          cVar2S9S70N047N012P069nsss(0) <='0';
          end if;
        if(cVar1S10S70P050P027P000P035(0)='1' AND  B(22)='0' AND A(18)='1' )then
          cVar2S10S70P032P003nsss(0) <='1';
          else
          cVar2S10S70P032P003nsss(0) <='0';
          end if;
        if(cVar1S11S70P050P027P000P035(0)='1' AND  B(22)='0' AND A(18)='0' AND D(20)='1' )then
          cVar2S11S70P032N003P051nsss(0) <='1';
          else
          cVar2S11S70P032N003P051nsss(0) <='0';
          end if;
        if(cVar1S13S70P050P043P027N009(0)='1' AND  E(12)='0' )then
          cVar2S13S70P052nsss(0) <='1';
          else
          cVar2S13S70P052nsss(0) <='0';
          end if;
        if(cVar1S14S70P050P043N027P020(0)='1' AND  B(13)='1' )then
          cVar2S14S70P031nsss(0) <='1';
          else
          cVar2S14S70P031nsss(0) <='0';
          end if;
        if(cVar1S15S70P050P043N027P020(0)='1' AND  B(13)='0' AND E(12)='1' AND A(24)='1' )then
          cVar2S15S70N031P052P010nsss(0) <='1';
          else
          cVar2S15S70N031P052P010nsss(0) <='0';
          end if;
        if(cVar1S2S71P021N040P048N039(0)='1' AND  E(10)='0' AND E( 9)='1' )then
          cVar2S2S71P060P064nsss(0) <='1';
          else
          cVar2S2S71P060P064nsss(0) <='0';
          end if;
        if(cVar1S3S71N021P038P040P057(0)='1' AND  B(23)='1' AND A(26)='0' )then
          cVar2S3S71P030P006nsss(0) <='1';
          else
          cVar2S3S71P030P006nsss(0) <='0';
          end if;
        if(cVar1S4S71N021P038P040P057(0)='1' AND  B(23)='0' AND E(23)='0' AND B(13)='1' )then
          cVar2S4S71N030P041P031nsss(0) <='1';
          else
          cVar2S4S71N030P041P031nsss(0) <='0';
          end if;
        if(cVar1S5S71N021P038P040N057(0)='1' AND  B(23)='0' AND A(21)='1' AND A(28)='0' )then
          cVar2S5S71P030P016P002nsss(0) <='1';
          else
          cVar2S5S71P030P016P002nsss(0) <='0';
          end if;
        if(cVar1S6S71N021P038P040N057(0)='1' AND  B(23)='0' AND A(21)='0' AND B(22)='1' )then
          cVar2S6S71P030N016P032nsss(0) <='1';
          else
          cVar2S6S71P030N016P032nsss(0) <='0';
          end if;
        if(cVar1S7S71N021P038P040N057(0)='1' AND  B(23)='1' AND D(19)='0' AND D(11)='1' )then
          cVar2S7S71P030P055P054nsss(0) <='1';
          else
          cVar2S7S71P030P055P054nsss(0) <='0';
          end if;
        if(cVar1S8S71N021P038P040P059(0)='1' AND  A(28)='1' )then
          cVar2S8S71P002nsss(0) <='1';
          else
          cVar2S8S71P002nsss(0) <='0';
          end if;
        if(cVar1S9S71N021P038P040P059(0)='1' AND  A(28)='0' AND A(20)='1' AND A(12)='0' )then
          cVar2S9S71N002P018P015nsss(0) <='1';
          else
          cVar2S9S71N002P018P015nsss(0) <='0';
          end if;
        if(cVar1S10S71N021P038P040P059(0)='1' AND  A(28)='0' AND A(20)='0' AND B(10)='1' )then
          cVar2S10S71N002N018P037nsss(0) <='1';
          else
          cVar2S10S71N002N018P037nsss(0) <='0';
          end if;
        if(cVar1S12S71N021P038P040N015(0)='1' AND  A(20)='0' )then
          cVar2S12S71P018nsss(0) <='1';
          else
          cVar2S12S71P018nsss(0) <='0';
          end if;
        if(cVar1S1S72P016P021N038P011(0)='1' AND  A(10)='1' AND A(13)='0' AND A(11)='0' )then
          cVar2S1S72P019P013P017nsss(0) <='1';
          else
          cVar2S1S72P019P013P017nsss(0) <='0';
          end if;
        if(cVar1S2S72P016P021N038P011(0)='1' AND  A(10)='0' AND A(24)='0' AND E( 8)='0' )then
          cVar2S2S72N019P010P068nsss(0) <='1';
          else
          cVar2S2S72N019P010P068nsss(0) <='0';
          end if;
        if(cVar1S3S72P016N021P040P038(0)='1' AND  E(14)='1' AND B(17)='1' )then
          cVar2S3S72P044P023nsss(0) <='1';
          else
          cVar2S3S72P044P023nsss(0) <='0';
          end if;
        if(cVar1S4S72P016N021P040P038(0)='1' AND  E(14)='1' AND B(17)='0' AND A(13)='0' )then
          cVar2S4S72P044N023P013nsss(0) <='1';
          else
          cVar2S4S72P044N023P013nsss(0) <='0';
          end if;
        if(cVar1S5S72P016N021P040P038(0)='1' AND  E(14)='0' AND D(14)='0' AND A(17)='0' )then
          cVar2S5S72N044P042P005nsss(0) <='1';
          else
          cVar2S5S72N044P042P005nsss(0) <='0';
          end if;
        if(cVar1S6S72P016N021P040P038(0)='1' AND  A(24)='1' )then
          cVar2S6S72P010nsss(0) <='1';
          else
          cVar2S6S72P010nsss(0) <='0';
          end if;
        if(cVar1S8S72P016N021P040N002(0)='1' AND  E(17)='0' AND E(16)='1' )then
          cVar2S8S72P065P069nsss(0) <='1';
          else
          cVar2S8S72P065P069nsss(0) <='0';
          end if;
        if(cVar1S9S72P016P039P041P022(0)='1' AND  D(22)='0' AND B(10)='1' AND A(26)='0' )then
          cVar2S9S72P043P037P006nsss(0) <='1';
          else
          cVar2S9S72P043P037P006nsss(0) <='0';
          end if;
        if(cVar1S10S72P016P039P041P022(0)='1' AND  D(22)='1' AND E(17)='0' AND A(10)='0' )then
          cVar2S10S72P043P065P019nsss(0) <='1';
          else
          cVar2S10S72P043P065P019nsss(0) <='0';
          end if;
        if(cVar1S11S72P016P039P041P022(0)='1' AND  A(10)='1' AND A(14)='1' )then
          cVar2S11S72P019P011nsss(0) <='1';
          else
          cVar2S11S72P019P011nsss(0) <='0';
          end if;
        if(cVar1S12S72P016P039P041P069(0)='1' AND  A(24)='0' AND A(12)='1' )then
          cVar2S12S72P010P015nsss(0) <='1';
          else
          cVar2S12S72P010P015nsss(0) <='0';
          end if;
        if(cVar1S14S72P016P039P054N005(0)='1' AND  E(18)='1' )then
          cVar2S14S72P061nsss(0) <='1';
          else
          cVar2S14S72P061nsss(0) <='0';
          end if;
        if(cVar1S1S73P021N040P048P056(0)='1' AND  A(14)='0' AND B(28)='0' )then
          cVar2S1S73P011P020nsss(0) <='1';
          else
          cVar2S1S73P011P020nsss(0) <='0';
          end if;
        if(cVar1S2S73P021N040P048P056(0)='1' AND  A(14)='1' AND A(13)='0' AND A(21)='1' )then
          cVar2S2S73P011P013P016nsss(0) <='1';
          else
          cVar2S2S73P011P013P016nsss(0) <='0';
          end if;
        if(cVar1S3S73N021P038P040P057(0)='1' AND  E(23)='0' AND B(23)='1' AND A(22)='0' )then
          cVar2S3S73P041P030P014nsss(0) <='1';
          else
          cVar2S3S73P041P030P014nsss(0) <='0';
          end if;
        if(cVar1S4S73N021P038P040P057(0)='1' AND  E(23)='0' AND B(23)='0' AND B(13)='1' )then
          cVar2S4S73P041N030P031nsss(0) <='1';
          else
          cVar2S4S73P041N030P031nsss(0) <='0';
          end if;
        if(cVar1S5S73N021P038P040N057(0)='1' AND  B(23)='0' AND D(20)='1' AND B(24)='1' )then
          cVar2S5S73P030P051P028nsss(0) <='1';
          else
          cVar2S5S73P030P051P028nsss(0) <='0';
          end if;
        if(cVar1S6S73N021P038P040N057(0)='1' AND  B(23)='1' AND D(19)='0' AND D(11)='1' )then
          cVar2S6S73P030P055P054nsss(0) <='1';
          else
          cVar2S6S73P030P055P054nsss(0) <='0';
          end if;
        if(cVar1S7S73N021P038P040P059(0)='1' AND  A(28)='1' )then
          cVar2S7S73P002nsss(0) <='1';
          else
          cVar2S7S73P002nsss(0) <='0';
          end if;
        if(cVar1S8S73N021P038P040P059(0)='1' AND  A(28)='0' AND A(20)='1' AND A(23)='1' )then
          cVar2S8S73N002P018P012nsss(0) <='1';
          else
          cVar2S8S73N002P018P012nsss(0) <='0';
          end if;
        if(cVar1S9S73N021P038P040P059(0)='1' AND  A(28)='0' AND A(20)='0' AND B(10)='1' )then
          cVar2S9S73N002N018P037nsss(0) <='1';
          else
          cVar2S9S73N002N018P037nsss(0) <='0';
          end if;
        if(cVar1S11S73N021P038N020P063(0)='1' AND  A(23)='1' AND A(21)='0' )then
          cVar2S11S73P012P016nsss(0) <='1';
          else
          cVar2S11S73P012P016nsss(0) <='0';
          end if;
        if(cVar1S12S73N021P038N020P063(0)='1' AND  A(23)='0' AND A(20)='1' AND A(10)='1' )then
          cVar2S12S73N012P018P019nsss(0) <='1';
          else
          cVar2S12S73N012P018P019nsss(0) <='0';
          end if;
        if(cVar1S1S74P014P027P002N009(0)='1' AND  A(24)='0' AND A(25)='1' )then
          cVar2S1S74P010P008nsss(0) <='1';
          else
          cVar2S1S74P010P008nsss(0) <='0';
          end if;
        if(cVar1S2S74P014P027P002N009(0)='1' AND  A(24)='0' AND A(25)='0' AND A(23)='1' )then
          cVar2S2S74P010N008P012nsss(0) <='1';
          else
          cVar2S2S74P010N008P012nsss(0) <='0';
          end if;
        if(cVar1S3S74P014N027P010P028(0)='1' AND  D( 8)='0' )then
          cVar2S3S74P066nsss(0) <='1';
          else
          cVar2S3S74P066nsss(0) <='0';
          end if;
        if(cVar1S4S74P014N027P010P028(0)='1' AND  D( 8)='1' AND B(10)='1' )then
          cVar2S4S74P066P037nsss(0) <='1';
          else
          cVar2S4S74P066P037nsss(0) <='0';
          end if;
        if(cVar1S5S74P014N027P010N028(0)='1' AND  A(13)='1' AND D(23)='0' AND E(20)='0' )then
          cVar2S5S74P013P039P053nsss(0) <='1';
          else
          cVar2S5S74P013P039P053nsss(0) <='0';
          end if;
        if(cVar1S6S74P014N027P010N028(0)='1' AND  A(13)='0' AND B(22)='0' AND B(13)='1' )then
          cVar2S6S74N013P032P031nsss(0) <='1';
          else
          cVar2S6S74N013P032P031nsss(0) <='0';
          end if;
        if(cVar1S7S74P014N027N010P024(0)='1' AND  D(21)='1' )then
          cVar2S7S74P047nsss(0) <='1';
          else
          cVar2S7S74P047nsss(0) <='0';
          end if;
        if(cVar1S8S74P014N027N010P024(0)='1' AND  D(21)='0' AND D(11)='0' )then
          cVar2S8S74N047P054nsss(0) <='1';
          else
          cVar2S8S74N047P054nsss(0) <='0';
          end if;
        if(cVar1S9S74P014N027N010N024(0)='1' AND  D(21)='0' AND E(13)='0' AND B(16)='0' )then
          cVar2S9S74P047P048P025nsss(0) <='1';
          else
          cVar2S9S74P047P048P025nsss(0) <='0';
          end if;
        if(cVar1S10S74P014N027N010N024(0)='1' AND  D(21)='0' AND E(13)='1' AND B(16)='1' )then
          cVar2S10S74P047P048P025nsss(0) <='1';
          else
          cVar2S10S74P047P048P025nsss(0) <='0';
          end if;
        if(cVar1S11S74P014N027N010N024(0)='1' AND  D(21)='1' AND B(25)='1' )then
          cVar2S11S74P047P026nsss(0) <='1';
          else
          cVar2S11S74P047P026nsss(0) <='0';
          end if;
        if(cVar1S12S74P014N027N010N024(0)='1' AND  D(21)='1' AND B(25)='0' AND A(14)='1' )then
          cVar2S12S74P047N026P011nsss(0) <='1';
          else
          cVar2S12S74P047N026P011nsss(0) <='0';
          end if;
        if(cVar1S13S74P014P024P044P037(0)='1' AND  B(23)='0' AND E(13)='0' )then
          cVar2S13S74P030P048nsss(0) <='1';
          else
          cVar2S13S74P030P048nsss(0) <='0';
          end if;
        if(cVar1S14S74P014P024P044N037(0)='1' AND  E(13)='1' AND D( 9)='1' )then
          cVar2S14S74P048P062nsss(0) <='1';
          else
          cVar2S14S74P048P062nsss(0) <='0';
          end if;
        if(cVar1S15S74P014P024P044N037(0)='1' AND  E(13)='1' AND D( 9)='0' AND A(11)='0' )then
          cVar2S15S74P048N062P017nsss(0) <='1';
          else
          cVar2S15S74P048N062P017nsss(0) <='0';
          end if;
        if(cVar1S16S74P014P024P044N037(0)='1' AND  E(13)='0' AND B(15)='0' AND B(18)='1' )then
          cVar2S16S74N048P027P021nsss(0) <='1';
          else
          cVar2S16S74N048P027P021nsss(0) <='0';
          end if;
        if(cVar1S17S74P014P024P044P065(0)='1' AND  A(20)='1' AND A(11)='0' )then
          cVar2S17S74P018P017nsss(0) <='1';
          else
          cVar2S17S74P018P017nsss(0) <='0';
          end if;
        if(cVar1S19S74P014P024P031N045(0)='1' AND  A(23)='0' AND A(18)='0' AND E( 9)='1' )then
          cVar2S19S74P012P003P064nsss(0) <='1';
          else
          cVar2S19S74P012P003P064nsss(0) <='0';
          end if;
        if(cVar1S20S74P014P024P031N045(0)='1' AND  A(23)='1' AND A(29)='1' )then
          cVar2S20S74P012P000nsss(0) <='1';
          else
          cVar2S20S74P012P000nsss(0) <='0';
          end if;
        if(cVar1S0S75P010P024P028P003(0)='1' AND  B(21)='0' )then
          cVar2S0S75P034nsss(0) <='1';
          else
          cVar2S0S75P034nsss(0) <='0';
          end if;
        if(cVar1S1S75P010P024N028P045(0)='1' AND  B(13)='1' AND A(22)='0' )then
          cVar2S1S75P031P014nsss(0) <='1';
          else
          cVar2S1S75P031P014nsss(0) <='0';
          end if;
        if(cVar1S2S75P010P024N028P045(0)='1' AND  B(13)='0' AND B(14)='1' )then
          cVar2S2S75N031P029nsss(0) <='1';
          else
          cVar2S2S75N031P029nsss(0) <='0';
          end if;
        if(cVar1S3S75P010P024N028P045(0)='1' AND  B(13)='0' AND B(14)='0' AND D(10)='1' )then
          cVar2S3S75N031N029P058nsss(0) <='1';
          else
          cVar2S3S75N031N029P058nsss(0) <='0';
          end if;
        if(cVar1S4S75P010P024N028P045(0)='1' AND  A(20)='1' )then
          cVar2S4S75P018nsss(0) <='1';
          else
          cVar2S4S75P018nsss(0) <='0';
          end if;
        if(cVar1S5S75P010P024P064P019(0)='1' AND  B(20)='0' AND B(21)='1' )then
          cVar2S5S75P036P034nsss(0) <='1';
          else
          cVar2S5S75P036P034nsss(0) <='0';
          end if;
        if(cVar1S6S75P010P024P064P019(0)='1' AND  B(20)='0' AND B(21)='0' AND A(11)='0' )then
          cVar2S6S75P036N034P017nsss(0) <='1';
          else
          cVar2S6S75P036N034P017nsss(0) <='0';
          end if;
        if(cVar1S7S75N010P014P024P056(0)='1' AND  E(10)='1' AND B(21)='1' )then
          cVar2S7S75P060P034nsss(0) <='1';
          else
          cVar2S7S75P060P034nsss(0) <='0';
          end if;
        if(cVar1S8S75N010P014P024P056(0)='1' AND  E(10)='1' AND B(21)='0' AND B(20)='0' )then
          cVar2S8S75P060N034P036nsss(0) <='1';
          else
          cVar2S8S75P060N034P036nsss(0) <='0';
          end if;
        if(cVar1S9S75N010P014P024P056(0)='1' AND  E(10)='0' AND B(13)='0' AND D(10)='0' )then
          cVar2S9S75N060P031P058nsss(0) <='1';
          else
          cVar2S9S75N060P031P058nsss(0) <='0';
          end if;
        if(cVar1S10S75N010P014P024P056(0)='1' AND  E(10)='0' AND B(13)='1' AND D(16)='1' )then
          cVar2S10S75N060P031P067nsss(0) <='1';
          else
          cVar2S10S75N060P031P067nsss(0) <='0';
          end if;
        if(cVar1S11S75N010P014P024P056(0)='1' AND  A(13)='1' AND B(13)='1' )then
          cVar2S11S75P013P031nsss(0) <='1';
          else
          cVar2S11S75P013P031nsss(0) <='0';
          end if;
        if(cVar1S12S75N010P014P024P056(0)='1' AND  A(13)='0' AND A(23)='1' AND A(10)='1' )then
          cVar2S12S75N013P012P019nsss(0) <='1';
          else
          cVar2S12S75N013P012P019nsss(0) <='0';
          end if;
        if(cVar1S13S75N010P014P024P051(0)='1' AND  E( 8)='0' AND B(25)='0' AND D(16)='0' )then
          cVar2S13S75P068P026P067nsss(0) <='1';
          else
          cVar2S13S75P068P026P067nsss(0) <='0';
          end if;
        if(cVar1S15S75N010N014P027N050(0)='1' AND  D(13)='1' )then
          cVar2S15S75P046nsss(0) <='1';
          else
          cVar2S15S75P046nsss(0) <='0';
          end if;
        if(cVar1S16S75N010N014P027N050(0)='1' AND  D(13)='0' AND E(21)='1' )then
          cVar2S16S75N046P049nsss(0) <='1';
          else
          cVar2S16S75N046P049nsss(0) <='0';
          end if;
        if(cVar1S17S75N010N014P027N050(0)='1' AND  D(13)='0' AND E(21)='0' AND E(16)='0' )then
          cVar2S17S75N046N049P069nsss(0) <='1';
          else
          cVar2S17S75N046N049P069nsss(0) <='0';
          end if;
        if(cVar1S18S75N010N014N027P024(0)='1' AND  D(21)='1' )then
          cVar2S18S75P047nsss(0) <='1';
          else
          cVar2S18S75P047nsss(0) <='0';
          end if;
        if(cVar1S19S75N010N014N027P024(0)='1' AND  D(21)='0' AND D(11)='0' AND D(22)='1' )then
          cVar2S19S75N047P054P043nsss(0) <='1';
          else
          cVar2S19S75N047P054P043nsss(0) <='0';
          end if;
        if(cVar1S20S75N010N014N027N024(0)='1' AND  D(21)='0' AND E(14)='1' AND B(17)='1' )then
          cVar2S20S75P047P044P023nsss(0) <='1';
          else
          cVar2S20S75P047P044P023nsss(0) <='0';
          end if;
        if(cVar1S21S75N010N014N027N024(0)='1' AND  D(21)='0' AND E(14)='0' AND E(23)='1' )then
          cVar2S21S75P047N044P041nsss(0) <='1';
          else
          cVar2S21S75P047N044P041nsss(0) <='0';
          end if;
        if(cVar1S22S75N010N014N027N024(0)='1' AND  D(21)='1' AND B(25)='1' )then
          cVar2S22S75P047P026nsss(0) <='1';
          else
          cVar2S22S75P047P026nsss(0) <='0';
          end if;
        if(cVar1S0S76P014P010P032P021(0)='1' AND  B(24)='1' )then
          cVar2S0S76P028nsss(0) <='1';
          else
          cVar2S0S76P028nsss(0) <='0';
          end if;
        if(cVar1S1S76P014P010P032P021(0)='1' AND  B(24)='0' AND B(26)='0' )then
          cVar2S1S76N028P024nsss(0) <='1';
          else
          cVar2S1S76N028P024nsss(0) <='0';
          end if;
        if(cVar1S2S76P014P010P032P017(0)='1' AND  A(13)='1' )then
          cVar2S2S76P013nsss(0) <='1';
          else
          cVar2S2S76P013nsss(0) <='0';
          end if;
        if(cVar1S4S76P014N010P027N050(0)='1' AND  D(13)='1' )then
          cVar2S4S76P046nsss(0) <='1';
          else
          cVar2S4S76P046nsss(0) <='0';
          end if;
        if(cVar1S5S76P014N010P027N050(0)='1' AND  D(13)='0' AND E(21)='1' )then
          cVar2S5S76N046P049nsss(0) <='1';
          else
          cVar2S5S76N046P049nsss(0) <='0';
          end if;
        if(cVar1S6S76P014N010N027P050(0)='1' AND  E(12)='0' AND B(26)='1' )then
          cVar2S6S76P052P024nsss(0) <='1';
          else
          cVar2S6S76P052P024nsss(0) <='0';
          end if;
        if(cVar1S7S76P014N010N027P050(0)='1' AND  E(12)='0' AND B(26)='0' AND D(21)='0' )then
          cVar2S7S76P052N024P047nsss(0) <='1';
          else
          cVar2S7S76P052N024P047nsss(0) <='0';
          end if;
        if(cVar1S8S76P014N010N027P050(0)='1' AND  E(12)='1' AND D( 9)='1' )then
          cVar2S8S76P052P062nsss(0) <='1';
          else
          cVar2S8S76P052P062nsss(0) <='0';
          end if;
        if(cVar1S9S76P014N010N027P050(0)='1' AND  E(12)='1' AND D( 9)='0' AND E( 8)='1' )then
          cVar2S9S76P052N062P068nsss(0) <='1';
          else
          cVar2S9S76P052N062P068nsss(0) <='0';
          end if;
        if(cVar1S10S76P014N010N027P050(0)='1' AND  A(27)='0' AND A(25)='1' AND B(25)='1' )then
          cVar2S10S76P004P008P026nsss(0) <='1';
          else
          cVar2S10S76P004P008P026nsss(0) <='0';
          end if;
        if(cVar1S11S76P014N010N027P050(0)='1' AND  A(27)='0' AND A(25)='0' AND D(10)='1' )then
          cVar2S11S76P004N008P058nsss(0) <='1';
          else
          cVar2S11S76P004N008P058nsss(0) <='0';
          end if;
        if(cVar1S12S76P014P024P044P027(0)='1' AND  D(22)='0' AND B(27)='0' AND D(16)='1' )then
          cVar2S12S76P043P022P067nsss(0) <='1';
          else
          cVar2S12S76P043P022P067nsss(0) <='0';
          end if;
        if(cVar1S13S76P014P024P044P027(0)='1' AND  D(22)='1' AND B(20)='0' AND D( 8)='0' )then
          cVar2S13S76P043P036P066nsss(0) <='1';
          else
          cVar2S13S76P043P036P066nsss(0) <='0';
          end if;
        if(cVar1S14S76P014P024P044P027(0)='1' AND  B(20)='1' )then
          cVar2S14S76P036nsss(0) <='1';
          else
          cVar2S14S76P036nsss(0) <='0';
          end if;
        if(cVar1S15S76P014P024P044P027(0)='1' AND  B(20)='0' AND A(10)='0' AND A(20)='1' )then
          cVar2S15S76N036P019P018nsss(0) <='1';
          else
          cVar2S15S76N036P019P018nsss(0) <='0';
          end if;
        if(cVar1S16S76P014P024P044P062(0)='1' AND  A(11)='0' AND A(10)='1' )then
          cVar2S16S76P017P019nsss(0) <='1';
          else
          cVar2S16S76P017P019nsss(0) <='0';
          end if;
        if(cVar1S18S76P014P024P031N045(0)='1' AND  A(23)='0' AND A(18)='0' AND E(21)='1' )then
          cVar2S18S76P012P003P049nsss(0) <='1';
          else
          cVar2S18S76P012P003P049nsss(0) <='0';
          end if;
        if(cVar1S19S76P014P024P031N045(0)='1' AND  A(23)='1' AND A(29)='1' )then
          cVar2S19S76P012P000nsss(0) <='1';
          else
          cVar2S19S76P012P000nsss(0) <='0';
          end if;
        if(cVar1S0S77P010P024P028P003(0)='1' AND  E(19)='1' )then
          cVar2S0S77P057nsss(0) <='1';
          else
          cVar2S0S77P057nsss(0) <='0';
          end if;
        if(cVar1S1S77P010P024P028P003(0)='1' AND  E(19)='0' AND E(20)='1' )then
          cVar2S1S77N057P053nsss(0) <='1';
          else
          cVar2S1S77N057P053nsss(0) <='0';
          end if;
        if(cVar1S2S77P010P024P028P003(0)='1' AND  E(19)='0' AND E(20)='0' AND A(13)='0' )then
          cVar2S2S77N057N053P013nsss(0) <='1';
          else
          cVar2S2S77N057N053P013nsss(0) <='0';
          end if;
        if(cVar1S3S77P010P024N028P045(0)='1' AND  B(13)='1' )then
          cVar2S3S77P031nsss(0) <='1';
          else
          cVar2S3S77P031nsss(0) <='0';
          end if;
        if(cVar1S4S77P010P024N028P045(0)='1' AND  B(13)='0' AND B(16)='0' )then
          cVar2S4S77N031P025nsss(0) <='1';
          else
          cVar2S4S77N031P025nsss(0) <='0';
          end if;
        if(cVar1S5S77P010P024N028P045(0)='1' AND  A(20)='1' )then
          cVar2S5S77P018nsss(0) <='1';
          else
          cVar2S5S77P018nsss(0) <='0';
          end if;
        if(cVar1S6S77P010P024P064P019(0)='1' AND  B(20)='0' AND B(21)='1' )then
          cVar2S6S77P036P034nsss(0) <='1';
          else
          cVar2S6S77P036P034nsss(0) <='0';
          end if;
        if(cVar1S7S77P010P024P064P019(0)='1' AND  B(20)='0' AND B(21)='0' AND A(11)='0' )then
          cVar2S7S77P036N034P017nsss(0) <='1';
          else
          cVar2S7S77P036N034P017nsss(0) <='0';
          end if;
        if(cVar1S10S77N010P025N046N007(0)='1' AND  B(26)='1' )then
          cVar2S10S77P024nsss(0) <='1';
          else
          cVar2S10S77P024nsss(0) <='0';
          end if;
        if(cVar1S11S77N010P025N046N007(0)='1' AND  B(26)='0' AND A(11)='0' AND A(22)='1' )then
          cVar2S11S77N024P017P014nsss(0) <='1';
          else
          cVar2S11S77N024P017P014nsss(0) <='0';
          end if;
        if(cVar1S12S77N010N025P046P002(0)='1' AND  E(15)='1' )then
          cVar2S12S77P040nsss(0) <='1';
          else
          cVar2S12S77P040nsss(0) <='0';
          end if;
        if(cVar1S13S77N010N025P046P002(0)='1' AND  E(15)='0' AND A(14)='0' )then
          cVar2S13S77N040P011nsss(0) <='1';
          else
          cVar2S13S77N040P011nsss(0) <='0';
          end if;
        if(cVar1S14S77N010N025P046P002(0)='1' AND  E(15)='0' AND A(14)='1' AND A(26)='1' )then
          cVar2S14S77N040P011P006nsss(0) <='1';
          else
          cVar2S14S77N040P011P006nsss(0) <='0';
          end if;
        if(cVar1S15S77N010N025P046N002(0)='1' AND  B(28)='1' AND D(23)='1' )then
          cVar2S15S77P020P039nsss(0) <='1';
          else
          cVar2S15S77P020P039nsss(0) <='0';
          end if;
        if(cVar1S17S77N010N025P046N047(0)='1' AND  D(16)='1' AND A(20)='1' )then
          cVar2S17S77P067P018nsss(0) <='1';
          else
          cVar2S17S77P067P018nsss(0) <='0';
          end if;
        if(cVar1S18S77N010N025P046N047(0)='1' AND  D(16)='0' AND A(15)='1' )then
          cVar2S18S77N067P009nsss(0) <='1';
          else
          cVar2S18S77N067P009nsss(0) <='0';
          end if;
        if(cVar1S19S77N010N025P046N047(0)='1' AND  D(16)='0' AND A(15)='0' AND A(25)='1' )then
          cVar2S19S77N067N009P008nsss(0) <='1';
          else
          cVar2S19S77N067N009P008nsss(0) <='0';
          end if;
        if(cVar1S0S78P039P041P020P050(0)='1' AND  D(22)='0' AND B(18)='0' )then
          cVar2S0S78P043P021nsss(0) <='1';
          else
          cVar2S0S78P043P021nsss(0) <='0';
          end if;
        if(cVar1S1S78P039P041P020N050(0)='1' AND  B(18)='1' AND E(15)='1' )then
          cVar2S1S78P021P040nsss(0) <='1';
          else
          cVar2S1S78P021P040nsss(0) <='0';
          end if;
        if(cVar1S2S78P039P041P020N050(0)='1' AND  B(18)='1' AND E(15)='0' AND A(26)='1' )then
          cVar2S2S78P021N040P006nsss(0) <='1';
          else
          cVar2S2S78P021N040P006nsss(0) <='0';
          end if;
        if(cVar1S3S78P039P041P020N050(0)='1' AND  B(18)='0' AND D(15)='0' AND E(15)='0' )then
          cVar2S3S78N021P038P040nsss(0) <='1';
          else
          cVar2S3S78N021P038P040nsss(0) <='0';
          end if;
        if(cVar1S5S78P039P041P020N040(0)='1' AND  B(27)='0' AND E( 9)='0' AND A(16)='1' )then
          cVar2S5S78P022P064P007nsss(0) <='1';
          else
          cVar2S5S78P022P064P007nsss(0) <='0';
          end if;
        if(cVar1S6S78P039P041P020N040(0)='1' AND  B(27)='0' AND E( 9)='1' AND A(22)='1' )then
          cVar2S6S78P022P064P014nsss(0) <='1';
          else
          cVar2S6S78P022P064P014nsss(0) <='0';
          end if;
        if(cVar1S9S78P039N020P012P060(0)='1' AND  B(18)='1' )then
          cVar2S9S78P021nsss(0) <='1';
          else
          cVar2S9S78P021nsss(0) <='0';
          end if;
        if(cVar1S10S78P039N020P012P060(0)='1' AND  B(18)='0' AND A(25)='0' AND A(15)='1' )then
          cVar2S10S78N021P008P009nsss(0) <='1';
          else
          cVar2S10S78N021P008P009nsss(0) <='0';
          end if;
        if(cVar1S1S79P021N040P048P060(0)='1' AND  E(19)='0' AND B(28)='0' )then
          cVar2S1S79P057P020nsss(0) <='1';
          else
          cVar2S1S79P057P020nsss(0) <='0';
          end if;
        if(cVar1S2S79N021P038P040P050(0)='1' AND  D(22)='0' AND E(13)='1' )then
          cVar2S2S79P043P048nsss(0) <='1';
          else
          cVar2S2S79P043P048nsss(0) <='0';
          end if;
        if(cVar1S3S79N021P038P040P050(0)='1' AND  D(22)='0' AND E(13)='0' AND E(12)='1' )then
          cVar2S3S79P043N048P052nsss(0) <='1';
          else
          cVar2S3S79P043N048P052nsss(0) <='0';
          end if;
        if(cVar1S4S79N021P038P040N050(0)='1' AND  D(21)='1' AND B(26)='1' AND A(21)='0' )then
          cVar2S4S79P047P024P016nsss(0) <='1';
          else
          cVar2S4S79P047P024P016nsss(0) <='0';
          end if;
        if(cVar1S5S79N021P038P040N050(0)='1' AND  D(21)='1' AND B(26)='0' AND E(11)='0' )then
          cVar2S5S79P047N024P056nsss(0) <='1';
          else
          cVar2S5S79P047N024P056nsss(0) <='0';
          end if;
        if(cVar1S6S79N021P038P040N050(0)='1' AND  D(21)='0' AND E(21)='0' AND D(10)='1' )then
          cVar2S6S79N047P049P058nsss(0) <='1';
          else
          cVar2S6S79N047P049P058nsss(0) <='0';
          end if;
        if(cVar1S7S79N021P038P040N050(0)='1' AND  D(21)='0' AND E(21)='1' AND A(20)='1' )then
          cVar2S7S79N047P049P018nsss(0) <='1';
          else
          cVar2S7S79N047P049P018nsss(0) <='0';
          end if;
        if(cVar1S8S79N021P038P040P059(0)='1' AND  A(20)='1' AND D(14)='1' )then
          cVar2S8S79P018P042nsss(0) <='1';
          else
          cVar2S8S79P018P042nsss(0) <='0';
          end if;
        if(cVar1S9S79N021P038P040P059(0)='1' AND  A(20)='1' AND D(14)='0' AND A(12)='0' )then
          cVar2S9S79P018N042P015nsss(0) <='1';
          else
          cVar2S9S79P018N042P015nsss(0) <='0';
          end if;
        if(cVar1S10S79N021P038P040P059(0)='1' AND  A(20)='0' AND B(10)='1' )then
          cVar2S10S79N018P037nsss(0) <='1';
          else
          cVar2S10S79N018P037nsss(0) <='0';
          end if;
        if(cVar1S12S79N021P038P065N020(0)='1' AND  B(20)='0' AND A(20)='1' AND A(12)='1' )then
          cVar2S12S79P036P018P015nsss(0) <='1';
          else
          cVar2S12S79P036P018P015nsss(0) <='0';
          end if;
        if(cVar1S13S79N021P038P065N020(0)='1' AND  B(20)='0' AND A(20)='0' AND A(23)='1' )then
          cVar2S13S79P036N018P012nsss(0) <='1';
          else
          cVar2S13S79P036N018P012nsss(0) <='0';
          end if;
        if(cVar1S2S80P037P048N025N027(0)='1' AND  D( 9)='1' AND A(10)='0' )then
          cVar2S2S80P062P019nsss(0) <='1';
          else
          cVar2S2S80P062P019nsss(0) <='0';
          end if;
        if(cVar1S3S80P037P048N025N027(0)='1' AND  D( 9)='0' AND D(21)='1' )then
          cVar2S3S80N062P047nsss(0) <='1';
          else
          cVar2S3S80N062P047nsss(0) <='0';
          end if;
        if(cVar1S4S80P037P048N025N027(0)='1' AND  D( 9)='0' AND D(21)='0' AND A(20)='1' )then
          cVar2S4S80N062N047P018nsss(0) <='1';
          else
          cVar2S4S80N062N047P018nsss(0) <='0';
          end if;
        if(cVar1S5S80P037N048P046P064(0)='1' AND  A(10)='1' AND D(16)='0' AND E(17)='0' )then
          cVar2S5S80P019P067P065nsss(0) <='1';
          else
          cVar2S5S80P019P067P065nsss(0) <='0';
          end if;
        if(cVar1S6S80P037N048P046P064(0)='1' AND  A(10)='0' AND E(19)='1' AND E(20)='0' )then
          cVar2S6S80N019P057P053nsss(0) <='1';
          else
          cVar2S6S80N019P057P053nsss(0) <='0';
          end if;
        if(cVar1S7S80P037N048P046P064(0)='1' AND  A(10)='0' AND E(19)='0' AND B(13)='0' )then
          cVar2S7S80N019N057P031nsss(0) <='1';
          else
          cVar2S7S80N019N057P031nsss(0) <='0';
          end if;
        if(cVar1S8S80P037N048P046P064(0)='1' AND  A(11)='0' AND D(16)='1' AND E(17)='0' )then
          cVar2S8S80P017P067P065nsss(0) <='1';
          else
          cVar2S8S80P017P067P065nsss(0) <='0';
          end if;
        if(cVar1S9S80P037N048P046P064(0)='1' AND  A(11)='0' AND D(16)='0' AND D( 8)='1' )then
          cVar2S9S80P017N067P066nsss(0) <='1';
          else
          cVar2S9S80P017N067P066nsss(0) <='0';
          end if;
        if(cVar1S10S80P037N048P046P064(0)='1' AND  A(11)='1' AND B(11)='1' AND D(17)='1' )then
          cVar2S10S80P017P035P063nsss(0) <='1';
          else
          cVar2S10S80P017P035P063nsss(0) <='0';
          end if;
        if(cVar1S11S80P037N048P046P003(0)='1' AND  E(14)='1' AND A(11)='0' )then
          cVar2S11S80P044P017nsss(0) <='1';
          else
          cVar2S11S80P044P017nsss(0) <='0';
          end if;
        if(cVar1S12S80P037N048P046P003(0)='1' AND  E(14)='0' AND A(11)='1' )then
          cVar2S12S80N044P017nsss(0) <='1';
          else
          cVar2S12S80N044P017nsss(0) <='0';
          end if;
        if(cVar1S13S80P037P013P048P064(0)='1' AND  A(18)='0' AND D(10)='0' )then
          cVar2S13S80P003P058nsss(0) <='1';
          else
          cVar2S13S80P003P058nsss(0) <='0';
          end if;
        if(cVar1S14S80P037P013P048P064(0)='1' AND  A(18)='0' AND D(10)='1' AND E(10)='1' )then
          cVar2S14S80P003P058P060nsss(0) <='1';
          else
          cVar2S14S80P003P058P060nsss(0) <='0';
          end if;
        if(cVar1S15S80P037P013P048N064(0)='1' AND  E(23)='1' )then
          cVar2S15S80P041nsss(0) <='1';
          else
          cVar2S15S80P041nsss(0) <='0';
          end if;
        if(cVar1S16S80P037P013P048N064(0)='1' AND  E(23)='0' AND D(23)='0' AND A(25)='1' )then
          cVar2S16S80N041P039P008nsss(0) <='1';
          else
          cVar2S16S80N041P039P008nsss(0) <='0';
          end if;
        if(cVar1S17S80P037P013P048P035(0)='1' AND  D(13)='1' )then
          cVar2S17S80P046nsss(0) <='1';
          else
          cVar2S17S80P046nsss(0) <='0';
          end if;
        if(cVar1S18S80P037P013P018P015(0)='1' AND  A(22)='1' )then
          cVar2S18S80P014nsss(0) <='1';
          else
          cVar2S18S80P014nsss(0) <='0';
          end if;
        if(cVar1S19S80P037P013P018P015(0)='1' AND  A(22)='0' AND A(10)='0' )then
          cVar2S19S80N014P019nsss(0) <='1';
          else
          cVar2S19S80N014P019nsss(0) <='0';
          end if;
        if(cVar1S20S80P037P013P018P015(0)='1' AND  A(22)='0' AND A(25)='0' AND A(11)='0' )then
          cVar2S20S80P014P008P017nsss(0) <='1';
          else
          cVar2S20S80P014P008P017nsss(0) <='0';
          end if;
        if(cVar1S21S80P037P013P018P015(0)='1' AND  A(22)='1' AND A(10)='1' AND E(16)='1' )then
          cVar2S21S80P014P019P069nsss(0) <='1';
          else
          cVar2S21S80P014P019P069nsss(0) <='0';
          end if;
        if(cVar1S23S80P037P013N018N031(0)='1' AND  A(23)='1' AND D(20)='0' AND A(24)='0' )then
          cVar2S23S80P012P051P010nsss(0) <='1';
          else
          cVar2S23S80P012P051P010nsss(0) <='0';
          end if;
        if(cVar1S24S80P037P013N018N031(0)='1' AND  A(23)='0' AND E(16)='1' AND A(25)='0' )then
          cVar2S24S80N012P069P008nsss(0) <='1';
          else
          cVar2S24S80N012P069P008nsss(0) <='0';
          end if;
        if(cVar1S0S81P019P017P055P053(0)='1' AND  E(18)='0' )then
          cVar2S0S81P061nsss(0) <='1';
          else
          cVar2S0S81P061nsss(0) <='0';
          end if;
        if(cVar1S1S81P019P017N055P057(0)='1' AND  E(20)='1' AND A(22)='1' )then
          cVar2S1S81P053P014nsss(0) <='1';
          else
          cVar2S1S81P053P014nsss(0) <='0';
          end if;
        if(cVar1S2S81P019P017N055P057(0)='1' AND  E(20)='1' AND A(22)='0' AND A(23)='0' )then
          cVar2S2S81P053N014P012nsss(0) <='1';
          else
          cVar2S2S81P053N014P012nsss(0) <='0';
          end if;
        if(cVar1S3S81P019P017N055P057(0)='1' AND  E(20)='0' AND B(11)='1' )then
          cVar2S3S81N053P035nsss(0) <='1';
          else
          cVar2S3S81N053P035nsss(0) <='0';
          end if;
        if(cVar1S4S81P019P017N055P057(0)='1' AND  E(20)='0' AND B(11)='0' AND A(12)='0' )then
          cVar2S4S81N053N035P015nsss(0) <='1';
          else
          cVar2S4S81N053N035P015nsss(0) <='0';
          end if;
        if(cVar1S5S81P019P017N055P057(0)='1' AND  A(21)='0' AND D(18)='1' )then
          cVar2S5S81P016P059nsss(0) <='1';
          else
          cVar2S5S81P016P059nsss(0) <='0';
          end if;
        if(cVar1S6S81P019P017P064P029(0)='1' AND  D(17)='0' AND E(11)='0' AND E(17)='0' )then
          cVar2S6S81P063P056P065nsss(0) <='1';
          else
          cVar2S6S81P063P056P065nsss(0) <='0';
          end if;
        if(cVar1S7S81P019P017P064P029(0)='1' AND  D(17)='0' AND E(11)='1' AND D( 8)='1' )then
          cVar2S7S81P063P056P066nsss(0) <='1';
          else
          cVar2S7S81P063P056P066nsss(0) <='0';
          end if;
        if(cVar1S8S81P019P017P064P029(0)='1' AND  D(17)='1' AND B(26)='0' AND A(18)='1' )then
          cVar2S8S81P063P024P003nsss(0) <='1';
          else
          cVar2S8S81P063P024P003nsss(0) <='0';
          end if;
        if(cVar1S9S81P019P017P064P029(0)='1' AND  A(23)='0' AND A(20)='1' )then
          cVar2S9S81P012P018nsss(0) <='1';
          else
          cVar2S9S81P012P018nsss(0) <='0';
          end if;
        if(cVar1S10S81P019P017P064P011(0)='1' AND  B(20)='1' )then
          cVar2S10S81P036nsss(0) <='1';
          else
          cVar2S10S81P036nsss(0) <='0';
          end if;
        if(cVar1S11S81P019P017P064P011(0)='1' AND  B(20)='0' AND A(20)='1' )then
          cVar2S11S81N036P018nsss(0) <='1';
          else
          cVar2S11S81N036P018nsss(0) <='0';
          end if;
        if(cVar1S12S81P019P017P064N011(0)='1' AND  D( 9)='1' AND D(17)='1' AND A(20)='1' )then
          cVar2S12S81P062P063P018nsss(0) <='1';
          else
          cVar2S12S81P062P063P018nsss(0) <='0';
          end if;
        if(cVar1S13S81N019P037P003P035(0)='1' AND  B(13)='1' )then
          cVar2S13S81P031nsss(0) <='1';
          else
          cVar2S13S81P031nsss(0) <='0';
          end if;
        if(cVar1S14S81N019P037P003P035(0)='1' AND  B(13)='0' AND A(13)='0' AND E(10)='0' )then
          cVar2S14S81N031P013P060nsss(0) <='1';
          else
          cVar2S14S81N031P013P060nsss(0) <='0';
          end if;
        if(cVar1S15S81N019P037P003P035(0)='1' AND  B(13)='0' AND A(13)='1' AND D(16)='1' )then
          cVar2S15S81N031P013P067nsss(0) <='1';
          else
          cVar2S15S81N031P013P067nsss(0) <='0';
          end if;
        if(cVar1S16S81N019P037P003P035(0)='1' AND  A(17)='0' AND D(16)='0' AND D( 8)='1' )then
          cVar2S16S81P005P067P066nsss(0) <='1';
          else
          cVar2S16S81P005P067P066nsss(0) <='0';
          end if;
        if(cVar1S17S81N019P037P003P035(0)='1' AND  A(17)='0' AND D(16)='1' AND D( 9)='1' )then
          cVar2S17S81P005P067P062nsss(0) <='1';
          else
          cVar2S17S81P005P067P062nsss(0) <='0';
          end if;
        if(cVar1S19S81N019P037P003N034(0)='1' AND  B(20)='0' AND A(21)='0' AND A(13)='1' )then
          cVar2S19S81P036N016P013nsss(0) <='1';
          else
          cVar2S19S81P036N016P013nsss(0) <='0';
          end if;
        if(cVar1S21S81N019N037P048N062(0)='1' AND  B(15)='1' )then
          cVar2S21S81P027nsss(0) <='1';
          else
          cVar2S21S81P027nsss(0) <='0';
          end if;
        if(cVar1S22S81N019N037P048N062(0)='1' AND  B(15)='0' AND B(16)='1' )then
          cVar2S22S81N027P025nsss(0) <='1';
          else
          cVar2S22S81N027P025nsss(0) <='0';
          end if;
        if(cVar1S23S81N019N037P048N062(0)='1' AND  B(15)='0' AND B(16)='0' AND D(11)='1' )then
          cVar2S23S81N027N025P054nsss(0) <='1';
          else
          cVar2S23S81N027N025P054nsss(0) <='0';
          end if;
        if(cVar1S24S81N019N037N048P057(0)='1' AND  A(13)='1' AND A(23)='0' )then
          cVar2S24S81P013P012nsss(0) <='1';
          else
          cVar2S24S81P013P012nsss(0) <='0';
          end if;
        if(cVar1S25S81N019N037N048P057(0)='1' AND  A(13)='0' AND A(14)='1' )then
          cVar2S25S81N013P011nsss(0) <='1';
          else
          cVar2S25S81N013P011nsss(0) <='0';
          end if;
        if(cVar1S26S81N019N037N048P057(0)='1' AND  A(13)='0' AND A(14)='0' AND A(12)='0' )then
          cVar2S26S81N013N011P015nsss(0) <='1';
          else
          cVar2S26S81N013N011P015nsss(0) <='0';
          end if;
        if(cVar1S27S81N019N037N048N057(0)='1' AND  A(12)='1' AND A(27)='0' AND B(11)='1' )then
          cVar2S27S81P015P004P035nsss(0) <='1';
          else
          cVar2S27S81P015P004P035nsss(0) <='0';
          end if;
        if(cVar1S28S81N019N037N048N057(0)='1' AND  A(12)='1' AND A(27)='1' AND A(13)='1' )then
          cVar2S28S81P015P004P013nsss(0) <='1';
          else
          cVar2S28S81P015P004P013nsss(0) <='0';
          end if;
        if(cVar1S29S81N019N037N048N057(0)='1' AND  A(12)='0' AND D(20)='1' AND A(14)='1' )then
          cVar2S29S81N015P051P011nsss(0) <='1';
          else
          cVar2S29S81N015P051P011nsss(0) <='0';
          end if;
        if(cVar1S1S82P019P030P040N021(0)='1' AND  A(28)='1' )then
          cVar2S1S82P002nsss(0) <='1';
          else
          cVar2S1S82P002nsss(0) <='0';
          end if;
        if(cVar1S2S82P019P030P040N021(0)='1' AND  A(28)='0' AND D( 8)='0' AND A(20)='1' )then
          cVar2S2S82N002P066P018nsss(0) <='1';
          else
          cVar2S2S82N002P066P018nsss(0) <='0';
          end if;
        if(cVar1S3S82P019P030N040P038(0)='1' AND  B(18)='0' AND D(12)='1' )then
          cVar2S3S82P021P050nsss(0) <='1';
          else
          cVar2S3S82P021P050nsss(0) <='0';
          end if;
        if(cVar1S4S82P019P030N040P038(0)='1' AND  B(18)='0' AND D(12)='0' AND D(19)='0' )then
          cVar2S4S82P021N050P055nsss(0) <='1';
          else
          cVar2S4S82P021N050P055nsss(0) <='0';
          end if;
        if(cVar1S5S82P019P030N040P038(0)='1' AND  B(18)='1' AND A(26)='1' )then
          cVar2S5S82P021P006nsss(0) <='1';
          else
          cVar2S5S82P021P006nsss(0) <='0';
          end if;
        if(cVar1S7S82P019P030P045N056(0)='1' AND  A(28)='1' )then
          cVar2S7S82P002nsss(0) <='1';
          else
          cVar2S7S82P002nsss(0) <='0';
          end if;
        if(cVar1S8S82P019P030P045N056(0)='1' AND  A(28)='0' AND E(19)='1' AND A(22)='0' )then
          cVar2S8S82N002P057P014nsss(0) <='1';
          else
          cVar2S8S82N002P057P014nsss(0) <='0';
          end if;
        if(cVar1S9S82P019P030P045N056(0)='1' AND  A(28)='0' AND E(19)='0' AND A(16)='1' )then
          cVar2S9S82N002N057P007nsss(0) <='1';
          else
          cVar2S9S82N002N057P007nsss(0) <='0';
          end if;
        if(cVar1S11S82P019P017P055N065(0)='1' AND  D(18)='0' AND E(20)='0' )then
          cVar2S11S82P059P053nsss(0) <='1';
          else
          cVar2S11S82P059P053nsss(0) <='0';
          end if;
        if(cVar1S12S82P019P017N055P057(0)='1' AND  E(20)='1' AND A(22)='1' )then
          cVar2S12S82P053P014nsss(0) <='1';
          else
          cVar2S12S82P053P014nsss(0) <='0';
          end if;
        if(cVar1S13S82P019P017N055P057(0)='1' AND  E(20)='1' AND A(22)='0' AND A(21)='0' )then
          cVar2S13S82P053N014P016nsss(0) <='1';
          else
          cVar2S13S82P053N014P016nsss(0) <='0';
          end if;
        if(cVar1S14S82P019P017N055P057(0)='1' AND  E(20)='0' AND E(18)='1' )then
          cVar2S14S82N053P061nsss(0) <='1';
          else
          cVar2S14S82N053P061nsss(0) <='0';
          end if;
        if(cVar1S15S82P019P017N055P057(0)='1' AND  A(21)='0' AND D(18)='1' )then
          cVar2S15S82P016P059nsss(0) <='1';
          else
          cVar2S15S82P016P059nsss(0) <='0';
          end if;
        if(cVar1S16S82P019P017P053P029(0)='1' AND  B(13)='1' AND A(25)='0' )then
          cVar2S16S82P031P008nsss(0) <='1';
          else
          cVar2S16S82P031P008nsss(0) <='0';
          end if;
        if(cVar1S17S82P019P017P053P029(0)='1' AND  B(13)='0' AND B(26)='1' AND A(21)='0' )then
          cVar2S17S82N031P024P016nsss(0) <='1';
          else
          cVar2S17S82N031P024P016nsss(0) <='0';
          end if;
        if(cVar1S18S82P019P017P053P037(0)='1' AND  A(22)='0' )then
          cVar2S18S82P014nsss(0) <='1';
          else
          cVar2S18S82P014nsss(0) <='0';
          end if;
        if(cVar1S19S82P019P017P053N037(0)='1' AND  A(25)='1' )then
          cVar2S19S82P008nsss(0) <='1';
          else
          cVar2S19S82P008nsss(0) <='0';
          end if;
        if(cVar1S0S83P015P051P017P012(0)='1' AND  A(18)='0' AND B(21)='0' AND B(26)='0' )then
          cVar2S0S83P003P034P024nsss(0) <='1';
          else
          cVar2S0S83P003P034P024nsss(0) <='0';
          end if;
        if(cVar1S1S83P015P051P017P012(0)='1' AND  A(18)='1' AND A(20)='0' AND A(21)='1' )then
          cVar2S1S83P003P018P016nsss(0) <='1';
          else
          cVar2S1S83P003P018P016nsss(0) <='0';
          end if;
        if(cVar1S2S83P015P051P017N012(0)='1' AND  E(18)='1' AND B(12)='1' )then
          cVar2S2S83P061P033nsss(0) <='1';
          else
          cVar2S2S83P061P033nsss(0) <='0';
          end if;
        if(cVar1S3S83P015P051P017N012(0)='1' AND  E(18)='1' AND B(12)='0' AND A(20)='1' )then
          cVar2S3S83P061N033P018nsss(0) <='1';
          else
          cVar2S3S83P061N033P018nsss(0) <='0';
          end if;
        if(cVar1S4S83P015P051P017N012(0)='1' AND  E(18)='0' AND B(22)='1' AND A(14)='0' )then
          cVar2S4S83N061P032P011nsss(0) <='1';
          else
          cVar2S4S83N061P032P011nsss(0) <='0';
          end if;
        if(cVar1S5S83P015P051P017N012(0)='1' AND  E(18)='0' AND B(22)='0' AND B(21)='1' )then
          cVar2S5S83N061N032P034nsss(0) <='1';
          else
          cVar2S5S83N061N032P034nsss(0) <='0';
          end if;
        if(cVar1S6S83P015P051P017P061(0)='1' AND  B(12)='0' AND A(15)='0' AND E(17)='0' )then
          cVar2S6S83P033P009P065nsss(0) <='1';
          else
          cVar2S6S83P033P009P065nsss(0) <='0';
          end if;
        if(cVar1S7S83P015P051P017P061(0)='1' AND  B(12)='1' AND B(10)='0' AND E( 8)='1' )then
          cVar2S7S83P033P037P068nsss(0) <='1';
          else
          cVar2S7S83P033P037P068nsss(0) <='0';
          end if;
        if(cVar1S8S83P015P051P017P061(0)='1' AND  E(10)='1' )then
          cVar2S8S83P060nsss(0) <='1';
          else
          cVar2S8S83P060nsss(0) <='0';
          end if;
        if(cVar1S9S83P015P051P053P000(0)='1' AND  B(20)='1' )then
          cVar2S9S83P036nsss(0) <='1';
          else
          cVar2S9S83P036nsss(0) <='0';
          end if;
        if(cVar1S10S83P015P051P053P000(0)='1' AND  B(20)='0' AND E(16)='0' AND A(14)='1' )then
          cVar2S10S83N036P069P011nsss(0) <='1';
          else
          cVar2S10S83N036P069P011nsss(0) <='0';
          end if;
        if(cVar1S11S83P015P051N053P014(0)='1' AND  B(11)='1' )then
          cVar2S11S83P035nsss(0) <='1';
          else
          cVar2S11S83P035nsss(0) <='0';
          end if;
        if(cVar1S13S83N015P021N038P069(0)='1' AND  A(13)='0' AND A(23)='1' )then
          cVar2S13S83P013P012nsss(0) <='1';
          else
          cVar2S13S83P013P012nsss(0) <='0';
          end if;
        if(cVar1S14S83N015P021N038P069(0)='1' AND  A(13)='0' AND A(23)='0' AND A(10)='1' )then
          cVar2S14S83P013N012P019nsss(0) <='1';
          else
          cVar2S14S83P013N012P019nsss(0) <='0';
          end if;
        if(cVar1S15S83N015N021P038P067(0)='1' AND  B(25)='0' AND B(11)='0' )then
          cVar2S15S83P026P035nsss(0) <='1';
          else
          cVar2S15S83P026P035nsss(0) <='0';
          end if;
        if(cVar1S16S83N015N021P038P067(0)='1' AND  B(25)='0' AND B(11)='1' AND A(22)='1' )then
          cVar2S16S83P026P035P014nsss(0) <='1';
          else
          cVar2S16S83P026P035P014nsss(0) <='0';
          end if;
        if(cVar1S17S83N015N021P038P067(0)='1' AND  B(25)='1' AND E( 8)='0' AND A(20)='1' )then
          cVar2S17S83P026P068P018nsss(0) <='1';
          else
          cVar2S17S83P026P068P018nsss(0) <='0';
          end if;
        if(cVar1S18S83N015N021P038N067(0)='1' AND  D(20)='1' AND A(14)='1' AND D( 8)='0' )then
          cVar2S18S83P051P011P066nsss(0) <='1';
          else
          cVar2S18S83P051P011P066nsss(0) <='0';
          end if;
        if(cVar1S19S83N015N021P038N067(0)='1' AND  D(20)='1' AND A(14)='0' AND A(25)='1' )then
          cVar2S19S83P051N011P008nsss(0) <='1';
          else
          cVar2S19S83P051N011P008nsss(0) <='0';
          end if;
        if(cVar1S20S83N015N021P038N067(0)='1' AND  D(20)='0' AND E(20)='0' AND D(21)='1' )then
          cVar2S20S83N051P053P047nsss(0) <='1';
          else
          cVar2S20S83N051P053P047nsss(0) <='0';
          end if;
        if(cVar1S21S83N015N021P038P069(0)='1' AND  A(22)='0' AND A(23)='1' )then
          cVar2S21S83P014P012nsss(0) <='1';
          else
          cVar2S21S83P014P012nsss(0) <='0';
          end if;
        if(cVar1S22S83N015N021P038P069(0)='1' AND  A(22)='0' AND A(23)='0' AND E(15)='1' )then
          cVar2S22S83P014N012P040nsss(0) <='1';
          else
          cVar2S22S83P014N012P040nsss(0) <='0';
          end if;
        if(cVar1S1S84P067P037P021N040(0)='1' AND  E( 9)='1' )then
          cVar2S1S84P064nsss(0) <='1';
          else
          cVar2S1S84P064nsss(0) <='0';
          end if;
        if(cVar1S2S84P067P037P021N040(0)='1' AND  E( 9)='0' AND A(14)='0' AND D( 8)='0' )then
          cVar2S2S84N064P011P066nsss(0) <='1';
          else
          cVar2S2S84N064P011P066nsss(0) <='0';
          end if;
        if(cVar1S3S84P067P037N021P013(0)='1' AND  B(13)='1' AND A(14)='0' )then
          cVar2S3S84P031P011nsss(0) <='1';
          else
          cVar2S3S84P031P011nsss(0) <='0';
          end if;
        if(cVar1S4S84P067P037N021P013(0)='1' AND  B(13)='0' AND B(14)='1' AND A(12)='0' )then
          cVar2S4S84N031P029P015nsss(0) <='1';
          else
          cVar2S4S84N031P029P015nsss(0) <='0';
          end if;
        if(cVar1S5S84P067P037N021P013(0)='1' AND  B(13)='0' AND B(14)='0' AND E(11)='0' )then
          cVar2S5S84N031N029P056nsss(0) <='1';
          else
          cVar2S5S84N031N029P056nsss(0) <='0';
          end if;
        if(cVar1S6S84P067P037N021N013(0)='1' AND  B(13)='0' AND B(22)='0' AND D(10)='0' )then
          cVar2S6S84P031P032P058nsss(0) <='1';
          else
          cVar2S6S84P031P032P058nsss(0) <='0';
          end if;
        if(cVar1S7S84P067P037N021N013(0)='1' AND  B(13)='0' AND B(22)='1' AND D(18)='0' )then
          cVar2S7S84P031P032P059nsss(0) <='1';
          else
          cVar2S7S84P031P032P059nsss(0) <='0';
          end if;
        if(cVar1S8S84P067P037N021N013(0)='1' AND  B(13)='1' AND A(23)='1' AND A(22)='0' )then
          cVar2S8S84P031P012P014nsss(0) <='1';
          else
          cVar2S8S84P031P012P014nsss(0) <='0';
          end if;
        if(cVar1S10S84P067P037N028P013(0)='1' AND  E(13)='0' AND A(29)='1' AND A(11)='0' )then
          cVar2S10S84P048P000P017nsss(0) <='1';
          else
          cVar2S10S84P048P000P017nsss(0) <='0';
          end if;
        if(cVar1S11S84P067P037N028P013(0)='1' AND  E(13)='0' AND A(29)='0' AND D(20)='1' )then
          cVar2S11S84P048N000P051nsss(0) <='1';
          else
          cVar2S11S84P048N000P051nsss(0) <='0';
          end if;
        if(cVar1S12S84P067P037N028P013(0)='1' AND  E(13)='1' AND D(13)='1' )then
          cVar2S12S84P048P046nsss(0) <='1';
          else
          cVar2S12S84P048P046nsss(0) <='0';
          end if;
        if(cVar1S13S84P067P037N028P013(0)='1' AND  A(20)='1' AND A(27)='0' AND A(15)='1' )then
          cVar2S13S84P018P004P009nsss(0) <='1';
          else
          cVar2S13S84P018P004P009nsss(0) <='0';
          end if;
        if(cVar1S14S84P067P037N028P013(0)='1' AND  A(20)='0' AND B(13)='1' )then
          cVar2S14S84N018P031nsss(0) <='1';
          else
          cVar2S14S84N018P031nsss(0) <='0';
          end if;
        if(cVar1S15S84P067P051P065P010(0)='1' AND  E( 8)='0' AND B(22)='0' )then
          cVar2S15S84P068P032nsss(0) <='1';
          else
          cVar2S15S84P068P032nsss(0) <='0';
          end if;
        if(cVar1S16S84P067P051P065P010(0)='1' AND  E( 8)='1' AND A(23)='1' )then
          cVar2S16S84P068P012nsss(0) <='1';
          else
          cVar2S16S84P068P012nsss(0) <='0';
          end if;
        if(cVar1S17S84P067P051P065P010(0)='1' AND  A(12)='1' AND A(20)='1' )then
          cVar2S17S84P015P018nsss(0) <='1';
          else
          cVar2S17S84P015P018nsss(0) <='0';
          end if;
        if(cVar1S18S84P067P051N065P064(0)='1' AND  D(10)='0' AND A(15)='0' AND A(23)='0' )then
          cVar2S18S84P058P009P012nsss(0) <='1';
          else
          cVar2S18S84P058P009P012nsss(0) <='0';
          end if;
        if(cVar1S19S84P067P051N065N064(0)='1' AND  E(12)='1' AND A(14)='0' )then
          cVar2S19S84P052P011nsss(0) <='1';
          else
          cVar2S19S84P052P011nsss(0) <='0';
          end if;
        if(cVar1S20S84P067P051N065N064(0)='1' AND  E(12)='0' AND D(17)='0' AND D(18)='1' )then
          cVar2S20S84N052P063P059nsss(0) <='1';
          else
          cVar2S20S84N052P063P059nsss(0) <='0';
          end if;
        if(cVar1S21S84P067P051N065N064(0)='1' AND  E(12)='0' AND D(17)='1' AND B(26)='1' )then
          cVar2S21S84N052P063P024nsss(0) <='1';
          else
          cVar2S21S84N052P063P024nsss(0) <='0';
          end if;
        if(cVar1S22S84P067P051P006P034(0)='1' AND  A(29)='0' AND B(24)='1' )then
          cVar2S22S84P000P028nsss(0) <='1';
          else
          cVar2S22S84P000P028nsss(0) <='0';
          end if;
        if(cVar1S0S85P037P013P048P055(0)='1' AND  A(10)='1' AND A(22)='0' )then
          cVar2S0S85P019P014nsss(0) <='1';
          else
          cVar2S0S85P019P014nsss(0) <='0';
          end if;
        if(cVar1S1S85P037P013P048P055(0)='1' AND  A(10)='0' AND A(23)='1' )then
          cVar2S1S85N019P012nsss(0) <='1';
          else
          cVar2S1S85N019P012nsss(0) <='0';
          end if;
        if(cVar1S2S85P037P013P048N055(0)='1' AND  E(19)='0' AND B(11)='0' AND B(23)='0' )then
          cVar2S2S85P057P035P030nsss(0) <='1';
          else
          cVar2S2S85P057P035P030nsss(0) <='0';
          end if;
        if(cVar1S3S85P037P013P048N055(0)='1' AND  E(19)='0' AND B(11)='1' AND D( 9)='1' )then
          cVar2S3S85P057P035P062nsss(0) <='1';
          else
          cVar2S3S85P057P035P062nsss(0) <='0';
          end if;
        if(cVar1S4S85P037P013P048N055(0)='1' AND  E(19)='1' AND A(20)='1' )then
          cVar2S4S85P057P018nsss(0) <='1';
          else
          cVar2S4S85P057P018nsss(0) <='0';
          end if;
        if(cVar1S5S85P037P013P048P035(0)='1' AND  D(13)='1' )then
          cVar2S5S85P046nsss(0) <='1';
          else
          cVar2S5S85P046nsss(0) <='0';
          end if;
        if(cVar1S6S85P037P013P018P050(0)='1' AND  A(11)='0' AND D( 8)='1' )then
          cVar2S6S85P017P066nsss(0) <='1';
          else
          cVar2S6S85P017P066nsss(0) <='0';
          end if;
        if(cVar1S7S85P037P013P018P050(0)='1' AND  A(11)='0' AND D( 8)='0' AND B(20)='1' )then
          cVar2S7S85P017N066P036nsss(0) <='1';
          else
          cVar2S7S85P017N066P036nsss(0) <='0';
          end if;
        if(cVar1S8S85P037P013P018P050(0)='1' AND  A(11)='1' AND A(12)='0' AND A(10)='0' )then
          cVar2S8S85P017P015P019nsss(0) <='1';
          else
          cVar2S8S85P017P015P019nsss(0) <='0';
          end if;
        if(cVar1S9S85P037P013P018P050(0)='1' AND  A(11)='1' AND A(12)='1' AND B(11)='1' )then
          cVar2S9S85P017P015P035nsss(0) <='1';
          else
          cVar2S9S85P017P015P035nsss(0) <='0';
          end if;
        if(cVar1S10S85P037P013N018P041(0)='1' AND  B(13)='1' )then
          cVar2S10S85P031nsss(0) <='1';
          else
          cVar2S10S85P031nsss(0) <='0';
          end if;
        if(cVar1S11S85P037P013N018P041(0)='1' AND  B(13)='0' AND A(23)='1' AND D( 8)='0' )then
          cVar2S11S85N031P012P066nsss(0) <='1';
          else
          cVar2S11S85N031P012P066nsss(0) <='0';
          end if;
        if(cVar1S13S85N037P058P011N031(0)='1' AND  B(12)='1' AND D( 9)='1' )then
          cVar2S13S85P033P062nsss(0) <='1';
          else
          cVar2S13S85P033P062nsss(0) <='0';
          end if;
        if(cVar1S14S85N037P058P011N031(0)='1' AND  B(12)='1' AND D( 9)='0' AND A(23)='0' )then
          cVar2S14S85P033N062P012nsss(0) <='1';
          else
          cVar2S14S85P033N062P012nsss(0) <='0';
          end if;
        if(cVar1S15S85N037P058P011N031(0)='1' AND  B(12)='0' AND A(24)='1' AND A(21)='0' )then
          cVar2S15S85N033P010P016nsss(0) <='1';
          else
          cVar2S15S85N033P010P016nsss(0) <='0';
          end if;
        if(cVar1S16S85N037P058P011N031(0)='1' AND  B(12)='0' AND A(24)='0' AND B(11)='1' )then
          cVar2S16S85N033N010P035nsss(0) <='1';
          else
          cVar2S16S85N033N010P035nsss(0) <='0';
          end if;
        if(cVar1S17S85N037P058P011P009(0)='1' AND  A(13)='0' AND A(11)='1' )then
          cVar2S17S85P013P017nsss(0) <='1';
          else
          cVar2S17S85P013P017nsss(0) <='0';
          end if;
        if(cVar1S18S85N037P058P011P009(0)='1' AND  A(13)='0' AND A(11)='0' AND A(22)='1' )then
          cVar2S18S85P013N017P014nsss(0) <='1';
          else
          cVar2S18S85P013N017P014nsss(0) <='0';
          end if;
        if(cVar1S20S85N037N058P021N040(0)='1' AND  E(18)='0' AND E( 9)='1' )then
          cVar2S20S85P061P064nsss(0) <='1';
          else
          cVar2S20S85P061P064nsss(0) <='0';
          end if;
        if(cVar1S21S85N037N058P021N040(0)='1' AND  E(18)='0' AND E( 9)='0' AND A(14)='0' )then
          cVar2S21S85P061N064P011nsss(0) <='1';
          else
          cVar2S21S85P061N064P011nsss(0) <='0';
          end if;
        if(cVar1S22S85N037N058N021P048(0)='1' AND  B(16)='1' )then
          cVar2S22S85P025nsss(0) <='1';
          else
          cVar2S22S85P025nsss(0) <='0';
          end if;
        if(cVar1S23S85N037N058N021P048(0)='1' AND  B(16)='0' AND B(15)='1' )then
          cVar2S23S85N025P027nsss(0) <='1';
          else
          cVar2S23S85N025P027nsss(0) <='0';
          end if;
        if(cVar1S24S85N037N058N021P048(0)='1' AND  B(16)='0' AND B(15)='0' AND B(25)='1' )then
          cVar2S24S85N025N027P026nsss(0) <='1';
          else
          cVar2S24S85N025N027P026nsss(0) <='0';
          end if;
        if(cVar1S25S85N037N058N021N048(0)='1' AND  D(13)='0' AND B(28)='1' AND D(23)='1' )then
          cVar2S25S85P046P020P039nsss(0) <='1';
          else
          cVar2S25S85P046P020P039nsss(0) <='0';
          end if;
        if(cVar1S1S86P037P048N025P050(0)='1' AND  B(15)='1' )then
          cVar2S1S86P027nsss(0) <='1';
          else
          cVar2S1S86P027nsss(0) <='0';
          end if;
        if(cVar1S2S86P037P048N025P050(0)='1' AND  B(15)='0' AND A(23)='0' )then
          cVar2S2S86N027P012nsss(0) <='1';
          else
          cVar2S2S86N027P012nsss(0) <='0';
          end if;
        if(cVar1S3S86P037P048N025N050(0)='1' AND  D(21)='1' )then
          cVar2S3S86P047nsss(0) <='1';
          else
          cVar2S3S86P047nsss(0) <='0';
          end if;
        if(cVar1S4S86P037P048N025N050(0)='1' AND  D(21)='0' AND D( 9)='1' )then
          cVar2S4S86N047P062nsss(0) <='1';
          else
          cVar2S4S86N047P062nsss(0) <='0';
          end if;
        if(cVar1S5S86P037N048P046P036(0)='1' AND  B(22)='0' AND E(11)='1' )then
          cVar2S5S86P032P056nsss(0) <='1';
          else
          cVar2S5S86P032P056nsss(0) <='0';
          end if;
        if(cVar1S6S86P037N048P046P036(0)='1' AND  B(22)='0' AND E(11)='0' AND A(19)='0' )then
          cVar2S6S86P032N056P001nsss(0) <='1';
          else
          cVar2S6S86P032N056P001nsss(0) <='0';
          end if;
        if(cVar1S7S86P037N048P046P036(0)='1' AND  B(22)='1' AND E(16)='1' AND A(12)='1' )then
          cVar2S7S86P032P069P015nsss(0) <='1';
          else
          cVar2S7S86P032P069P015nsss(0) <='0';
          end if;
        if(cVar1S8S86P037N048P046N036(0)='1' AND  A(15)='0' AND A(10)='1' AND E(14)='0' )then
          cVar2S8S86P009P019P044nsss(0) <='1';
          else
          cVar2S8S86P009P019P044nsss(0) <='0';
          end if;
        if(cVar1S9S86P037N048P046N036(0)='1' AND  A(15)='0' AND A(10)='0' )then
          cVar2S9S86P009N019psss(0) <='1';
          else
          cVar2S9S86P009N019psss(0) <='0';
          end if;
        if(cVar1S10S86P037N048P046N036(0)='1' AND  A(15)='1' AND A(21)='1' AND A(10)='0' )then
          cVar2S10S86P009P016P019nsss(0) <='1';
          else
          cVar2S10S86P009P016P019nsss(0) <='0';
          end if;
        if(cVar1S11S86P037N048P046P062(0)='1' AND  A(10)='0' AND A(20)='1' )then
          cVar2S11S86P019P018nsss(0) <='1';
          else
          cVar2S11S86P019P018nsss(0) <='0';
          end if;
        if(cVar1S12S86P037N048P046P062(0)='1' AND  A(10)='0' AND A(20)='0' AND E(14)='1' )then
          cVar2S12S86P019N018P044nsss(0) <='1';
          else
          cVar2S12S86P019N018P044nsss(0) <='0';
          end if;
        if(cVar1S13S86P037P004P031P035(0)='1' AND  A(22)='0' )then
          cVar2S13S86P014nsss(0) <='1';
          else
          cVar2S13S86P014nsss(0) <='0';
          end if;
        if(cVar1S14S86P037P004N031P055(0)='1' AND  A(10)='1' AND A(22)='0' )then
          cVar2S14S86P019P014nsss(0) <='1';
          else
          cVar2S14S86P019P014nsss(0) <='0';
          end if;
        if(cVar1S15S86P037P004N031P055(0)='1' AND  A(10)='0' AND E(19)='1' )then
          cVar2S15S86N019P057nsss(0) <='1';
          else
          cVar2S15S86N019P057nsss(0) <='0';
          end if;
        if(cVar1S16S86P037P004N031N055(0)='1' AND  E(19)='0' AND A(22)='1' )then
          cVar2S16S86P057P014nsss(0) <='1';
          else
          cVar2S16S86P057P014nsss(0) <='0';
          end if;
        if(cVar1S17S86P037P004N031N055(0)='1' AND  E(19)='0' AND A(22)='0' AND D(20)='1' )then
          cVar2S17S86P057N014P051nsss(0) <='1';
          else
          cVar2S17S86P057N014P051nsss(0) <='0';
          end if;
        if(cVar1S18S86P037P004P051P036(0)='1' AND  D( 8)='0' AND A(11)='0' )then
          cVar2S18S86P066P017nsss(0) <='1';
          else
          cVar2S18S86P066P017nsss(0) <='0';
          end if;
        if(cVar1S19S86P037P004P051P036(0)='1' AND  D( 8)='1' AND D( 9)='0' AND A(11)='1' )then
          cVar2S19S86P066P062P017nsss(0) <='1';
          else
          cVar2S19S86P066P062P017nsss(0) <='0';
          end if;
        if(cVar1S0S87P019P017P035P026(0)='1' AND  A(21)='1' AND E( 9)='1' )then
          cVar2S0S87P016P064nsss(0) <='1';
          else
          cVar2S0S87P016P064nsss(0) <='0';
          end if;
        if(cVar1S1S87P019P017P035P026(0)='1' AND  A(21)='1' AND E( 9)='0' AND B(20)='0' )then
          cVar2S1S87P016N064P036nsss(0) <='1';
          else
          cVar2S1S87P016N064P036nsss(0) <='0';
          end if;
        if(cVar1S2S87P019P017P035P026(0)='1' AND  A(21)='0' AND A(14)='1' )then
          cVar2S2S87N016P011nsss(0) <='1';
          else
          cVar2S2S87N016P011nsss(0) <='0';
          end if;
        if(cVar1S3S87P019P017P035P026(0)='1' AND  A(21)='0' AND A(14)='0' AND A(22)='1' )then
          cVar2S3S87N016N011P014nsss(0) <='1';
          else
          cVar2S3S87N016N011P014nsss(0) <='0';
          end if;
        if(cVar1S4S87P019P017N035P066(0)='1' AND  B(20)='1' AND A(24)='0' AND A(15)='0' )then
          cVar2S4S87P036P010P009nsss(0) <='1';
          else
          cVar2S4S87P036P010P009nsss(0) <='0';
          end if;
        if(cVar1S5S87P019P017N035P066(0)='1' AND  B(20)='0' AND D(16)='1' AND B(21)='0' )then
          cVar2S5S87N036P067P034nsss(0) <='1';
          else
          cVar2S5S87N036P067P034nsss(0) <='0';
          end if;
        if(cVar1S6S87P019P017N035P066(0)='1' AND  B(20)='0' AND D(16)='0' AND E(10)='1' )then
          cVar2S6S87N036N067P060nsss(0) <='1';
          else
          cVar2S6S87N036N067P060nsss(0) <='0';
          end if;
        if(cVar1S7S87P019P017N035N066(0)='1' AND  B(12)='0' AND E(22)='1' AND A(22)='0' )then
          cVar2S7S87P033P045P014nsss(0) <='1';
          else
          cVar2S7S87P033P045P014nsss(0) <='0';
          end if;
        if(cVar1S8S87P019P017N035N066(0)='1' AND  B(12)='0' AND E(22)='0' AND D(22)='0' )then
          cVar2S8S87P033N045P043nsss(0) <='1';
          else
          cVar2S8S87P033N045P043nsss(0) <='0';
          end if;
        if(cVar1S9S87P019P017N035N066(0)='1' AND  B(12)='1' AND A(23)='0' AND A(12)='1' )then
          cVar2S9S87P033P012P015nsss(0) <='1';
          else
          cVar2S9S87P033P012P015nsss(0) <='0';
          end if;
        if(cVar1S10S87P019P017P053P029(0)='1' AND  B(11)='0' AND B(13)='1' AND A(12)='0' )then
          cVar2S10S87P035P031P015nsss(0) <='1';
          else
          cVar2S10S87P035P031P015nsss(0) <='0';
          end if;
        if(cVar1S11S87P019P017P053P029(0)='1' AND  B(11)='1' AND B(22)='0' AND D(17)='1' )then
          cVar2S11S87P035P032P063nsss(0) <='1';
          else
          cVar2S11S87P035P032P063nsss(0) <='0';
          end if;
        if(cVar1S12S87P019P017P053P029(0)='1' AND  A(14)='1' )then
          cVar2S12S87P011nsss(0) <='1';
          else
          cVar2S12S87P011nsss(0) <='0';
          end if;
        if(cVar1S13S87P019P017P053P037(0)='1' AND  A(22)='0' )then
          cVar2S13S87P014nsss(0) <='1';
          else
          cVar2S13S87P014nsss(0) <='0';
          end if;
        if(cVar1S14S87N019P009P068P039(0)='1' AND  B(21)='1' AND B(11)='0' )then
          cVar2S14S87P034P035nsss(0) <='1';
          else
          cVar2S14S87P034P035nsss(0) <='0';
          end if;
        if(cVar1S15S87N019P009P068P039(0)='1' AND  B(21)='0' AND A(26)='1' AND A(14)='0' )then
          cVar2S15S87N034P006P011nsss(0) <='1';
          else
          cVar2S15S87N034P006P011nsss(0) <='0';
          end if;
        if(cVar1S16S87N019P009P068P039(0)='1' AND  B(21)='0' AND A(26)='0' AND B(15)='1' )then
          cVar2S16S87N034N006P027nsss(0) <='1';
          else
          cVar2S16S87N034N006P027nsss(0) <='0';
          end if;
        if(cVar1S19S87N019N009P040N021(0)='1' AND  B(28)='1' )then
          cVar2S19S87P020nsss(0) <='1';
          else
          cVar2S19S87P020nsss(0) <='0';
          end if;
        if(cVar1S20S87N019N009P040N021(0)='1' AND  B(28)='0' AND A(11)='1' AND A(20)='0' )then
          cVar2S20S87N020P017P018nsss(0) <='1';
          else
          cVar2S20S87N020P017P018nsss(0) <='0';
          end if;
        if(cVar1S21S87N019N009P040N021(0)='1' AND  B(28)='0' AND A(11)='0' AND A(20)='1' )then
          cVar2S21S87N020N017P018nsss(0) <='1';
          else
          cVar2S21S87N020N017P018nsss(0) <='0';
          end if;
        if(cVar1S22S87N019N009N040P038(0)='1' AND  B(18)='0' AND E( 8)='1' AND D(21)='0' )then
          cVar2S22S87P021P068P047nsss(0) <='1';
          else
          cVar2S22S87P021P068P047nsss(0) <='0';
          end if;
        if(cVar1S23S87N019N009N040P038(0)='1' AND  B(18)='0' AND E( 8)='0' AND E(10)='1' )then
          cVar2S23S87P021N068P060nsss(0) <='1';
          else
          cVar2S23S87P021N068P060nsss(0) <='0';
          end if;
        if(cVar1S24S87N019N009N040P038(0)='1' AND  B(18)='1' AND D(23)='1' )then
          cVar2S24S87P021P039nsss(0) <='1';
          else
          cVar2S24S87P021P039nsss(0) <='0';
          end if;
        if(cVar1S25S87N019N009N040P038(0)='1' AND  A(12)='1' )then
          cVar2S25S87P015nsss(0) <='1';
          else
          cVar2S25S87P015nsss(0) <='0';
          end if;
        if(cVar1S0S88P060P009P068P063(0)='1' AND  A(16)='1' AND A(17)='0' AND A(13)='0' )then
          cVar2S0S88P007P005P013nsss(0) <='1';
          else
          cVar2S0S88P007P005P013nsss(0) <='0';
          end if;
        if(cVar1S1S88P060P009P068P063(0)='1' AND  A(16)='0' AND A(23)='0' )then
          cVar2S1S88N007P012nsss(0) <='1';
          else
          cVar2S1S88N007P012nsss(0) <='0';
          end if;
        if(cVar1S2S88P060P009P068P063(0)='1' AND  A(16)='0' AND A(23)='1' AND A(13)='1' )then
          cVar2S2S88N007P012P013nsss(0) <='1';
          else
          cVar2S2S88N007P012P013nsss(0) <='0';
          end if;
        if(cVar1S3S88P060P009P068P063(0)='1' AND  A(25)='0' AND A(21)='1' AND A(23)='0' )then
          cVar2S3S88P008P016P012nsss(0) <='1';
          else
          cVar2S3S88P008P016P012nsss(0) <='0';
          end if;
        if(cVar1S4S88P060P009P068P063(0)='1' AND  A(25)='0' AND A(21)='0' AND B(20)='1' )then
          cVar2S4S88P008N016P036nsss(0) <='1';
          else
          cVar2S4S88P008N016P036nsss(0) <='0';
          end if;
        if(cVar1S5S88P060P009P068P002(0)='1' AND  D(18)='1' AND A(20)='1' )then
          cVar2S5S88P059P018nsss(0) <='1';
          else
          cVar2S5S88P059P018nsss(0) <='0';
          end if;
        if(cVar1S6S88P060P009P068P002(0)='1' AND  D(18)='0' AND D( 8)='1' AND D( 9)='1' )then
          cVar2S6S88N059P066P062nsss(0) <='1';
          else
          cVar2S6S88N059P066P062nsss(0) <='0';
          end if;
        if(cVar1S7S88P060N009P053P055(0)='1' AND  A(16)='0' )then
          cVar2S7S88P007nsss(0) <='1';
          else
          cVar2S7S88P007nsss(0) <='0';
          end if;
        if(cVar1S8S88P060N009P053N055(0)='1' AND  D(10)='0' AND B(24)='0' AND E(12)='0' )then
          cVar2S8S88P058P028P052nsss(0) <='1';
          else
          cVar2S8S88P058P028P052nsss(0) <='0';
          end if;
        if(cVar1S9S88P060N009P053N055(0)='1' AND  D(10)='0' AND B(24)='1' AND D(11)='1' )then
          cVar2S9S88P058P028P054nsss(0) <='1';
          else
          cVar2S9S88P058P028P054nsss(0) <='0';
          end if;
        if(cVar1S10S88P060N009P053N055(0)='1' AND  D(10)='1' AND B(10)='0' AND E(12)='1' )then
          cVar2S10S88P058P037P052nsss(0) <='1';
          else
          cVar2S10S88P058P037P052nsss(0) <='0';
          end if;
        if(cVar1S12S88P060N009P053N028(0)='1' AND  A(25)='1' AND B(25)='1' )then
          cVar2S12S88P008P026nsss(0) <='1';
          else
          cVar2S12S88P008P026nsss(0) <='0';
          end if;
        if(cVar1S13S88P060N009P053N028(0)='1' AND  A(25)='0' AND B(14)='1' )then
          cVar2S13S88N008P029nsss(0) <='1';
          else
          cVar2S13S88N008P029nsss(0) <='0';
          end if;
        if(cVar1S14S88P060N009P053N028(0)='1' AND  A(25)='0' AND B(14)='0' AND E(13)='1' )then
          cVar2S14S88N008N029P048nsss(0) <='1';
          else
          cVar2S14S88N008N029P048nsss(0) <='0';
          end if;
        if(cVar1S15S88P060P039P062P051(0)='1' AND  B(21)='1' )then
          cVar2S15S88P034nsss(0) <='1';
          else
          cVar2S15S88P034nsss(0) <='0';
          end if;
        if(cVar1S16S88P060P039P062P051(0)='1' AND  B(21)='0' AND A(15)='0' AND A(21)='0' )then
          cVar2S16S88N034P009P016nsss(0) <='1';
          else
          cVar2S16S88N034P009P016nsss(0) <='0';
          end if;
        if(cVar1S17S88P060P039N062P031(0)='1' AND  A(23)='1' )then
          cVar2S17S88P012nsss(0) <='1';
          else
          cVar2S17S88P012nsss(0) <='0';
          end if;
        if(cVar1S18S88P060P039N062P031(0)='1' AND  A(23)='0' AND A(13)='1' )then
          cVar2S18S88N012P013nsss(0) <='1';
          else
          cVar2S18S88N012P013nsss(0) <='0';
          end if;
        if(cVar1S19S88P060P039N062N031(0)='1' AND  E(16)='1' AND A(22)='0' )then
          cVar2S19S88P069P014nsss(0) <='1';
          else
          cVar2S19S88P069P014nsss(0) <='0';
          end if;
        if(cVar1S20S88P060P039N062N031(0)='1' AND  E(16)='0' AND E(17)='0' AND D( 8)='1' )then
          cVar2S20S88N069P065P066nsss(0) <='1';
          else
          cVar2S20S88N069P065P066nsss(0) <='0';
          end if;
        if(cVar1S0S89P009P068P063P007(0)='1' AND  A(17)='0' AND A(13)='0' )then
          cVar2S0S89P005P013nsss(0) <='1';
          else
          cVar2S0S89P005P013nsss(0) <='0';
          end if;
        if(cVar1S1S89P009P068P063P007(0)='1' AND  A(17)='0' AND A(13)='1' AND A(10)='0' )then
          cVar2S1S89P005P013P019nsss(0) <='1';
          else
          cVar2S1S89P005P013P019nsss(0) <='0';
          end if;
        if(cVar1S2S89P009P068P063N007(0)='1' AND  B(23)='0' AND A(23)='0' )then
          cVar2S2S89P030P012nsss(0) <='1';
          else
          cVar2S2S89P030P012nsss(0) <='0';
          end if;
        if(cVar1S3S89P009P068P063P008(0)='1' AND  D( 8)='0' AND A(21)='1' )then
          cVar2S3S89P066P016nsss(0) <='1';
          else
          cVar2S3S89P066P016nsss(0) <='0';
          end if;
        if(cVar1S5S89P009P068P002N047(0)='1' AND  D(18)='1' AND A(11)='0' )then
          cVar2S5S89P059P017nsss(0) <='1';
          else
          cVar2S5S89P059P017nsss(0) <='0';
          end if;
        if(cVar1S6S89P009P068P002N047(0)='1' AND  D(18)='0' AND D( 8)='1' AND D(12)='1' )then
          cVar2S6S89N059P066P050nsss(0) <='1';
          else
          cVar2S6S89N059P066P050nsss(0) <='0';
          end if;
        if(cVar1S8S89N009P049P023N005(0)='1' AND  D(14)='1' )then
          cVar2S8S89P042nsss(0) <='1';
          else
          cVar2S8S89P042nsss(0) <='0';
          end if;
        if(cVar1S9S89N009P049P023N005(0)='1' AND  D(14)='0' AND A(16)='1' )then
          cVar2S9S89N042P007nsss(0) <='1';
          else
          cVar2S9S89N042P007nsss(0) <='0';
          end if;
        if(cVar1S10S89N009P049P023N005(0)='1' AND  D(14)='0' AND A(16)='0' AND B(20)='1' )then
          cVar2S10S89N042N007P036nsss(0) <='1';
          else
          cVar2S10S89N042N007P036nsss(0) <='0';
          end if;
        if(cVar1S11S89N009P049N023P043(0)='1' AND  B(27)='0' AND E(22)='1' AND A(23)='1' )then
          cVar2S11S89P022P045P012nsss(0) <='1';
          else
          cVar2S11S89P022P045P012nsss(0) <='0';
          end if;
        if(cVar1S12S89N009P049N023P043(0)='1' AND  B(27)='1' AND A(22)='0' AND D(14)='1' )then
          cVar2S12S89P022P014P042nsss(0) <='1';
          else
          cVar2S12S89P022P014P042nsss(0) <='0';
          end if;
        if(cVar1S13S89N009P049N023P043(0)='1' AND  B(27)='1' )then
          cVar2S13S89P022nsss(0) <='1';
          else
          cVar2S13S89P022nsss(0) <='0';
          end if;
        if(cVar1S14S89N009P049N023P043(0)='1' AND  B(27)='0' AND B(26)='1' AND E(22)='1' )then
          cVar2S14S89N022P024P045nsss(0) <='1';
          else
          cVar2S14S89N022P024P045nsss(0) <='0';
          end if;
        if(cVar1S15S89N009P049N023P043(0)='1' AND  B(27)='0' AND B(26)='0' AND A(16)='1' )then
          cVar2S15S89N022N024P007nsss(0) <='1';
          else
          cVar2S15S89N022N024P007nsss(0) <='0';
          end if;
        if(cVar1S17S89N009P049N026P024(0)='1' AND  D(21)='1' )then
          cVar2S17S89P047nsss(0) <='1';
          else
          cVar2S17S89P047nsss(0) <='0';
          end if;
        if(cVar1S18S89N009P049N026N024(0)='1' AND  D(13)='1' )then
          cVar2S18S89P046nsss(0) <='1';
          else
          cVar2S18S89P046nsss(0) <='0';
          end if;
        if(cVar1S19S89N009P049N026N024(0)='1' AND  D(13)='0' AND A(17)='1' )then
          cVar2S19S89N046P005nsss(0) <='1';
          else
          cVar2S19S89N046P005nsss(0) <='0';
          end if;
        if(cVar1S20S89N009P049N026N024(0)='1' AND  D(13)='0' AND A(17)='0' AND A(16)='1' )then
          cVar2S20S89N046N005P007nsss(0) <='1';
          else
          cVar2S20S89N046N005P007nsss(0) <='0';
          end if;
        if(cVar1S1S90P049P052N065P062(0)='1' AND  B(11)='0' )then
          cVar2S1S90P035nsss(0) <='1';
          else
          cVar2S1S90P035nsss(0) <='0';
          end if;
        if(cVar1S2S90P049P052N065N062(0)='1' AND  D(12)='1' AND A(20)='0' AND A(21)='0' )then
          cVar2S2S90P050P018P016nsss(0) <='1';
          else
          cVar2S2S90P050P018P016nsss(0) <='0';
          end if;
        if(cVar1S3S90P049P052N065N062(0)='1' AND  D(12)='1' AND A(20)='1' AND B(14)='1' )then
          cVar2S3S90P050P018P029nsss(0) <='1';
          else
          cVar2S3S90P050P018P029nsss(0) <='0';
          end if;
        if(cVar1S4S90P049P052N065N062(0)='1' AND  D(12)='0' AND D( 8)='1' )then
          cVar2S4S90N050P066nsss(0) <='1';
          else
          cVar2S4S90N050P066nsss(0) <='0';
          end if;
        if(cVar1S5S90P049P052N065N062(0)='1' AND  D(12)='0' AND D( 8)='0' AND A(13)='1' )then
          cVar2S5S90N050N066P013nsss(0) <='1';
          else
          cVar2S5S90N050N066P013nsss(0) <='0';
          end if;
        if(cVar1S6S90P049N052P029P055(0)='1' AND  B(25)='0' AND A(24)='1' AND E(19)='1' )then
          cVar2S6S90P026P010P057nsss(0) <='1';
          else
          cVar2S6S90P026P010P057nsss(0) <='0';
          end if;
        if(cVar1S7S90P049N052P029P055(0)='1' AND  B(25)='0' AND A(24)='0' AND A(26)='0' )then
          cVar2S7S90P026N010P006nsss(0) <='1';
          else
          cVar2S7S90P026N010P006nsss(0) <='0';
          end if;
        if(cVar1S8S90P049N052P029N055(0)='1' AND  D(22)='0' AND B(27)='0' AND E(22)='0' )then
          cVar2S8S90P043P022P045nsss(0) <='1';
          else
          cVar2S8S90P043P022P045nsss(0) <='0';
          end if;
        if(cVar1S9S90P049N052P029N055(0)='1' AND  D(22)='0' AND B(27)='1' AND A(28)='1' )then
          cVar2S9S90P043P022P002nsss(0) <='1';
          else
          cVar2S9S90P043P022P002nsss(0) <='0';
          end if;
        if(cVar1S10S90P049N052P029N055(0)='1' AND  D(22)='1' AND B(27)='1' )then
          cVar2S10S90P043P022nsss(0) <='1';
          else
          cVar2S10S90P043P022nsss(0) <='0';
          end if;
        if(cVar1S11S90P049N052P029N055(0)='1' AND  D(22)='1' AND B(27)='0' AND B(17)='1' )then
          cVar2S11S90P043N022P023nsss(0) <='1';
          else
          cVar2S11S90P043N022P023nsss(0) <='0';
          end if;
        if(cVar1S12S90P049N052P029P056(0)='1' AND  A(10)='0' )then
          cVar2S12S90P019nsss(0) <='1';
          else
          cVar2S12S90P019nsss(0) <='0';
          end if;
        if(cVar1S13S90P049N052P029N056(0)='1' AND  D(20)='1' )then
          cVar2S13S90P051nsss(0) <='1';
          else
          cVar2S13S90P051nsss(0) <='0';
          end if;
        if(cVar1S16S90P049N026N027P024(0)='1' AND  D(21)='1' )then
          cVar2S16S90P047nsss(0) <='1';
          else
          cVar2S16S90P047nsss(0) <='0';
          end if;
        if(cVar1S17S90P049N026N027N024(0)='1' AND  D(13)='1' )then
          cVar2S17S90P046nsss(0) <='1';
          else
          cVar2S17S90P046nsss(0) <='0';
          end if;
        if(cVar1S18S90P049N026N027N024(0)='1' AND  D(13)='0' AND A(21)='1' AND D(20)='0' )then
          cVar2S18S90N046P016P051nsss(0) <='1';
          else
          cVar2S18S90N046P016P051nsss(0) <='0';
          end if;
        if(cVar1S19S90P049N026N027N024(0)='1' AND  D(13)='0' AND A(21)='0' AND A(17)='1' )then
          cVar2S19S90N046N016P005nsss(0) <='1';
          else
          cVar2S19S90N046N016P005nsss(0) <='0';
          end if;
        if(cVar1S2S91P052N065N062P050(0)='1' AND  B(21)='0' AND A(21)='0' )then
          cVar2S2S91P034P016nsss(0) <='1';
          else
          cVar2S2S91P034P016nsss(0) <='0';
          end if;
        if(cVar1S3S91P052N065N062P050(0)='1' AND  B(21)='0' AND A(21)='1' AND A(12)='1' )then
          cVar2S3S91P034P016P015nsss(0) <='1';
          else
          cVar2S3S91P034P016P015nsss(0) <='0';
          end if;
        if(cVar1S4S91P052N065N062N050(0)='1' AND  D(16)='1' )then
          cVar2S4S91P067nsss(0) <='1';
          else
          cVar2S4S91P067nsss(0) <='0';
          end if;
        if(cVar1S5S91P052N065N062N050(0)='1' AND  D(16)='0' AND D( 8)='1' )then
          cVar2S5S91N067P066nsss(0) <='1';
          else
          cVar2S5S91N067P066nsss(0) <='0';
          end if;
        if(cVar1S6S91P052N065N062N050(0)='1' AND  D(16)='0' AND D( 8)='0' AND A(13)='1' )then
          cVar2S6S91N067N066P013nsss(0) <='1';
          else
          cVar2S6S91N067N066P013nsss(0) <='0';
          end if;
        if(cVar1S7S91N052P048P061P007(0)='1' AND  B(16)='1' )then
          cVar2S7S91P025nsss(0) <='1';
          else
          cVar2S7S91P025nsss(0) <='0';
          end if;
        if(cVar1S8S91N052P048P061P007(0)='1' AND  B(16)='0' AND A(20)='1' )then
          cVar2S8S91N025P018nsss(0) <='1';
          else
          cVar2S8S91N025P018nsss(0) <='0';
          end if;
        if(cVar1S9S91N052P048P061N007(0)='1' AND  B(10)='0' AND D( 9)='1' )then
          cVar2S9S91P037P062nsss(0) <='1';
          else
          cVar2S9S91P037P062nsss(0) <='0';
          end if;
        if(cVar1S10S91N052P048P061N007(0)='1' AND  B(10)='0' AND D( 9)='0' AND D(16)='1' )then
          cVar2S10S91P037N062P067nsss(0) <='1';
          else
          cVar2S10S91P037N062P067nsss(0) <='0';
          end if;
        if(cVar1S11S91N052P048P061N007(0)='1' AND  B(10)='1' AND A(20)='0' AND D( 8)='0' )then
          cVar2S11S91P037P018P066nsss(0) <='1';
          else
          cVar2S11S91P037P018P066nsss(0) <='0';
          end if;
        if(cVar1S13S91N052N048P050P055(0)='1' AND  B(25)='0' AND A(27)='0' )then
          cVar2S13S91P026P004nsss(0) <='1';
          else
          cVar2S13S91P026P004nsss(0) <='0';
          end if;
        if(cVar1S14S91N052N048P050N055(0)='1' AND  E(19)='0' AND E(15)='1' AND B(18)='1' )then
          cVar2S14S91P057P040P021nsss(0) <='1';
          else
          cVar2S14S91P057P040P021nsss(0) <='0';
          end if;
        if(cVar1S15S91N052N048P050P004(0)='1' AND  E(17)='0' AND A(19)='0' AND A(21)='1' )then
          cVar2S15S91P065P001P016nsss(0) <='1';
          else
          cVar2S15S91P065P001P016nsss(0) <='0';
          end if;
        if(cVar1S1S92P019P068P029N054(0)='1' AND  D(20)='1' )then
          cVar2S1S92P051nsss(0) <='1';
          else
          cVar2S1S92P051nsss(0) <='0';
          end if;
        if(cVar1S2S92P019P068P029N054(0)='1' AND  D(20)='0' AND E(12)='1' )then
          cVar2S2S92N051P052nsss(0) <='1';
          else
          cVar2S2S92N051P052nsss(0) <='0';
          end if;
        if(cVar1S3S92P019P068P029N054(0)='1' AND  D(20)='0' AND E(12)='0' AND A(12)='1' )then
          cVar2S3S92N051N052P015nsss(0) <='1';
          else
          cVar2S3S92N051N052P015nsss(0) <='0';
          end if;
        if(cVar1S4S92P019P068N029P054(0)='1' AND  B(10)='1' AND A(16)='0' AND A(18)='0' )then
          cVar2S4S92P037P007P003nsss(0) <='1';
          else
          cVar2S4S92P037P007P003nsss(0) <='0';
          end if;
        if(cVar1S5S92P019P068N029P054(0)='1' AND  B(10)='1' AND A(16)='1' AND A(15)='1' )then
          cVar2S5S92P037P007P009nsss(0) <='1';
          else
          cVar2S5S92P037P007P009nsss(0) <='0';
          end if;
        if(cVar1S6S92P019P068N029P054(0)='1' AND  B(10)='0' AND E(22)='1' )then
          cVar2S6S92N037P045nsss(0) <='1';
          else
          cVar2S6S92N037P045nsss(0) <='0';
          end if;
        if(cVar1S7S92P019P068N029P054(0)='1' AND  B(10)='0' AND E(22)='0' AND D(22)='0' )then
          cVar2S7S92N037N045P043nsss(0) <='1';
          else
          cVar2S7S92N037N045P043nsss(0) <='0';
          end if;
        if(cVar1S8S92P019P068N029P054(0)='1' AND  B(21)='1' )then
          cVar2S8S92P034nsss(0) <='1';
          else
          cVar2S8S92P034nsss(0) <='0';
          end if;
        if(cVar1S9S92P019P068N029P054(0)='1' AND  B(21)='0' AND B(25)='0' AND B(23)='1' )then
          cVar2S9S92N034P026P030nsss(0) <='1';
          else
          cVar2S9S92N034P026P030nsss(0) <='0';
          end if;
        if(cVar1S10S92P019P068P055P050(0)='1' AND  A(24)='0' )then
          cVar2S10S92P010nsss(0) <='1';
          else
          cVar2S10S92P010nsss(0) <='0';
          end if;
        if(cVar1S11S92P019P068P055N050(0)='1' AND  A(14)='0' AND B(14)='0' AND E(11)='1' )then
          cVar2S11S92P011P029P056nsss(0) <='1';
          else
          cVar2S11S92P011P029P056nsss(0) <='0';
          end if;
        if(cVar1S14S92P019P066P009N046(0)='1' AND  D(12)='0' AND E(18)='1' AND D(18)='1' )then
          cVar2S14S92P050P061P059nsss(0) <='1';
          else
          cVar2S14S92P050P061P059nsss(0) <='0';
          end if;
        if(cVar1S15S92P019P066P009N046(0)='1' AND  D(12)='0' AND E(18)='0' AND E(13)='0' )then
          cVar2S15S92P050N061P048nsss(0) <='1';
          else
          cVar2S15S92P050N061P048nsss(0) <='0';
          end if;
        if(cVar1S16S92P019P066P009N046(0)='1' AND  D(12)='1' AND E(12)='1' )then
          cVar2S16S92P050P052nsss(0) <='1';
          else
          cVar2S16S92P050P052nsss(0) <='0';
          end if;
        if(cVar1S17S92P019P066P009P068(0)='1' AND  A(27)='0' AND A(26)='1' )then
          cVar2S17S92P004P006nsss(0) <='1';
          else
          cVar2S17S92P004P006nsss(0) <='0';
          end if;
        if(cVar1S18S92P019P066P009P068(0)='1' AND  A(27)='0' AND A(26)='0' AND A(13)='1' )then
          cVar2S18S92P004N006P013nsss(0) <='1';
          else
          cVar2S18S92P004N006P013nsss(0) <='0';
          end if;
        if(cVar1S19S92P019N066P051P061(0)='1' AND  A(12)='1' AND A(14)='0' )then
          cVar2S19S92P015P011nsss(0) <='1';
          else
          cVar2S19S92P015P011nsss(0) <='0';
          end if;
        if(cVar1S20S92P019N066P051P061(0)='1' AND  A(12)='0' AND B(24)='1' AND A(20)='0' )then
          cVar2S20S92N015P028P018nsss(0) <='1';
          else
          cVar2S20S92N015P028P018nsss(0) <='0';
          end if;
        if(cVar1S21S92P019N066P051P061(0)='1' AND  A(12)='0' AND B(24)='0' AND E(13)='1' )then
          cVar2S21S92N015N028P048nsss(0) <='1';
          else
          cVar2S21S92N015N028P048nsss(0) <='0';
          end if;
        if(cVar1S22S92P019N066P051P061(0)='1' AND  D(10)='1' AND A(12)='0' )then
          cVar2S22S92P058P015nsss(0) <='1';
          else
          cVar2S22S92P058P015nsss(0) <='0';
          end if;
        if(cVar1S23S92P019N066P051P061(0)='1' AND  D(10)='0' AND D(16)='1' AND A(12)='0' )then
          cVar2S23S92N058P067P015nsss(0) <='1';
          else
          cVar2S23S92N058P067P015nsss(0) <='0';
          end if;
        if(cVar1S24S92P019N066P051P016(0)='1' AND  B(20)='0' AND D(17)='1' )then
          cVar2S24S92P036P063nsss(0) <='1';
          else
          cVar2S24S92P036P063nsss(0) <='0';
          end if;
        if(cVar1S25S92P019N066P051P016(0)='1' AND  B(20)='0' AND D(17)='0' AND A(25)='1' )then
          cVar2S25S92P036N063P008nsss(0) <='1';
          else
          cVar2S25S92P036N063P008nsss(0) <='0';
          end if;
        if(cVar1S26S92P019N066P051P016(0)='1' AND  A(13)='0' AND E(17)='0' AND A(22)='1' )then
          cVar2S26S92P013P065P014nsss(0) <='1';
          else
          cVar2S26S92P013P065P014nsss(0) <='0';
          end if;
        if(cVar1S0S93P019P051P002P000(0)='1' AND  A(23)='0' AND B(20)='1' )then
          cVar2S0S93P012P036nsss(0) <='1';
          else
          cVar2S0S93P012P036nsss(0) <='0';
          end if;
        if(cVar1S1S93P019P051P002P000(0)='1' AND  A(23)='0' AND B(20)='0' AND E(16)='0' )then
          cVar2S1S93P012N036P069nsss(0) <='1';
          else
          cVar2S1S93P012N036P069nsss(0) <='0';
          end if;
        if(cVar1S2S93P019P051P002P000(0)='1' AND  A(23)='1' AND A(24)='1' )then
          cVar2S2S93P012P010nsss(0) <='1';
          else
          cVar2S2S93P012P010nsss(0) <='0';
          end if;
        if(cVar1S3S93P019P051P002N000(0)='1' AND  E(16)='1' AND E(17)='1' AND D(18)='0' )then
          cVar2S3S93P069P065P059nsss(0) <='1';
          else
          cVar2S3S93P069P065P059nsss(0) <='0';
          end if;
        if(cVar1S4S93P019P051P002N000(0)='1' AND  E(16)='1' AND E(17)='0' AND B(23)='1' )then
          cVar2S4S93P069N065P030nsss(0) <='1';
          else
          cVar2S4S93P069N065P030nsss(0) <='0';
          end if;
        if(cVar1S5S93P019P051P002N000(0)='1' AND  E(16)='0' AND D(21)='1' )then
          cVar2S5S93N069P047nsss(0) <='1';
          else
          cVar2S5S93N069P047nsss(0) <='0';
          end if;
        if(cVar1S6S93P019P051P002N000(0)='1' AND  E(16)='0' AND D(21)='0' AND B(20)='0' )then
          cVar2S6S93N069N047P036nsss(0) <='1';
          else
          cVar2S6S93N069N047P036nsss(0) <='0';
          end if;
        if(cVar1S7S93P019P051P002P054(0)='1' AND  B(20)='1' AND A(24)='0' )then
          cVar2S7S93P036P010nsss(0) <='1';
          else
          cVar2S7S93P036P010nsss(0) <='0';
          end if;
        if(cVar1S8S93P019P051P024P037(0)='1' AND  D(16)='0' AND A(22)='0' )then
          cVar2S8S93P067P014nsss(0) <='1';
          else
          cVar2S8S93P067P014nsss(0) <='0';
          end if;
        if(cVar1S9S93P019P051P024N037(0)='1' AND  A(25)='1' AND A(13)='0' )then
          cVar2S9S93P008P013nsss(0) <='1';
          else
          cVar2S9S93P008P013nsss(0) <='0';
          end if;
        if(cVar1S10S93P019P051P024N037(0)='1' AND  A(25)='0' AND A(11)='0' AND A(13)='1' )then
          cVar2S10S93N008P017P013nsss(0) <='1';
          else
          cVar2S10S93N008P017P013nsss(0) <='0';
          end if;
        if(cVar1S12S93N019P056P054N013(0)='1' AND  A(21)='0' )then
          cVar2S12S93P016nsss(0) <='1';
          else
          cVar2S12S93P016nsss(0) <='0';
          end if;
        if(cVar1S13S93N019P056N054P058(0)='1' AND  A(23)='1' )then
          cVar2S13S93P012nsss(0) <='1';
          else
          cVar2S13S93P012nsss(0) <='0';
          end if;
        if(cVar1S14S93N019P056N054P058(0)='1' AND  A(23)='0' AND E(10)='0' )then
          cVar2S14S93N012P060nsss(0) <='1';
          else
          cVar2S14S93N012P060nsss(0) <='0';
          end if;
        if(cVar1S15S93N019P056N054N058(0)='1' AND  B(10)='0' AND A(11)='0' AND A(12)='1' )then
          cVar2S15S93P037P017P015nsss(0) <='1';
          else
          cVar2S15S93P037P017P015nsss(0) <='0';
          end if;
        if(cVar1S16S93N019N056P054P037(0)='1' AND  B(14)='0' AND B(24)='1' )then
          cVar2S16S93P029P028nsss(0) <='1';
          else
          cVar2S16S93P029P028nsss(0) <='0';
          end if;
        if(cVar1S17S93N019N056P054P037(0)='1' AND  B(14)='0' AND B(24)='0' AND A(18)='0' )then
          cVar2S17S93P029N028P003nsss(0) <='1';
          else
          cVar2S17S93P029N028P003nsss(0) <='0';
          end if;
        if(cVar1S18S93N019N056P054N037(0)='1' AND  A(16)='1' AND B(16)='1' )then
          cVar2S18S93P007P025nsss(0) <='1';
          else
          cVar2S18S93P007P025nsss(0) <='0';
          end if;
        if(cVar1S19S93N019N056P054N037(0)='1' AND  A(16)='1' AND B(16)='0' AND A(28)='1' )then
          cVar2S19S93P007N025P002nsss(0) <='1';
          else
          cVar2S19S93P007N025P002nsss(0) <='0';
          end if;
        if(cVar1S20S93N019N056P054N037(0)='1' AND  A(16)='0' AND E(20)='1' AND A(15)='1' )then
          cVar2S20S93N007P053P009nsss(0) <='1';
          else
          cVar2S20S93N007P053P009nsss(0) <='0';
          end if;
        if(cVar1S21S93N019N056P054P005(0)='1' AND  B(21)='1' )then
          cVar2S21S93P034nsss(0) <='1';
          else
          cVar2S21S93P034nsss(0) <='0';
          end if;
        if(cVar1S22S93N019N056P054P005(0)='1' AND  B(21)='0' AND D(17)='0' AND B(20)='1' )then
          cVar2S22S93N034P063P036nsss(0) <='1';
          else
          cVar2S22S93N034P063P036nsss(0) <='0';
          end if;
        if(cVar1S0S94P019P037P029P011(0)='1' AND  D(11)='1' )then
          cVar2S0S94P054nsss(0) <='1';
          else
          cVar2S0S94P054nsss(0) <='0';
          end if;
        if(cVar1S1S94P019P037P029P011(0)='1' AND  D(11)='0' AND D(20)='1' )then
          cVar2S1S94N054P051nsss(0) <='1';
          else
          cVar2S1S94N054P051nsss(0) <='0';
          end if;
        if(cVar1S2S94P019P037P029P011(0)='1' AND  D(11)='0' AND D(20)='0' AND E(12)='1' )then
          cVar2S2S94N054N051P052nsss(0) <='1';
          else
          cVar2S2S94N054N051P052nsss(0) <='0';
          end if;
        if(cVar1S3S94P019P037P029N011(0)='1' AND  B(21)='1' )then
          cVar2S3S94P034nsss(0) <='1';
          else
          cVar2S3S94P034nsss(0) <='0';
          end if;
        if(cVar1S4S94P019P037P029N011(0)='1' AND  B(21)='0' AND A(12)='1' )then
          cVar2S4S94N034P015nsss(0) <='1';
          else
          cVar2S4S94N034P015nsss(0) <='0';
          end if;
        if(cVar1S5S94P019P037P029N011(0)='1' AND  B(21)='0' AND A(12)='0' AND E(12)='1' )then
          cVar2S5S94N034N015P052nsss(0) <='1';
          else
          cVar2S5S94N034N015P052nsss(0) <='0';
          end if;
        if(cVar1S6S94P019P037N029P045(0)='1' AND  A(17)='1' )then
          cVar2S6S94P005nsss(0) <='1';
          else
          cVar2S6S94P005nsss(0) <='0';
          end if;
        if(cVar1S7S94P019P037N029P045(0)='1' AND  A(17)='0' AND B(26)='1' )then
          cVar2S7S94N005P024nsss(0) <='1';
          else
          cVar2S7S94N005P024nsss(0) <='0';
          end if;
        if(cVar1S8S94P019P037N029P045(0)='1' AND  A(17)='0' AND B(26)='0' AND A(16)='1' )then
          cVar2S8S94N005N024P007nsss(0) <='1';
          else
          cVar2S8S94N005N024P007nsss(0) <='0';
          end if;
        if(cVar1S9S94P019P037N029N045(0)='1' AND  B(27)='0' AND D(22)='0' )then
          cVar2S9S94P022P043nsss(0) <='1';
          else
          cVar2S9S94P022P043nsss(0) <='0';
          end if;
        if(cVar1S10S94P019P037N029N045(0)='1' AND  B(27)='0' AND D(22)='1' AND A(25)='1' )then
          cVar2S10S94P022P043P008nsss(0) <='1';
          else
          cVar2S10S94P022P043P008nsss(0) <='0';
          end if;
        if(cVar1S12S94P019P037P059N028(0)='1' AND  D(19)='0' AND A(25)='0' AND E(19)='0' )then
          cVar2S12S94P055P008P057nsss(0) <='1';
          else
          cVar2S12S94P055P008P057nsss(0) <='0';
          end if;
        if(cVar1S13S94P019P037P059P064(0)='1' AND  A(11)='1' )then
          cVar2S13S94P017nsss(0) <='1';
          else
          cVar2S13S94P017nsss(0) <='0';
          end if;
        if(cVar1S14S94P019P037P059P064(0)='1' AND  A(11)='0' AND E(18)='1' )then
          cVar2S14S94N017P061nsss(0) <='1';
          else
          cVar2S14S94N017P061nsss(0) <='0';
          end if;
        if(cVar1S15S94P019P069P051P029(0)='1' AND  D(14)='1' )then
          cVar2S15S94P042nsss(0) <='1';
          else
          cVar2S15S94P042nsss(0) <='0';
          end if;
        if(cVar1S16S94P019P069P051P029(0)='1' AND  D(14)='0' AND A(28)='0' )then
          cVar2S16S94N042P002nsss(0) <='1';
          else
          cVar2S16S94N042P002nsss(0) <='0';
          end if;
        if(cVar1S17S94P019P069P051P013(0)='1' AND  E(20)='1' )then
          cVar2S17S94P053nsss(0) <='1';
          else
          cVar2S17S94P053nsss(0) <='0';
          end if;
        if(cVar1S18S94P019N069P057P030(0)='1' AND  A(25)='1' AND D(17)='1' AND D( 8)='1' )then
          cVar2S18S94P008P063P066nsss(0) <='1';
          else
          cVar2S18S94P008P063P066nsss(0) <='0';
          end if;
        if(cVar1S19S94P019N069P057P030(0)='1' AND  A(25)='1' AND D(17)='0' AND B(22)='0' )then
          cVar2S19S94P008N063P032nsss(0) <='1';
          else
          cVar2S19S94P008N063P032nsss(0) <='0';
          end if;
        if(cVar1S20S94P019N069P057P030(0)='1' AND  A(25)='0' AND A(20)='1' AND E(18)='1' )then
          cVar2S20S94N008P018P061nsss(0) <='1';
          else
          cVar2S20S94N008P018P061nsss(0) <='0';
          end if;
        if(cVar1S21S94P019N069P057P061(0)='1' AND  A(20)='0' AND B(23)='1' )then
          cVar2S21S94P018P030nsss(0) <='1';
          else
          cVar2S21S94P018P030nsss(0) <='0';
          end if;
        if(cVar1S22S94P019N069P057P061(0)='1' AND  A(20)='0' AND B(23)='0' AND B(20)='0' )then
          cVar2S22S94P018N030P036nsss(0) <='1';
          else
          cVar2S22S94P018N030P036nsss(0) <='0';
          end if;
        if(cVar1S23S94P019N069P057P061(0)='1' AND  A(20)='1' AND E( 8)='0' AND D(19)='1' )then
          cVar2S23S94P018P068P055nsss(0) <='1';
          else
          cVar2S23S94P018P068P055nsss(0) <='0';
          end if;
        if(cVar1S0S95P019P057P036P009(0)='1' AND  D( 8)='0' AND A(23)='0' )then
          cVar2S0S95P066P012nsss(0) <='1';
          else
          cVar2S0S95P066P012nsss(0) <='0';
          end if;
        if(cVar1S1S95P019P057P036P009(0)='1' AND  D( 8)='0' AND A(23)='1' AND E(16)='0' )then
          cVar2S1S95P066P012P069nsss(0) <='1';
          else
          cVar2S1S95P066P012P069nsss(0) <='0';
          end if;
        if(cVar1S2S95P019P057P036P009(0)='1' AND  D( 8)='1' AND A(22)='1' )then
          cVar2S2S95P066P014nsss(0) <='1';
          else
          cVar2S2S95P066P014nsss(0) <='0';
          end if;
        if(cVar1S3S95P019P057P036N009(0)='1' AND  B(22)='0' AND A(27)='0' AND A(21)='1' )then
          cVar2S3S95P032P004P016nsss(0) <='1';
          else
          cVar2S3S95P032P004P016nsss(0) <='0';
          end if;
        if(cVar1S4S95P019P057P036N009(0)='1' AND  B(22)='1' AND A(23)='0' AND A(22)='1' )then
          cVar2S4S95P032P012P014nsss(0) <='1';
          else
          cVar2S4S95P032P012P014nsss(0) <='0';
          end if;
        if(cVar1S5S95P019P057N036P056(0)='1' AND  A(15)='0' AND A(27)='1' AND A(23)='0' )then
          cVar2S5S95P009P004P012nsss(0) <='1';
          else
          cVar2S5S95P009P004P012nsss(0) <='0';
          end if;
        if(cVar1S6S95P019P057N036P056(0)='1' AND  A(15)='0' AND A(27)='0' AND E(14)='0' )then
          cVar2S6S95P009N004P044nsss(0) <='1';
          else
          cVar2S6S95P009N004P044nsss(0) <='0';
          end if;
        if(cVar1S7S95P019P057N036P056(0)='1' AND  A(15)='1' AND A(11)='0' AND D(17)='0' )then
          cVar2S7S95P009P017P063nsss(0) <='1';
          else
          cVar2S7S95P009P017P063nsss(0) <='0';
          end if;
        if(cVar1S8S95P019P057N036P056(0)='1' AND  A(16)='1' )then
          cVar2S8S95P007nsss(0) <='1';
          else
          cVar2S8S95P007nsss(0) <='0';
          end if;
        if(cVar1S9S95P019P057N036P056(0)='1' AND  A(16)='0' AND A(24)='1' AND A(12)='0' )then
          cVar2S9S95N007P010P015nsss(0) <='1';
          else
          cVar2S9S95N007P010P015nsss(0) <='0';
          end if;
        if(cVar1S11S95P019P057P030N056(0)='1' AND  A(11)='0' AND E( 8)='0' )then
          cVar2S11S95P017P068nsss(0) <='1';
          else
          cVar2S11S95P017P068nsss(0) <='0';
          end if;
        if(cVar1S12S95P019P057N030P004(0)='1' AND  E(10)='0' AND A(22)='0' AND B(10)='1' )then
          cVar2S12S95P060P014P037nsss(0) <='1';
          else
          cVar2S12S95P060P014P037nsss(0) <='0';
          end if;
        if(cVar1S14S95N019P045P062N005(0)='1' AND  A(16)='1' )then
          cVar2S14S95P007nsss(0) <='1';
          else
          cVar2S14S95P007nsss(0) <='0';
          end if;
        if(cVar1S15S95N019P045P062N005(0)='1' AND  A(16)='0' AND E(16)='0' AND B(26)='1' )then
          cVar2S15S95N007P069P024nsss(0) <='1';
          else
          cVar2S15S95N007P069P024nsss(0) <='0';
          end if;
        if(cVar1S16S95N019N045P029P011(0)='1' AND  D(11)='1' )then
          cVar2S16S95P054nsss(0) <='1';
          else
          cVar2S16S95P054nsss(0) <='0';
          end if;
        if(cVar1S17S95N019N045P029P011(0)='1' AND  D(11)='0' AND D(20)='1' )then
          cVar2S17S95N054P051nsss(0) <='1';
          else
          cVar2S17S95N054P051nsss(0) <='0';
          end if;
        if(cVar1S18S95N019N045P029P011(0)='1' AND  D(11)='0' AND D(20)='0' AND E(12)='1' )then
          cVar2S18S95N054N051P052nsss(0) <='1';
          else
          cVar2S18S95N054N051P052nsss(0) <='0';
          end if;
        if(cVar1S19S95N019N045P029N011(0)='1' AND  D(19)='0' AND A(25)='1' )then
          cVar2S19S95P055P008nsss(0) <='1';
          else
          cVar2S19S95P055P008nsss(0) <='0';
          end if;
        if(cVar1S20S95N019N045P029N011(0)='1' AND  D(19)='0' AND A(25)='0' AND A(12)='1' )then
          cVar2S20S95P055N008P015nsss(0) <='1';
          else
          cVar2S20S95P055N008P015nsss(0) <='0';
          end if;
        if(cVar1S21S95N019N045N029P031(0)='1' AND  A(13)='1' AND A(14)='0' )then
          cVar2S21S95P013P011nsss(0) <='1';
          else
          cVar2S21S95P013P011nsss(0) <='0';
          end if;
        if(cVar1S22S95N019N045N029P031(0)='1' AND  A(13)='0' AND A(21)='0' AND A(23)='1' )then
          cVar2S22S95N013P016P012nsss(0) <='1';
          else
          cVar2S22S95N013P016P012nsss(0) <='0';
          end if;
        if(cVar1S23S95N019N045N029P031(0)='1' AND  A(13)='0' AND A(21)='1' AND A(23)='1' )then
          cVar2S23S95N013P016P012nsss(0) <='1';
          else
          cVar2S23S95N013P016P012nsss(0) <='0';
          end if;
        if(cVar1S24S95N019N045N029N031(0)='1' AND  D(11)='0' AND A(28)='1' AND B(25)='0' )then
          cVar2S24S95P054P002P026nsss(0) <='1';
          else
          cVar2S24S95P054P002P026nsss(0) <='0';
          end if;
        if(cVar1S25S95N019N045N029N031(0)='1' AND  D(11)='0' AND A(28)='0' AND B(24)='1' )then
          cVar2S25S95P054N002P028nsss(0) <='1';
          else
          cVar2S25S95P054N002P028nsss(0) <='0';
          end if;
        if(cVar1S26S95N019N045N029N031(0)='1' AND  D(11)='1' AND B(23)='1' )then
          cVar2S26S95P054P030nsss(0) <='1';
          else
          cVar2S26S95P054P030nsss(0) <='0';
          end if;
        if(cVar1S1S96P019P037P045N005(0)='1' AND  E(16)='0' AND B(26)='1' )then
          cVar2S1S96P069P024nsss(0) <='1';
          else
          cVar2S1S96P069P024nsss(0) <='0';
          end if;
        if(cVar1S2S96P019P037P045N005(0)='1' AND  E(16)='0' AND B(26)='0' AND A(14)='1' )then
          cVar2S2S96P069N024P011nsss(0) <='1';
          else
          cVar2S2S96P069N024P011nsss(0) <='0';
          end if;
        if(cVar1S3S96P019P037N045P029(0)='1' AND  A(14)='1' )then
          cVar2S3S96P011nsss(0) <='1';
          else
          cVar2S3S96P011nsss(0) <='0';
          end if;
        if(cVar1S4S96P019P037N045P029(0)='1' AND  A(14)='0' AND B(21)='1' )then
          cVar2S4S96N011P034nsss(0) <='1';
          else
          cVar2S4S96N011P034nsss(0) <='0';
          end if;
        if(cVar1S5S96P019P037N045P029(0)='1' AND  A(14)='0' AND B(21)='0' AND A(12)='1' )then
          cVar2S5S96N011N034P015nsss(0) <='1';
          else
          cVar2S5S96N011N034P015nsss(0) <='0';
          end if;
        if(cVar1S6S96P019P037N045N029(0)='1' AND  E(15)='1' AND D(15)='1' )then
          cVar2S6S96P040P038nsss(0) <='1';
          else
          cVar2S6S96P040P038nsss(0) <='0';
          end if;
        if(cVar1S7S96P019P037N045N029(0)='1' AND  E(15)='1' AND D(15)='0' AND D(14)='1' )then
          cVar2S7S96P040N038P042nsss(0) <='1';
          else
          cVar2S7S96P040N038P042nsss(0) <='0';
          end if;
        if(cVar1S8S96P019P037N045N029(0)='1' AND  E(15)='0' AND D(15)='0' AND B(27)='0' )then
          cVar2S8S96N040P038P022nsss(0) <='1';
          else
          cVar2S8S96N040P038P022nsss(0) <='0';
          end if;
        if(cVar1S10S96P019P037P059N028(0)='1' AND  E(21)='0' AND E( 9)='1' AND A(20)='1' )then
          cVar2S10S96P049P064P018nsss(0) <='1';
          else
          cVar2S10S96P049P064P018nsss(0) <='0';
          end if;
        if(cVar1S11S96P019P037P059N028(0)='1' AND  E(21)='0' AND E( 9)='0' AND E(23)='1' )then
          cVar2S11S96P049N064P041nsss(0) <='1';
          else
          cVar2S11S96P049N064P041nsss(0) <='0';
          end if;
        if(cVar1S12S96P019P037P059P064(0)='1' AND  A(11)='1' )then
          cVar2S12S96P017nsss(0) <='1';
          else
          cVar2S12S96P017nsss(0) <='0';
          end if;
        if(cVar1S13S96P019P037P059P064(0)='1' AND  A(11)='0' AND E(18)='1' )then
          cVar2S13S96N017P061nsss(0) <='1';
          else
          cVar2S13S96N017P061nsss(0) <='0';
          end if;
        if(cVar1S14S96P019P036P006P009(0)='1' AND  E(10)='0' AND B(21)='0' AND A(23)='0' )then
          cVar2S14S96P060P034P012nsss(0) <='1';
          else
          cVar2S14S96P060P034P012nsss(0) <='0';
          end if;
        if(cVar1S15S96P019P036P006N009(0)='1' AND  D(20)='0' AND E(11)='1' )then
          cVar2S15S96P051P056nsss(0) <='1';
          else
          cVar2S15S96P051P056nsss(0) <='0';
          end if;
        if(cVar1S16S96P019P036P006N009(0)='1' AND  D(20)='0' AND E(11)='0' AND A(14)='0' )then
          cVar2S16S96P051N056P011nsss(0) <='1';
          else
          cVar2S16S96P051N056P011nsss(0) <='0';
          end if;
        if(cVar1S17S96P019P036P006N009(0)='1' AND  D(20)='1' AND A(23)='0' AND A(21)='1' )then
          cVar2S17S96P051P012P016nsss(0) <='1';
          else
          cVar2S17S96P051P012P016nsss(0) <='0';
          end if;
        if(cVar1S18S96P019P036P006P004(0)='1' AND  B(21)='0' AND B(10)='1' )then
          cVar2S18S96P034P037nsss(0) <='1';
          else
          cVar2S18S96P034P037nsss(0) <='0';
          end if;
        if(cVar1S19S96P019P036P006P004(0)='1' AND  B(21)='0' AND B(10)='0' AND A(13)='1' )then
          cVar2S19S96P034N037P013nsss(0) <='1';
          else
          cVar2S19S96P034N037P013nsss(0) <='0';
          end if;
        if(cVar1S20S96P019N036P009P063(0)='1' AND  E( 9)='1' AND A(23)='1' )then
          cVar2S20S96P064P012nsss(0) <='1';
          else
          cVar2S20S96P064P012nsss(0) <='0';
          end if;
        if(cVar1S21S96P019N036P009P063(0)='1' AND  E( 9)='1' AND A(23)='0' AND E( 8)='1' )then
          cVar2S21S96P064N012P068nsss(0) <='1';
          else
          cVar2S21S96P064N012P068nsss(0) <='0';
          end if;
        if(cVar1S22S96P019N036P009P063(0)='1' AND  E( 9)='0' AND E(18)='0' AND D( 9)='0' )then
          cVar2S22S96N064P061P062nsss(0) <='1';
          else
          cVar2S22S96N064P061P062nsss(0) <='0';
          end if;
        if(cVar1S23S96P019N036P009N063(0)='1' AND  E(17)='0' AND B(13)='0' AND A(27)='1' )then
          cVar2S23S96P065P031P004nsss(0) <='1';
          else
          cVar2S23S96P065P031P004nsss(0) <='0';
          end if;
        if(cVar1S24S96P019N036P009N063(0)='1' AND  E(17)='0' AND B(13)='1' AND D(10)='1' )then
          cVar2S24S96P065P031P058nsss(0) <='1';
          else
          cVar2S24S96P065P031P058nsss(0) <='0';
          end if;
        if(cVar1S25S96P019N036P009N063(0)='1' AND  E(17)='1' AND B(21)='0' AND D( 8)='1' )then
          cVar2S25S96P065P034P066nsss(0) <='1';
          else
          cVar2S25S96P065P034P066nsss(0) <='0';
          end if;
        if(cVar1S26S96P019N036P009P028(0)='1' AND  B(28)='0' AND D(23)='1' )then
          cVar2S26S96P020P039nsss(0) <='1';
          else
          cVar2S26S96P020P039nsss(0) <='0';
          end if;
        if(cVar1S2S97P045P035N025N022(0)='1' AND  B(17)='1' )then
          cVar2S2S97P023nsss(0) <='1';
          else
          cVar2S2S97P023nsss(0) <='0';
          end if;
        if(cVar1S3S97P045P035N025N022(0)='1' AND  B(17)='0' AND B(26)='1' )then
          cVar2S3S97N023P024nsss(0) <='1';
          else
          cVar2S3S97N023P024nsss(0) <='0';
          end if;
        if(cVar1S4S97N045P043P019P023(0)='1' AND  A(27)='0' AND B(23)='1' AND B(13)='0' )then
          cVar2S4S97P004P030P031nsss(0) <='1';
          else
          cVar2S4S97P004P030P031nsss(0) <='0';
          end if;
        if(cVar1S5S97N045P043P019P023(0)='1' AND  A(27)='0' AND B(23)='0' AND E(19)='0' )then
          cVar2S5S97P004N030P057nsss(0) <='1';
          else
          cVar2S5S97P004N030P057nsss(0) <='0';
          end if;
        if(cVar1S6S97N045P043P019P023(0)='1' AND  A(23)='0' AND A(11)='0' )then
          cVar2S6S97P012P017nsss(0) <='1';
          else
          cVar2S6S97P012P017nsss(0) <='0';
          end if;
        if(cVar1S7S97N045P043N019P024(0)='1' AND  B(14)='1' AND A(14)='1' )then
          cVar2S7S97P029P011nsss(0) <='1';
          else
          cVar2S7S97P029P011nsss(0) <='0';
          end if;
        if(cVar1S8S97N045P043N019P024(0)='1' AND  B(14)='1' AND A(14)='0' AND A(25)='1' )then
          cVar2S8S97P029N011P008nsss(0) <='1';
          else
          cVar2S8S97P029N011P008nsss(0) <='0';
          end if;
        if(cVar1S9S97N045P043N019P024(0)='1' AND  B(14)='0' AND B(10)='1' AND B(16)='0' )then
          cVar2S9S97N029P037P025nsss(0) <='1';
          else
          cVar2S9S97N029P037P025nsss(0) <='0';
          end if;
        if(cVar1S10S97N045P043N019P024(0)='1' AND  B(14)='0' AND B(10)='0' AND E(15)='1' )then
          cVar2S10S97N029N037P040nsss(0) <='1';
          else
          cVar2S10S97N029N037P040nsss(0) <='0';
          end if;
        if(cVar1S11S97N045P043N019P024(0)='1' AND  A(22)='0' AND B(11)='0' AND A(26)='1' )then
          cVar2S11S97P014P035P006nsss(0) <='1';
          else
          cVar2S11S97P014P035P006nsss(0) <='0';
          end if;
        if(cVar1S14S97N045P043N022N057(0)='1' AND  B(21)='0' AND A(25)='1' AND A(12)='1' )then
          cVar2S14S97P034P008P015nsss(0) <='1';
          else
          cVar2S14S97P034P008P015nsss(0) <='0';
          end if;
        if(cVar1S0S98P019P045P026P062(0)='1' AND  A(17)='1' )then
          cVar2S0S98P005nsss(0) <='1';
          else
          cVar2S0S98P005nsss(0) <='0';
          end if;
        if(cVar1S1S98P019P045P026P062(0)='1' AND  A(17)='0' AND E(16)='0' )then
          cVar2S1S98N005P069nsss(0) <='1';
          else
          cVar2S1S98N005P069nsss(0) <='0';
          end if;
        if(cVar1S2S98P019N045P024P029(0)='1' AND  E(16)='1' )then
          cVar2S2S98P069nsss(0) <='1';
          else
          cVar2S2S98P069nsss(0) <='0';
          end if;
        if(cVar1S3S98P019N045P024P029(0)='1' AND  E(16)='0' AND D(11)='1' )then
          cVar2S3S98N069P054nsss(0) <='1';
          else
          cVar2S3S98N069P054nsss(0) <='0';
          end if;
        if(cVar1S4S98P019N045P024N029(0)='1' AND  E(21)='0' AND D(22)='0' AND B(16)='0' )then
          cVar2S4S98P049P043P025nsss(0) <='1';
          else
          cVar2S4S98P049P043P025nsss(0) <='0';
          end if;
        if(cVar1S5S98P019N045P024N029(0)='1' AND  E(21)='1' AND B(25)='1' )then
          cVar2S5S98P049P026nsss(0) <='1';
          else
          cVar2S5S98P049P026nsss(0) <='0';
          end if;
        if(cVar1S6S98P019N045P024N029(0)='1' AND  E(21)='1' AND B(25)='0' AND B(15)='1' )then
          cVar2S6S98P049N026P027nsss(0) <='1';
          else
          cVar2S6S98P049N026P027nsss(0) <='0';
          end if;
        if(cVar1S7S98P019N045P024P001(0)='1' AND  B(15)='0' AND E(21)='1' AND D(21)='1' )then
          cVar2S7S98P027P049P047nsss(0) <='1';
          else
          cVar2S7S98P027P049P047nsss(0) <='0';
          end if;
        if(cVar1S8S98P019P051P025P016(0)='1' AND  A(23)='1' )then
          cVar2S8S98P012nsss(0) <='1';
          else
          cVar2S8S98P012nsss(0) <='0';
          end if;
        if(cVar1S9S98P019P051P025P016(0)='1' AND  A(23)='0' AND A(12)='0' )then
          cVar2S9S98N012P015nsss(0) <='1';
          else
          cVar2S9S98N012P015nsss(0) <='0';
          end if;
        if(cVar1S10S98P019P051P025P016(0)='1' AND  A(12)='1' )then
          cVar2S10S98P015nsss(0) <='1';
          else
          cVar2S10S98P015nsss(0) <='0';
          end if;
        if(cVar1S11S98P019P051N025P029(0)='1' AND  A(29)='1' AND A(23)='0' AND B(12)='0' )then
          cVar2S11S98P000P012P033nsss(0) <='1';
          else
          cVar2S11S98P000P012P033nsss(0) <='0';
          end if;
        if(cVar1S12S98P019P051N025P029(0)='1' AND  A(29)='1' AND A(23)='1' AND A(24)='1' )then
          cVar2S12S98P000P012P010nsss(0) <='1';
          else
          cVar2S12S98P000P012P010nsss(0) <='0';
          end if;
        if(cVar1S13S98P019P051N025P029(0)='1' AND  A(29)='0' AND B(23)='1' AND B(13)='0' )then
          cVar2S13S98N000P030P031nsss(0) <='1';
          else
          cVar2S13S98N000P030P031nsss(0) <='0';
          end if;
        if(cVar1S14S98P019P051N025P029(0)='1' AND  A(29)='0' AND B(23)='0' AND B(13)='1' )then
          cVar2S14S98N000N030P031nsss(0) <='1';
          else
          cVar2S14S98N000N030P031nsss(0) <='0';
          end if;
        if(cVar1S15S98P019P051N025P029(0)='1' AND  E(12)='1' )then
          cVar2S15S98P052nsss(0) <='1';
          else
          cVar2S15S98P052nsss(0) <='0';
          end if;
        if(cVar1S16S98P019P051P037P024(0)='1' AND  D(16)='0' AND A(22)='0' )then
          cVar2S16S98P067P014nsss(0) <='1';
          else
          cVar2S16S98P067P014nsss(0) <='0';
          end if;
        if(cVar1S17S98P019P051N037P008(0)='1' AND  A(23)='0' )then
          cVar2S17S98P012nsss(0) <='1';
          else
          cVar2S17S98P012nsss(0) <='0';
          end if;
        if(cVar1S18S98P019P051N037N008(0)='1' AND  A(11)='0' AND A(22)='1' AND A(20)='0' )then
          cVar2S18S98P017P014P018nsss(0) <='1';
          else
          cVar2S18S98P017P014P018nsss(0) <='0';
          end if;
        if(cVar1S2S99P045P030N025N022(0)='1' AND  B(17)='1' )then
          cVar2S2S99P023nsss(0) <='1';
          else
          cVar2S2S99P023nsss(0) <='0';
          end if;
        if(cVar1S3S99P045P030N025N022(0)='1' AND  B(17)='0' AND B(26)='1' )then
          cVar2S3S99N023P024nsss(0) <='1';
          else
          cVar2S3S99N023P024nsss(0) <='0';
          end if;
        if(cVar1S4S99N045P019P043P051(0)='1' AND  B(14)='0' AND D(16)='1' AND B(26)='0' )then
          cVar2S4S99P029P067P024nsss(0) <='1';
          else
          cVar2S4S99P029P067P024nsss(0) <='0';
          end if;
        if(cVar1S5S99N045P019P043P051(0)='1' AND  B(14)='0' AND D(16)='0' AND E(12)='0' )then
          cVar2S5S99P029N067P052nsss(0) <='1';
          else
          cVar2S5S99P029N067P052nsss(0) <='0';
          end if;
        if(cVar1S6S99N045P019P043P051(0)='1' AND  B(14)='1' AND E(12)='1' )then
          cVar2S6S99P029P052nsss(0) <='1';
          else
          cVar2S6S99P029P052nsss(0) <='0';
          end if;
        if(cVar1S7S99N045P019P043P051(0)='1' AND  B(26)='0' AND B(10)='1' AND D(16)='0' )then
          cVar2S7S99P024P037P067nsss(0) <='1';
          else
          cVar2S7S99P024P037P067nsss(0) <='0';
          end if;
        if(cVar1S8S99N045P019P043P051(0)='1' AND  B(26)='0' AND B(10)='0' AND A(25)='1' )then
          cVar2S8S99P024N037P008nsss(0) <='1';
          else
          cVar2S8S99P024N037P008nsss(0) <='0';
          end if;
        if(cVar1S9S99N045P019P043P014(0)='1' AND  A(11)='1' )then
          cVar2S9S99P017nsss(0) <='1';
          else
          cVar2S9S99P017nsss(0) <='0';
          end if;
        if(cVar1S10S99N045P019P043P014(0)='1' AND  A(11)='0' AND A(20)='0' )then
          cVar2S10S99N017P018nsss(0) <='1';
          else
          cVar2S10S99N017P018nsss(0) <='0';
          end if;
        if(cVar1S11S99N045N019P029P011(0)='1' AND  D(11)='1' )then
          cVar2S11S99P054nsss(0) <='1';
          else
          cVar2S11S99P054nsss(0) <='0';
          end if;
        if(cVar1S12S99N045N019P029P011(0)='1' AND  D(11)='0' AND D(20)='1' )then
          cVar2S12S99N054P051nsss(0) <='1';
          else
          cVar2S12S99N054P051nsss(0) <='0';
          end if;
        if(cVar1S13S99N045N019P029P011(0)='1' AND  D(11)='0' AND D(20)='0' AND E(12)='1' )then
          cVar2S13S99N054N051P052nsss(0) <='1';
          else
          cVar2S13S99N054N051P052nsss(0) <='0';
          end if;
        if(cVar1S14S99N045N019P029N011(0)='1' AND  D(19)='0' AND A(25)='1' )then
          cVar2S14S99P055P008nsss(0) <='1';
          else
          cVar2S14S99P055P008nsss(0) <='0';
          end if;
        if(cVar1S15S99N045N019P029N011(0)='1' AND  D(19)='0' AND A(25)='0' AND A(24)='1' )then
          cVar2S15S99P055N008P010nsss(0) <='1';
          else
          cVar2S15S99P055N008P010nsss(0) <='0';
          end if;
        if(cVar1S16S99N045N019N029P032(0)='1' AND  B(20)='0' AND A(13)='1' AND D(17)='0' )then
          cVar2S16S99P036P013P063nsss(0) <='1';
          else
          cVar2S16S99P036P013P063nsss(0) <='0';
          end if;
        if(cVar1S17S99N045N019N029P032(0)='1' AND  B(20)='0' AND A(13)='0' AND A(24)='0' )then
          cVar2S17S99P036N013P010nsss(0) <='1';
          else
          cVar2S17S99P036N013P010nsss(0) <='0';
          end if;
        if(cVar1S18S99N045N019N029N032(0)='1' AND  E(13)='1' AND A(11)='0' AND A(18)='0' )then
          cVar2S18S99P048P017P003nsss(0) <='1';
          else
          cVar2S18S99P048P017P003nsss(0) <='0';
          end if;
        if(cVar1S19S99N045N019N029N032(0)='1' AND  E(13)='0' AND B(13)='1' AND A(13)='1' )then
          cVar2S19S99N048P031P013nsss(0) <='1';
          else
          cVar2S19S99N048P031P013nsss(0) <='0';
          end if;
        if(cVar1S0S100P019P045P026P062(0)='1' AND  A(17)='1' )then
          cVar2S0S100P005nsss(0) <='1';
          else
          cVar2S0S100P005nsss(0) <='0';
          end if;
        if(cVar1S1S100P019P045P026P062(0)='1' AND  A(17)='0' AND E(16)='0' )then
          cVar2S1S100N005P069nsss(0) <='1';
          else
          cVar2S1S100N005P069nsss(0) <='0';
          end if;
        if(cVar1S2S100P019N045P029P011(0)='1' AND  D(11)='1' )then
          cVar2S2S100P054nsss(0) <='1';
          else
          cVar2S2S100P054nsss(0) <='0';
          end if;
        if(cVar1S3S100P019N045P029P011(0)='1' AND  D(11)='0' AND D(20)='1' )then
          cVar2S3S100N054P051nsss(0) <='1';
          else
          cVar2S3S100N054P051nsss(0) <='0';
          end if;
        if(cVar1S4S100P019N045P029P011(0)='1' AND  D(11)='0' AND D(20)='0' AND E(12)='1' )then
          cVar2S4S100N054N051P052nsss(0) <='1';
          else
          cVar2S4S100N054N051P052nsss(0) <='0';
          end if;
        if(cVar1S5S100P019N045P029N011(0)='1' AND  D(19)='0' AND B(21)='1' )then
          cVar2S5S100P055P034nsss(0) <='1';
          else
          cVar2S5S100P055P034nsss(0) <='0';
          end if;
        if(cVar1S6S100P019N045P029N011(0)='1' AND  D(19)='0' AND B(21)='0' AND A(12)='1' )then
          cVar2S6S100P055N034P015nsss(0) <='1';
          else
          cVar2S6S100P055N034P015nsss(0) <='0';
          end if;
        if(cVar1S7S100P019N045N029P008(0)='1' AND  E(20)='0' AND A(23)='1' )then
          cVar2S7S100P053P012nsss(0) <='1';
          else
          cVar2S7S100P053P012nsss(0) <='0';
          end if;
        if(cVar1S8S100P019N045N029P008(0)='1' AND  E(20)='0' AND A(23)='0' AND A(29)='0' )then
          cVar2S8S100P053N012P000nsss(0) <='1';
          else
          cVar2S8S100P053N012P000nsss(0) <='0';
          end if;
        if(cVar1S9S100P019N045N029P008(0)='1' AND  E(20)='1' AND E(11)='0' AND A(15)='1' )then
          cVar2S9S100P053P056P009nsss(0) <='1';
          else
          cVar2S9S100P053P056P009nsss(0) <='0';
          end if;
        if(cVar1S10S100P019N045N029P008(0)='1' AND  E(20)='1' AND A(13)='0' )then
          cVar2S10S100P053P013nsss(0) <='1';
          else
          cVar2S10S100P053P013nsss(0) <='0';
          end if;
        if(cVar1S11S100P019N045N029P008(0)='1' AND  E(20)='0' AND A(26)='1' AND A(22)='0' )then
          cVar2S11S100N053P006P014nsss(0) <='1';
          else
          cVar2S11S100N053P006P014nsss(0) <='0';
          end if;
        if(cVar1S13S100P019P013P045N043(0)='1' AND  A(23)='1' )then
          cVar2S13S100P012nsss(0) <='1';
          else
          cVar2S13S100P012nsss(0) <='0';
          end if;
        if(cVar1S14S100P019P013P045N043(0)='1' AND  A(23)='0' AND D( 8)='0' AND A(20)='1' )then
          cVar2S14S100N012P066P018nsss(0) <='1';
          else
          cVar2S14S100N012P066P018nsss(0) <='0';
          end if;
        if(cVar1S15S100P019P013N045P067(0)='1' AND  A(20)='0' AND E(12)='1' )then
          cVar2S15S100P018P052nsss(0) <='1';
          else
          cVar2S15S100P018P052nsss(0) <='0';
          end if;
        if(cVar1S16S100P019P013N045P067(0)='1' AND  A(20)='0' AND E(12)='0' AND A(24)='0' )then
          cVar2S16S100P018N052P010nsss(0) <='1';
          else
          cVar2S16S100P018N052P010nsss(0) <='0';
          end if;
        if(cVar1S17S100P019P013N045N067(0)='1' AND  E(13)='0' AND D(10)='1' AND A(12)='0' )then
          cVar2S17S100P048P058P015nsss(0) <='1';
          else
          cVar2S17S100P048P058P015nsss(0) <='0';
          end if;
        if(cVar1S18S100P019P013N045N067(0)='1' AND  E(13)='1' AND A(21)='0' AND D(13)='1' )then
          cVar2S18S100P048P016P046nsss(0) <='1';
          else
          cVar2S18S100P048P016P046nsss(0) <='0';
          end if;
        if(cVar1S19S100P019P013P039P041(0)='1' AND  B(28)='0' AND B(14)='1' AND A(12)='0' )then
          cVar2S19S100P020P029P015nsss(0) <='1';
          else
          cVar2S19S100P020P029P015nsss(0) <='0';
          end if;
        if(cVar1S1S101P045P030P035N025(0)='1' AND  B(27)='1' )then
          cVar2S1S101P022nsss(0) <='1';
          else
          cVar2S1S101P022nsss(0) <='0';
          end if;
        if(cVar1S2S101P045P030P035N025(0)='1' AND  B(27)='0' AND B(17)='1' )then
          cVar2S2S101N022P023nsss(0) <='1';
          else
          cVar2S2S101N022P023nsss(0) <='0';
          end if;
        if(cVar1S3S101P045P030P035N025(0)='1' AND  B(27)='0' AND B(17)='0' AND B(26)='1' )then
          cVar2S3S101N022N023P024nsss(0) <='1';
          else
          cVar2S3S101N022N023P024nsss(0) <='0';
          end if;
        if(cVar1S4S101N045P019P043P023(0)='1' AND  A(26)='0' AND E(14)='0' AND A(28)='0' )then
          cVar2S4S101P006P044P002nsss(0) <='1';
          else
          cVar2S4S101P006P044P002nsss(0) <='0';
          end if;
        if(cVar1S5S101N045P019P043P023(0)='1' AND  A(26)='0' AND E(14)='1' AND A(21)='0' )then
          cVar2S5S101P006P044P016nsss(0) <='1';
          else
          cVar2S5S101P006P044P016nsss(0) <='0';
          end if;
        if(cVar1S6S101N045P019P043P023(0)='1' AND  A(26)='1' AND B(20)='0' AND B(23)='0' )then
          cVar2S6S101P006P036P030nsss(0) <='1';
          else
          cVar2S6S101P006P036P030nsss(0) <='0';
          end if;
        if(cVar1S7S101N045P019P043P023(0)='1' AND  A(23)='0' AND A(11)='0' )then
          cVar2S7S101P012P017nsss(0) <='1';
          else
          cVar2S7S101P012P017nsss(0) <='0';
          end if;
        if(cVar1S8S101N045P019P043P014(0)='1' AND  A(11)='1' )then
          cVar2S8S101P017nsss(0) <='1';
          else
          cVar2S8S101P017nsss(0) <='0';
          end if;
        if(cVar1S9S101N045P019P043P014(0)='1' AND  A(11)='0' AND A(20)='0' )then
          cVar2S9S101N017P018nsss(0) <='1';
          else
          cVar2S9S101N017P018nsss(0) <='0';
          end if;
        if(cVar1S10S101N045N019P029P024(0)='1' AND  E(16)='1' )then
          cVar2S10S101P069nsss(0) <='1';
          else
          cVar2S10S101P069nsss(0) <='0';
          end if;
        if(cVar1S11S101N045N019P029P024(0)='1' AND  E(16)='0' AND B(24)='0' AND A(20)='0' )then
          cVar2S11S101N069P028P018nsss(0) <='1';
          else
          cVar2S11S101N069P028P018nsss(0) <='0';
          end if;
        if(cVar1S12S101N045N019N029P040(0)='1' AND  A(28)='1' )then
          cVar2S12S101P002nsss(0) <='1';
          else
          cVar2S12S101P002nsss(0) <='0';
          end if;
        if(cVar1S13S101N045N019N029P040(0)='1' AND  A(28)='0' AND B(18)='1' )then
          cVar2S13S101N002P021nsss(0) <='1';
          else
          cVar2S13S101N002P021nsss(0) <='0';
          end if;
        if(cVar1S1S102P019P045P026N005(0)='1' AND  D( 9)='0' )then
          cVar2S1S102P062nsss(0) <='1';
          else
          cVar2S1S102P062nsss(0) <='0';
          end if;
        if(cVar1S2S102P019N045P029P061(0)='1' AND  E(16)='1' )then
          cVar2S2S102P069nsss(0) <='1';
          else
          cVar2S2S102P069nsss(0) <='0';
          end if;
        if(cVar1S3S102P019N045P029P061(0)='1' AND  E(16)='0' AND B(24)='0' AND B(25)='0' )then
          cVar2S3S102N069P028P026nsss(0) <='1';
          else
          cVar2S3S102N069P028P026nsss(0) <='0';
          end if;
        if(cVar1S4S102P019N045N029P054(0)='1' AND  E(11)='0' AND E(20)='1' )then
          cVar2S4S102P056P053nsss(0) <='1';
          else
          cVar2S4S102P056P053nsss(0) <='0';
          end if;
        if(cVar1S5S102P019N045N029P054(0)='1' AND  E(11)='0' AND E(20)='0' AND D(20)='0' )then
          cVar2S5S102P056N053P051nsss(0) <='1';
          else
          cVar2S5S102P056N053P051nsss(0) <='0';
          end if;
        if(cVar1S6S102P019N045N029P054(0)='1' AND  E(11)='1' AND D(10)='1' AND A(23)='1' )then
          cVar2S6S102P056P058P012nsss(0) <='1';
          else
          cVar2S6S102P056P058P012nsss(0) <='0';
          end if;
        if(cVar1S7S102P019N045N029P054(0)='1' AND  E(11)='1' AND D(10)='0' AND D( 9)='1' )then
          cVar2S7S102P056N058P062nsss(0) <='1';
          else
          cVar2S7S102P056N058P062nsss(0) <='0';
          end if;
        if(cVar1S8S102P019N045N029P054(0)='1' AND  B(13)='1' AND E( 8)='1' )then
          cVar2S8S102P031P068nsss(0) <='1';
          else
          cVar2S8S102P031P068nsss(0) <='0';
          end if;
        if(cVar1S9S102P019N045N029P054(0)='1' AND  B(13)='1' AND E( 8)='0' AND D(17)='1' )then
          cVar2S9S102P031N068P063nsss(0) <='1';
          else
          cVar2S9S102P031N068P063nsss(0) <='0';
          end if;
        if(cVar1S10S102P019N045N029P054(0)='1' AND  B(13)='0' AND A(27)='0' AND B(21)='1' )then
          cVar2S10S102N031P004P034nsss(0) <='1';
          else
          cVar2S10S102N031P004P034nsss(0) <='0';
          end if;
        if(cVar1S11S102P019P051P018P057(0)='1' AND  B(23)='0' AND B(12)='0' AND D(12)='0' )then
          cVar2S11S102P030P033P050nsss(0) <='1';
          else
          cVar2S11S102P030P033P050nsss(0) <='0';
          end if;
        if(cVar1S12S102P019P051P018P057(0)='1' AND  B(23)='0' AND B(12)='1' AND E(18)='1' )then
          cVar2S12S102P030P033P061nsss(0) <='1';
          else
          cVar2S12S102P030P033P061nsss(0) <='0';
          end if;
        if(cVar1S13S102P019P051P018P057(0)='1' AND  B(23)='1' AND A(21)='0' AND A(11)='1' )then
          cVar2S13S102P030P016P017nsss(0) <='1';
          else
          cVar2S13S102P030P016P017nsss(0) <='0';
          end if;
        if(cVar1S14S102P019P051P018P057(0)='1' AND  A(25)='0' AND D(19)='1' AND E( 8)='0' )then
          cVar2S14S102P008P055P068nsss(0) <='1';
          else
          cVar2S14S102P008P055P068nsss(0) <='0';
          end if;
        if(cVar1S15S102P019P051N018P053(0)='1' AND  D(12)='1' AND E(17)='0' AND A(13)='0' )then
          cVar2S15S102P050P065P013nsss(0) <='1';
          else
          cVar2S15S102P050P065P013nsss(0) <='0';
          end if;
        if(cVar1S16S102P019P051N018P053(0)='1' AND  D(12)='0' AND B(26)='1' AND A(21)='0' )then
          cVar2S16S102N050P024P016nsss(0) <='1';
          else
          cVar2S16S102N050P024P016nsss(0) <='0';
          end if;
        if(cVar1S17S102P019P051N018P053(0)='1' AND  D(12)='0' AND B(26)='0' AND D(19)='1' )then
          cVar2S17S102N050N024P055nsss(0) <='1';
          else
          cVar2S17S102N050N024P055nsss(0) <='0';
          end if;
        if(cVar1S18S102P019P051N018P053(0)='1' AND  A(11)='0' AND A(12)='1' )then
          cVar2S18S102P017P015nsss(0) <='1';
          else
          cVar2S18S102P017P015nsss(0) <='0';
          end if;
        if(cVar1S19S102P019P051P024P037(0)='1' AND  B(21)='0' AND B(20)='0' AND A(22)='0' )then
          cVar2S19S102P034P036P014nsss(0) <='1';
          else
          cVar2S19S102P034P036P014nsss(0) <='0';
          end if;
        if(cVar1S20S102P019P051P024N037(0)='1' AND  E( 9)='0' AND B(25)='1' )then
          cVar2S20S102P064P026nsss(0) <='1';
          else
          cVar2S20S102P064P026nsss(0) <='0';
          end if;
        if(cVar1S2S103P045P030N025N022(0)='1' AND  B(17)='1' )then
          cVar2S2S103P023nsss(0) <='1';
          else
          cVar2S2S103P023nsss(0) <='0';
          end if;
        if(cVar1S3S103P045P030N025N022(0)='1' AND  B(17)='0' AND B(26)='1' )then
          cVar2S3S103N023P024nsss(0) <='1';
          else
          cVar2S3S103N023P024nsss(0) <='0';
          end if;
        if(cVar1S6S103N045P052N065N062(0)='1' AND  A(25)='1' AND A(22)='0' )then
          cVar2S6S103P008P014nsss(0) <='1';
          else
          cVar2S6S103P008P014nsss(0) <='0';
          end if;
        if(cVar1S7S103N045P052N065N062(0)='1' AND  A(25)='0' AND A(24)='1' )then
          cVar2S7S103N008P010nsss(0) <='1';
          else
          cVar2S7S103N008P010nsss(0) <='0';
          end if;
        if(cVar1S8S103N045N052P043P018(0)='1' AND  A(17)='0' AND E(18)='0' AND A(10)='1' )then
          cVar2S8S103P005P061P019nsss(0) <='1';
          else
          cVar2S8S103P005P061P019nsss(0) <='0';
          end if;
        if(cVar1S9S103N045N052P043P018(0)='1' AND  A(17)='1' AND A(25)='0' AND D(14)='1' )then
          cVar2S9S103P005P008P042nsss(0) <='1';
          else
          cVar2S9S103P005P008P042nsss(0) <='0';
          end if;
        if(cVar1S10S103N045N052P043P018(0)='1' AND  D(23)='0' AND B(16)='0' AND D(16)='1' )then
          cVar2S10S103P039P025P067nsss(0) <='1';
          else
          cVar2S10S103P039P025P067nsss(0) <='0';
          end if;
        if(cVar1S11S103N045N052P043P018(0)='1' AND  D(23)='0' AND B(16)='1' AND A(16)='1' )then
          cVar2S11S103P039P025P007nsss(0) <='1';
          else
          cVar2S11S103P039P025P007nsss(0) <='0';
          end if;
        if(cVar1S12S103N045N052P043P018(0)='1' AND  D(23)='1' AND A(21)='0' AND A(11)='0' )then
          cVar2S12S103P039P016P017nsss(0) <='1';
          else
          cVar2S12S103P039P016P017nsss(0) <='0';
          end if;
        if(cVar1S13S103N045N052P043P063(0)='1' AND  A(18)='1' )then
          cVar2S13S103P003nsss(0) <='1';
          else
          cVar2S13S103P003nsss(0) <='0';
          end if;
        if(cVar1S14S103N045N052P043P063(0)='1' AND  A(18)='0' AND A(13)='0' AND B(26)='1' )then
          cVar2S14S103N003P013P024nsss(0) <='1';
          else
          cVar2S14S103N003P013P024nsss(0) <='0';
          end if;
        if(cVar1S1S104P019P045P026N005(0)='1' AND  D( 9)='0' AND E(16)='0' )then
          cVar2S1S104P062P069nsss(0) <='1';
          else
          cVar2S1S104P062P069nsss(0) <='0';
          end if;
        if(cVar1S2S104P019N045P029P011(0)='1' AND  A(13)='0' )then
          cVar2S2S104P013nsss(0) <='1';
          else
          cVar2S2S104P013nsss(0) <='0';
          end if;
        if(cVar1S3S104P019N045P029N011(0)='1' AND  D(19)='0' AND A(15)='1' )then
          cVar2S3S104P055P009nsss(0) <='1';
          else
          cVar2S3S104P055P009nsss(0) <='0';
          end if;
        if(cVar1S4S104P019N045P029N011(0)='1' AND  D(19)='0' AND A(15)='0' AND A(25)='1' )then
          cVar2S4S104P055N009P008nsss(0) <='1';
          else
          cVar2S4S104P055N009P008nsss(0) <='0';
          end if;
        if(cVar1S5S104P019N045N029P069(0)='1' AND  D(20)='1' AND A(14)='1' AND A(23)='0' )then
          cVar2S5S104P051P011P012nsss(0) <='1';
          else
          cVar2S5S104P051P011P012nsss(0) <='0';
          end if;
        if(cVar1S6S104P019N045N029P069(0)='1' AND  D(20)='1' AND A(14)='0' AND A(24)='1' )then
          cVar2S6S104P051N011P010nsss(0) <='1';
          else
          cVar2S6S104P051N011P010nsss(0) <='0';
          end if;
        if(cVar1S7S104P019N045N029P069(0)='1' AND  D(20)='0' AND E(20)='0' )then
          cVar2S7S104N051P053nsss(0) <='1';
          else
          cVar2S7S104N051P053nsss(0) <='0';
          end if;
        if(cVar1S8S104P019N045N029P069(0)='1' AND  A(15)='0' AND E(14)='1' )then
          cVar2S8S104P009P044nsss(0) <='1';
          else
          cVar2S8S104P009P044nsss(0) <='0';
          end if;
        if(cVar1S9S104P019N045N029P069(0)='1' AND  A(15)='1' AND B(20)='0' AND A(14)='0' )then
          cVar2S9S104P009P036P011nsss(0) <='1';
          else
          cVar2S9S104P009P036P011nsss(0) <='0';
          end if;
        if(cVar1S11S104P019P067P047N006(0)='1' AND  E(21)='0' )then
          cVar2S11S104P049nsss(0) <='1';
          else
          cVar2S11S104P049nsss(0) <='0';
          end if;
        if(cVar1S12S104P019P067P047N006(0)='1' AND  E(21)='1' AND A(20)='0' )then
          cVar2S12S104P049P018nsss(0) <='1';
          else
          cVar2S12S104P049P018nsss(0) <='0';
          end if;
        if(cVar1S13S104P019P067N047P069(0)='1' AND  A(20)='1' AND A(17)='1' AND A(23)='0' )then
          cVar2S13S104P018P005P012nsss(0) <='1';
          else
          cVar2S13S104P018P005P012nsss(0) <='0';
          end if;
        if(cVar1S14S104P019P067N047P069(0)='1' AND  A(20)='0' AND D(11)='1' AND A(23)='1' )then
          cVar2S14S104N018P054P012nsss(0) <='1';
          else
          cVar2S14S104N018P054P012nsss(0) <='0';
          end if;
        if(cVar1S15S104P019P067N047P069(0)='1' AND  A(22)='0' AND B(20)='1' )then
          cVar2S15S104P014P036nsss(0) <='1';
          else
          cVar2S15S104P014P036nsss(0) <='0';
          end if;
        if(cVar1S16S104P019P067N047P069(0)='1' AND  A(22)='0' AND B(20)='0' AND A(14)='0' )then
          cVar2S16S104P014N036P011nsss(0) <='1';
          else
          cVar2S16S104P014N036P011nsss(0) <='0';
          end if;
        if(cVar1S18S104P019P067P024N042(0)='1' AND  E(12)='1' )then
          cVar2S18S104P052nsss(0) <='1';
          else
          cVar2S18S104P052nsss(0) <='0';
          end if;
        if(cVar1S19S104P019P067P024P069(0)='1' AND  D(17)='0' AND A(20)='0' )then
          cVar2S19S104P063P018nsss(0) <='1';
          else
          cVar2S19S104P063P018nsss(0) <='0';
          end if;
        if(cVar1S1S105P045P030P035N025(0)='1' AND  B(27)='1' )then
          cVar2S1S105P022nsss(0) <='1';
          else
          cVar2S1S105P022nsss(0) <='0';
          end if;
        if(cVar1S2S105P045P030P035N025(0)='1' AND  B(27)='0' AND E(19)='0' )then
          cVar2S2S105N022P057nsss(0) <='1';
          else
          cVar2S2S105N022P057nsss(0) <='0';
          end if;
        if(cVar1S3S105N045P029P059P028(0)='1' AND  D(20)='1' )then
          cVar2S3S105P051nsss(0) <='1';
          else
          cVar2S3S105P051nsss(0) <='0';
          end if;
        if(cVar1S4S105N045P029P059P028(0)='1' AND  D(20)='0' AND A(29)='0' AND B(12)='0' )then
          cVar2S4S105N051P000P033nsss(0) <='1';
          else
          cVar2S4S105N051P000P033nsss(0) <='0';
          end if;
        if(cVar1S5S105N045N029P043P062(0)='1' AND  E(12)='1' AND A(25)='0' )then
          cVar2S5S105P052P008nsss(0) <='1';
          else
          cVar2S5S105P052P008nsss(0) <='0';
          end if;
        if(cVar1S6S105N045N029P043P062(0)='1' AND  E(12)='0' AND B(11)='1' AND D(20)='0' )then
          cVar2S6S105N052P035P051nsss(0) <='1';
          else
          cVar2S6S105N052P035P051nsss(0) <='0';
          end if;
        if(cVar1S7S105N045N029P043N062(0)='1' AND  E( 9)='0' AND A(29)='1' AND D(20)='0' )then
          cVar2S7S105P064P000P051nsss(0) <='1';
          else
          cVar2S7S105P064P000P051nsss(0) <='0';
          end if;
        if(cVar1S8S105N045N029P043N062(0)='1' AND  E( 9)='0' AND A(29)='0' AND B(28)='1' )then
          cVar2S8S105P064N000P020nsss(0) <='1';
          else
          cVar2S8S105P064N000P020nsss(0) <='0';
          end if;
        if(cVar1S9S105N045N029P043N062(0)='1' AND  E( 9)='1' AND E(19)='1' )then
          cVar2S9S105P064P057nsss(0) <='1';
          else
          cVar2S9S105P064P057nsss(0) <='0';
          end if;
        if(cVar1S11S105N045N029P043N022(0)='1' AND  D(12)='0' AND A(25)='1' AND A(10)='0' )then
          cVar2S11S105P050P008P019nsss(0) <='1';
          else
          cVar2S11S105P050P008P019nsss(0) <='0';
          end if;
        if(cVar1S0S106P020P039P041P002(0)='1' AND  D(20)='1' AND A(14)='1' AND E(16)='0' )then
          cVar2S0S106P051P011P069nsss(0) <='1';
          else
          cVar2S0S106P051P011P069nsss(0) <='0';
          end if;
        if(cVar1S1S106P020P039P041P002(0)='1' AND  D(20)='1' AND A(14)='0' AND A(25)='1' )then
          cVar2S1S106P051N011P008nsss(0) <='1';
          else
          cVar2S1S106P051N011P008nsss(0) <='0';
          end if;
        if(cVar1S2S106P020P039P041P002(0)='1' AND  D(20)='0' AND E(22)='1' )then
          cVar2S2S106N051P045nsss(0) <='1';
          else
          cVar2S2S106N051P045nsss(0) <='0';
          end if;
        if(cVar1S3S106P020P039P041P002(0)='1' AND  D(20)='0' AND E(22)='0' AND A(16)='0' )then
          cVar2S3S106N051N045P007nsss(0) <='1';
          else
          cVar2S3S106N051N045P007nsss(0) <='0';
          end if;
        if(cVar1S4S106P020P039P041P002(0)='1' AND  D(14)='1' )then
          cVar2S4S106P042nsss(0) <='1';
          else
          cVar2S4S106P042nsss(0) <='0';
          end if;
        if(cVar1S5S106P020P039P041P002(0)='1' AND  D(14)='0' AND A(16)='1' AND A(22)='0' )then
          cVar2S5S106N042P007P014nsss(0) <='1';
          else
          cVar2S5S106N042P007P014nsss(0) <='0';
          end if;
        if(cVar1S6S106P020P039P041P002(0)='1' AND  D(14)='0' AND A(16)='0' AND B(23)='1' )then
          cVar2S6S106N042N007P030nsss(0) <='1';
          else
          cVar2S6S106N042N007P030nsss(0) <='0';
          end if;
        if(cVar1S8S106P020P039P012P060(0)='1' AND  A(18)='1' )then
          cVar2S8S106P003nsss(0) <='1';
          else
          cVar2S8S106P003nsss(0) <='0';
          end if;
        if(cVar1S9S106P020P039P012P060(0)='1' AND  A(18)='0' AND B(12)='1' )then
          cVar2S9S106N003P033nsss(0) <='1';
          else
          cVar2S9S106N003P033nsss(0) <='0';
          end if;
        if(cVar1S10S106P020P039P012P060(0)='1' AND  A(18)='0' AND B(12)='0' AND A(22)='1' )then
          cVar2S10S106N003N033P014nsss(0) <='1';
          else
          cVar2S10S106N003N033P014nsss(0) <='0';
          end if;
        if(cVar1S12S106P020N039P000P017(0)='1' AND  A(14)='0' AND B(20)='1' )then
          cVar2S12S106P011P036nsss(0) <='1';
          else
          cVar2S12S106P011P036nsss(0) <='0';
          end if;
        if(cVar1S13S106P020N039P000P017(0)='1' AND  A(14)='0' AND B(20)='0' AND D( 9)='0' )then
          cVar2S13S106P011N036P062nsss(0) <='1';
          else
          cVar2S13S106P011N036P062nsss(0) <='0';
          end if;
        if(cVar1S14S106P020N039P000N017(0)='1' AND  B(11)='0' AND B(21)='1' )then
          cVar2S14S106P035P034nsss(0) <='1';
          else
          cVar2S14S106P035P034nsss(0) <='0';
          end if;
        if(cVar1S0S107P051P041P024P053(0)='1' AND  A(29)='0' )then
          cVar2S0S107P000nsss(0) <='1';
          else
          cVar2S0S107P000nsss(0) <='0';
          end if;
        if(cVar1S1S107P051P041P024N053(0)='1' AND  E(16)='0' AND A(12)='0' )then
          cVar2S1S107P069P015nsss(0) <='1';
          else
          cVar2S1S107P069P015nsss(0) <='0';
          end if;
        if(cVar1S2S107P051P041P024N053(0)='1' AND  E(16)='0' AND A(12)='1' AND E(21)='1' )then
          cVar2S2S107P069P015P049nsss(0) <='1';
          else
          cVar2S2S107P069P015P049nsss(0) <='0';
          end if;
        if(cVar1S3S107P051P041P024P067(0)='1' AND  A(20)='0' AND E(20)='1' )then
          cVar2S3S107P018P053nsss(0) <='1';
          else
          cVar2S3S107P018P053nsss(0) <='0';
          end if;
        if(cVar1S5S107N051P053P007N025(0)='1' AND  E(17)='0' AND A(15)='1' AND A(14)='0' )then
          cVar2S5S107P065P009P011nsss(0) <='1';
          else
          cVar2S5S107P065P009P011nsss(0) <='0';
          end if;
        if(cVar1S6S107N051P053P007N025(0)='1' AND  E(17)='0' AND A(15)='0' AND D(19)='0' )then
          cVar2S6S107P065N009P055nsss(0) <='1';
          else
          cVar2S6S107P065N009P055nsss(0) <='0';
          end if;
        if(cVar1S7S107N051P053P007N025(0)='1' AND  E(17)='1' AND A(26)='0' AND B(21)='1' )then
          cVar2S7S107P065P006P034nsss(0) <='1';
          else
          cVar2S7S107P065P006P034nsss(0) <='0';
          end if;
        if(cVar1S8S107N051P053N007P048(0)='1' AND  B(16)='0' AND D(18)='1' AND A(27)='0' )then
          cVar2S8S107P025P059P004nsss(0) <='1';
          else
          cVar2S8S107P025P059P004nsss(0) <='0';
          end if;
        if(cVar1S9S107N051P053N007P048(0)='1' AND  B(16)='1' AND A(24)='0' AND B(26)='1' )then
          cVar2S9S107P025P010P024nsss(0) <='1';
          else
          cVar2S9S107P025P010P024nsss(0) <='0';
          end if;
        if(cVar1S10S107N051P053N007P048(0)='1' AND  B(10)='0' AND D( 9)='1' )then
          cVar2S10S107P037P062nsss(0) <='1';
          else
          cVar2S10S107P037P062nsss(0) <='0';
          end if;
        if(cVar1S11S107N051P053P027P030(0)='1' AND  A(21)='1' AND A(13)='0' AND B(20)='0' )then
          cVar2S11S107P016P013P036nsss(0) <='1';
          else
          cVar2S11S107P016P013P036nsss(0) <='0';
          end if;
        if(cVar1S0S108P061P059P051P039(0)='1' AND  B(26)='0' )then
          cVar2S0S108P024nsss(0) <='1';
          else
          cVar2S0S108P024nsss(0) <='0';
          end if;
        if(cVar1S1S108P061P059P051P039(0)='1' AND  B(26)='1' AND A(23)='0' AND A(21)='0' )then
          cVar2S1S108P024P012P016nsss(0) <='1';
          else
          cVar2S1S108P024P012P016nsss(0) <='0';
          end if;
        if(cVar1S2S108P061P059N051P045(0)='1' AND  B(27)='1' )then
          cVar2S2S108P022nsss(0) <='1';
          else
          cVar2S2S108P022nsss(0) <='0';
          end if;
        if(cVar1S3S108P061P059N051P045(0)='1' AND  B(27)='0' AND B(16)='1' )then
          cVar2S3S108N022P025nsss(0) <='1';
          else
          cVar2S3S108N022P025nsss(0) <='0';
          end if;
        if(cVar1S4S108P061P059N051P045(0)='1' AND  B(27)='0' AND B(16)='0' AND B(23)='0' )then
          cVar2S4S108N022N025P030nsss(0) <='1';
          else
          cVar2S4S108N022N025P030nsss(0) <='0';
          end if;
        if(cVar1S5S108P061P059N051N045(0)='1' AND  E(23)='1' AND B(28)='1' )then
          cVar2S5S108P041P020nsss(0) <='1';
          else
          cVar2S5S108P041P020nsss(0) <='0';
          end if;
        if(cVar1S6S108P061P059N051N045(0)='1' AND  E(23)='1' AND B(28)='0' AND A(21)='0' )then
          cVar2S6S108P041N020P016nsss(0) <='1';
          else
          cVar2S6S108P041N020P016nsss(0) <='0';
          end if;
        if(cVar1S7S108P061P059N051N045(0)='1' AND  E(23)='0' AND D(22)='0' )then
          cVar2S7S108N041P043nsss(0) <='1';
          else
          cVar2S7S108N041P043nsss(0) <='0';
          end if;
        if(cVar1S8S108P061P059N051N045(0)='1' AND  E(23)='0' AND D(22)='1' AND A(18)='1' )then
          cVar2S8S108N041P043P003nsss(0) <='1';
          else
          cVar2S8S108N041P043P003nsss(0) <='0';
          end if;
        if(cVar1S9S108P061P059P052P062(0)='1' AND  E(19)='1' AND A(23)='1' )then
          cVar2S9S108P057P012nsss(0) <='1';
          else
          cVar2S9S108P057P012nsss(0) <='0';
          end if;
        if(cVar1S10S108P061P059P052P062(0)='1' AND  E(19)='1' AND A(23)='0' AND A(22)='1' )then
          cVar2S10S108P057N012P014nsss(0) <='1';
          else
          cVar2S10S108P057N012P014nsss(0) <='0';
          end if;
        if(cVar1S11S108P061P059P052P062(0)='1' AND  E(19)='0' AND A(26)='1' )then
          cVar2S11S108N057P006nsss(0) <='1';
          else
          cVar2S11S108N057P006nsss(0) <='0';
          end if;
        if(cVar1S12S108P061P040P033P015(0)='1' AND  B(22)='0' )then
          cVar2S12S108P032nsss(0) <='1';
          else
          cVar2S12S108P032nsss(0) <='0';
          end if;
        if(cVar1S13S108P061P040P033N015(0)='1' AND  D(10)='0' )then
          cVar2S13S108P058nsss(0) <='1';
          else
          cVar2S13S108P058nsss(0) <='0';
          end if;
        if(cVar1S14S108P061P040N033P041(0)='1' AND  D(18)='1' AND B(13)='1' )then
          cVar2S14S108P059P031nsss(0) <='1';
          else
          cVar2S14S108P059P031nsss(0) <='0';
          end if;
        if(cVar1S15S108P061P040N033P041(0)='1' AND  D(18)='0' AND B(22)='1' )then
          cVar2S15S108N059P032nsss(0) <='1';
          else
          cVar2S15S108N059P032nsss(0) <='0';
          end if;
        if(cVar1S16S108P061P040N033P041(0)='1' AND  D(18)='0' AND B(22)='0' AND D(19)='1' )then
          cVar2S16S108N059N032P055nsss(0) <='1';
          else
          cVar2S16S108N059N032P055nsss(0) <='0';
          end if;
        if(cVar1S2S109P022N043N002P003(0)='1' AND  B(12)='1' )then
          cVar2S2S109P033nsss(0) <='1';
          else
          cVar2S2S109P033nsss(0) <='0';
          end if;
        if(cVar1S3S109N022P043P000P056(0)='1' AND  B(23)='1' )then
          cVar2S3S109P030nsss(0) <='1';
          else
          cVar2S3S109P030nsss(0) <='0';
          end if;
        if(cVar1S4S109N022P043P000P056(0)='1' AND  B(23)='0' AND A(13)='1' AND B(13)='1' )then
          cVar2S4S109N030P013P031nsss(0) <='1';
          else
          cVar2S4S109N030P013P031nsss(0) <='0';
          end if;
        if(cVar1S5S109N022P043P000N056(0)='1' AND  D(11)='0' AND E(20)='1' AND B(24)='1' )then
          cVar2S5S109P054P053P028nsss(0) <='1';
          else
          cVar2S5S109P054P053P028nsss(0) <='0';
          end if;
        if(cVar1S6S109N022P043P000N056(0)='1' AND  D(11)='1' AND E(14)='1' )then
          cVar2S6S109P054P044nsss(0) <='1';
          else
          cVar2S6S109P054P044nsss(0) <='0';
          end if;
        if(cVar1S8S109N022P043N025P050(0)='1' AND  B(17)='1' )then
          cVar2S8S109P023nsss(0) <='1';
          else
          cVar2S8S109P023nsss(0) <='0';
          end if;
        if(cVar1S9S109N022P043N025P050(0)='1' AND  B(17)='0' AND B(21)='0' AND A(26)='1' )then
          cVar2S9S109N023P034P006nsss(0) <='1';
          else
          cVar2S9S109N023P034P006nsss(0) <='0';
          end if;
        if(cVar1S0S110P000P051P041P053(0)='1' AND  A(15)='1' AND E(16)='0' )then
          cVar2S0S110P009P069nsss(0) <='1';
          else
          cVar2S0S110P009P069nsss(0) <='0';
          end if;
        if(cVar1S1S110P000P051P041P053(0)='1' AND  A(15)='0' AND A(14)='1' AND A(23)='0' )then
          cVar2S1S110N009P011P012nsss(0) <='1';
          else
          cVar2S1S110N009P011P012nsss(0) <='0';
          end if;
        if(cVar1S2S110P000P051P041P053(0)='1' AND  A(15)='0' AND A(14)='0' AND A(25)='1' )then
          cVar2S2S110N009N011P008nsss(0) <='1';
          else
          cVar2S2S110N009N011P008nsss(0) <='0';
          end if;
        if(cVar1S3S110P000P051P041N053(0)='1' AND  E(16)='0' AND A(12)='0' )then
          cVar2S3S110P069P015nsss(0) <='1';
          else
          cVar2S3S110P069P015nsss(0) <='0';
          end if;
        if(cVar1S4S110P000P051P041N053(0)='1' AND  E(16)='0' AND A(12)='1' AND A(25)='1' )then
          cVar2S4S110P069P015P008nsss(0) <='1';
          else
          cVar2S4S110P069P015P008nsss(0) <='0';
          end if;
        if(cVar1S5S110P000N051P053P044(0)='1' AND  B(17)='1' )then
          cVar2S5S110P023nsss(0) <='1';
          else
          cVar2S5S110P023nsss(0) <='0';
          end if;
        if(cVar1S6S110P000N051P053P044(0)='1' AND  B(17)='0' AND B(16)='1' )then
          cVar2S6S110N023P025nsss(0) <='1';
          else
          cVar2S6S110N023P025nsss(0) <='0';
          end if;
        if(cVar1S7S110P000N051P053N044(0)='1' AND  D(14)='0' AND B(17)='0' )then
          cVar2S7S110P042P023nsss(0) <='1';
          else
          cVar2S7S110P042P023nsss(0) <='0';
          end if;
        if(cVar1S8S110P000N051P053N044(0)='1' AND  D(14)='0' AND B(17)='1' AND E(22)='1' )then
          cVar2S8S110P042P023P045nsss(0) <='1';
          else
          cVar2S8S110P042P023P045nsss(0) <='0';
          end if;
        if(cVar1S9S110P000N051P053N044(0)='1' AND  D(14)='1' AND A(17)='1' )then
          cVar2S9S110P042P005nsss(0) <='1';
          else
          cVar2S9S110P042P005nsss(0) <='0';
          end if;
        if(cVar1S10S110P000N051P053P030(0)='1' AND  E( 9)='1' AND D( 8)='0' )then
          cVar2S10S110P064P066nsss(0) <='1';
          else
          cVar2S10S110P064P066nsss(0) <='0';
          end if;
        if(cVar1S11S110P000P030P027P060(0)='1' AND  E(11)='0' AND E(13)='0' )then
          cVar2S11S110P056P048nsss(0) <='1';
          else
          cVar2S11S110P056P048nsss(0) <='0';
          end if;
        if(cVar1S0S111P053P004P051P000(0)='1' AND  A(14)='1' AND E(16)='0' )then
          cVar2S0S111P011P069nsss(0) <='1';
          else
          cVar2S0S111P011P069nsss(0) <='0';
          end if;
        if(cVar1S1S111P053P004P051P000(0)='1' AND  A(14)='0' AND A(25)='1' )then
          cVar2S1S111N011P008nsss(0) <='1';
          else
          cVar2S1S111N011P008nsss(0) <='0';
          end if;
        if(cVar1S2S111P053P004P051P000(0)='1' AND  A(14)='0' AND A(25)='0' AND A(15)='1' )then
          cVar2S2S111N011N008P009nsss(0) <='1';
          else
          cVar2S2S111N011N008P009nsss(0) <='0';
          end if;
        if(cVar1S3S111P053P004N051P030(0)='1' AND  E( 9)='1' )then
          cVar2S3S111P064nsss(0) <='1';
          else
          cVar2S3S111P064nsss(0) <='0';
          end if;
        if(cVar1S4S111P053P004N051P030(0)='1' AND  E( 9)='0' AND D(18)='0' AND D(11)='0' )then
          cVar2S4S111N064P059P054nsss(0) <='1';
          else
          cVar2S4S111N064P059P054nsss(0) <='0';
          end if;
        if(cVar1S7S111N053P044N025N023(0)='1' AND  B(25)='0' AND B(27)='1' )then
          cVar2S7S111P026P022nsss(0) <='1';
          else
          cVar2S7S111P026P022nsss(0) <='0';
          end if;
        if(cVar1S8S111N053N044P042P023(0)='1' AND  E(11)='1' AND A(27)='0' AND D(23)='0' )then
          cVar2S8S111P056P004P039nsss(0) <='1';
          else
          cVar2S8S111P056P004P039nsss(0) <='0';
          end if;
        if(cVar1S9S111N053N044P042P023(0)='1' AND  E(11)='0' AND D(11)='0' AND B(27)='1' )then
          cVar2S9S111N056P054P022nsss(0) <='1';
          else
          cVar2S9S111N056P054P022nsss(0) <='0';
          end if;
        if(cVar1S10S111N053N044P042P023(0)='1' AND  E(22)='1' )then
          cVar2S10S111P045nsss(0) <='1';
          else
          cVar2S10S111P045nsss(0) <='0';
          end if;
        if(cVar1S11S111N053N044P042P023(0)='1' AND  E(22)='0' AND E( 9)='1' )then
          cVar2S11S111N045P064nsss(0) <='1';
          else
          cVar2S11S111N045P064nsss(0) <='0';
          end if;
        if(cVar1S13S111N053N044P042N005(0)='1' AND  A(15)='0' AND A(21)='0' AND A(20)='1' )then
          cVar2S13S111P009P016P018nsss(0) <='1';
          else
          cVar2S13S111P009P016P018nsss(0) <='0';
          end if;
        if(cVar1S2S112P044N023N025P032(0)='1' AND  A(29)='0' AND A(13)='0' AND D(10)='1' )then
          cVar2S2S112P000P013P058nsss(0) <='1';
          else
          cVar2S2S112P000P013P058nsss(0) <='0';
          end if;
        if(cVar1S3S112P044N023N025P032(0)='1' AND  A(29)='0' AND A(13)='1' AND D(16)='1' )then
          cVar2S3S112P000P013P067nsss(0) <='1';
          else
          cVar2S3S112P000P013P067nsss(0) <='0';
          end if;
        if(cVar1S4S112N044P042P023P051(0)='1' AND  E(23)='0' AND E(20)='1' AND A(29)='0' )then
          cVar2S4S112P041P053P000nsss(0) <='1';
          else
          cVar2S4S112P041P053P000nsss(0) <='0';
          end if;
        if(cVar1S5S112N044P042P023P051(0)='1' AND  E(23)='0' AND E(20)='0' AND E(16)='0' )then
          cVar2S5S112P041N053P069nsss(0) <='1';
          else
          cVar2S5S112P041N053P069nsss(0) <='0';
          end if;
        if(cVar1S6S112N044P042P023N051(0)='1' AND  E(20)='0' AND E(23)='1' AND B(28)='1' )then
          cVar2S6S112P053P041P020nsss(0) <='1';
          else
          cVar2S6S112P053P041P020nsss(0) <='0';
          end if;
        if(cVar1S7S112N044P042P023N051(0)='1' AND  E(20)='0' AND E(23)='0' AND D(23)='0' )then
          cVar2S7S112P053N041P039nsss(0) <='1';
          else
          cVar2S7S112P053N041P039nsss(0) <='0';
          end if;
        if(cVar1S8S112N044P042P023P024(0)='1' AND  E(22)='1' )then
          cVar2S8S112P045nsss(0) <='1';
          else
          cVar2S8S112P045nsss(0) <='0';
          end if;
        if(cVar1S9S112N044P042P023P024(0)='1' AND  E(22)='0' AND E( 9)='1' )then
          cVar2S9S112N045P064nsss(0) <='1';
          else
          cVar2S9S112N045P064nsss(0) <='0';
          end if;
        if(cVar1S10S112N044P042P024P062(0)='1' AND  D(17)='1' )then
          cVar2S10S112P063nsss(0) <='1';
          else
          cVar2S10S112P063nsss(0) <='0';
          end if;
        if(cVar1S11S112N044P042P024P062(0)='1' AND  D(17)='0' AND E( 8)='1' )then
          cVar2S11S112N063P068nsss(0) <='1';
          else
          cVar2S11S112N063P068nsss(0) <='0';
          end if;
        if(cVar1S2S113P044N025N023P032(0)='1' AND  A(29)='0' AND A(13)='0' )then
          cVar2S2S113P000P013nsss(0) <='1';
          else
          cVar2S2S113P000P013nsss(0) <='0';
          end if;
        if(cVar1S3S113N044P042P023P051(0)='1' AND  E(23)='0' AND E(20)='1' AND A(29)='0' )then
          cVar2S3S113P041P053P000nsss(0) <='1';
          else
          cVar2S3S113P041P053P000nsss(0) <='0';
          end if;
        if(cVar1S4S113N044P042P023P051(0)='1' AND  E(23)='0' AND E(20)='0' AND E(16)='0' )then
          cVar2S4S113P041N053P069nsss(0) <='1';
          else
          cVar2S4S113P041N053P069nsss(0) <='0';
          end if;
        if(cVar1S5S113N044P042P023N051(0)='1' AND  E(23)='1' AND B(28)='1' )then
          cVar2S5S113P041P020nsss(0) <='1';
          else
          cVar2S5S113P041P020nsss(0) <='0';
          end if;
        if(cVar1S6S113N044P042P023N051(0)='1' AND  E(23)='1' AND B(28)='0' AND A(21)='0' )then
          cVar2S6S113P041N020P016nsss(0) <='1';
          else
          cVar2S6S113P041N020P016nsss(0) <='0';
          end if;
        if(cVar1S7S113N044P042P023N051(0)='1' AND  E(23)='0' AND D(23)='0' AND A(21)='1' )then
          cVar2S7S113N041P039P016nsss(0) <='1';
          else
          cVar2S7S113N041P039P016nsss(0) <='0';
          end if;
        if(cVar1S8S113N044P042P023P024(0)='1' AND  E(22)='1' )then
          cVar2S8S113P045nsss(0) <='1';
          else
          cVar2S8S113P045nsss(0) <='0';
          end if;
        if(cVar1S9S113N044P042P023P024(0)='1' AND  E(22)='0' AND B(21)='0' AND B(11)='1' )then
          cVar2S9S113N045P034P035nsss(0) <='1';
          else
          cVar2S9S113N045P034P035nsss(0) <='0';
          end if;
        if(cVar1S10S113N044P042P024P062(0)='1' AND  D(17)='1' )then
          cVar2S10S113P063nsss(0) <='1';
          else
          cVar2S10S113P063nsss(0) <='0';
          end if;
        if(cVar1S11S113N044P042P024P062(0)='1' AND  D(17)='0' AND E( 8)='1' )then
          cVar2S11S113N063P068nsss(0) <='1';
          else
          cVar2S11S113N063P068nsss(0) <='0';
          end if;
        if(cVar1S2S114P016P044N023N025(0)='1' AND  B(25)='0' AND E(13)='0' AND B(27)='1' )then
          cVar2S2S114P026P048P022nsss(0) <='1';
          else
          cVar2S2S114P026P048P022nsss(0) <='0';
          end if;
        if(cVar1S4S114P016N044P041N020(0)='1' AND  D( 9)='0' AND E(18)='0' )then
          cVar2S4S114P062P061nsss(0) <='1';
          else
          cVar2S4S114P062P061nsss(0) <='0';
          end if;
        if(cVar1S5S114P016N044N041P020(0)='1' AND  A(27)='0' AND A(25)='1' AND A(11)='1' )then
          cVar2S5S114P004P008P017nsss(0) <='1';
          else
          cVar2S5S114P004P008P017nsss(0) <='0';
          end if;
        if(cVar1S6S114P016N044N041P020(0)='1' AND  A(27)='0' AND A(25)='0' AND D(21)='0' )then
          cVar2S6S114P004N008P047nsss(0) <='1';
          else
          cVar2S6S114P004N008P047nsss(0) <='0';
          end if;
        if(cVar1S7S114P016N044N041P020(0)='1' AND  A(27)='1' AND A(18)='0' AND A(26)='0' )then
          cVar2S7S114P004P003P006nsss(0) <='1';
          else
          cVar2S7S114P004P003P006nsss(0) <='0';
          end if;
        if(cVar1S8S114P016N044N041P020(0)='1' AND  E(15)='1' )then
          cVar2S8S114P040nsss(0) <='1';
          else
          cVar2S8S114P040nsss(0) <='0';
          end if;
        if(cVar1S9S114P016N044N041P020(0)='1' AND  E(15)='0' AND E( 9)='0' AND A(16)='1' )then
          cVar2S9S114N040P064P007nsss(0) <='1';
          else
          cVar2S9S114N040P064P007nsss(0) <='0';
          end if;
        if(cVar1S10S114P016P039P022P041(0)='1' AND  A(28)='0' AND A(12)='0' AND A(18)='1' )then
          cVar2S10S114P002P015P003nsss(0) <='1';
          else
          cVar2S10S114P002P015P003nsss(0) <='0';
          end if;
        if(cVar1S11S114P016P039P022P041(0)='1' AND  A(28)='1' AND D( 8)='1' AND E( 8)='0' )then
          cVar2S11S114P002P066P068nsss(0) <='1';
          else
          cVar2S11S114P002P066P068nsss(0) <='0';
          end if;
        if(cVar1S12S114P016P039P022P041(0)='1' AND  A(28)='1' AND D( 8)='0' AND A(15)='1' )then
          cVar2S12S114P002N066P009nsss(0) <='1';
          else
          cVar2S12S114P002N066P009nsss(0) <='0';
          end if;
        if(cVar1S13S114P016P039P022P041(0)='1' AND  E(16)='0' AND A(24)='0' AND A(23)='1' )then
          cVar2S13S114P069P010P012nsss(0) <='1';
          else
          cVar2S13S114P069P010P012nsss(0) <='0';
          end if;
        if(cVar1S14S114P016P039P022P019(0)='1' AND  A(20)='1' )then
          cVar2S14S114P018nsss(0) <='1';
          else
          cVar2S14S114P018nsss(0) <='0';
          end if;
        if(cVar1S16S114P016P039N005P069(0)='1' AND  B(21)='1' )then
          cVar2S16S114P034nsss(0) <='1';
          else
          cVar2S16S114P034nsss(0) <='0';
          end if;
        if(cVar1S2S115P044N025N023P032(0)='1' AND  A(29)='0' AND E(11)='0' AND A(26)='1' )then
          cVar2S2S115P000P056P006nsss(0) <='1';
          else
          cVar2S2S115P000P056P006nsss(0) <='0';
          end if;
        if(cVar1S3S115N044P042P023P008(0)='1' AND  B(13)='0' AND B(22)='0' )then
          cVar2S3S115P031P032nsss(0) <='1';
          else
          cVar2S3S115P031P032nsss(0) <='0';
          end if;
        if(cVar1S4S115N044P042P023P008(0)='1' AND  B(13)='0' AND B(22)='1' AND E( 8)='1' )then
          cVar2S4S115P031P032P068nsss(0) <='1';
          else
          cVar2S4S115P031P032P068nsss(0) <='0';
          end if;
        if(cVar1S5S115N044P042P023P008(0)='1' AND  B(13)='1' AND D(18)='1' )then
          cVar2S5S115P031P059nsss(0) <='1';
          else
          cVar2S5S115P031P059nsss(0) <='0';
          end if;
        if(cVar1S6S115N044P042P023N008(0)='1' AND  A(21)='1' AND B(27)='0' )then
          cVar2S6S115P016P022nsss(0) <='1';
          else
          cVar2S6S115P016P022nsss(0) <='0';
          end if;
        if(cVar1S7S115N044P042P023N008(0)='1' AND  A(21)='1' AND B(27)='1' AND A(20)='1' )then
          cVar2S7S115P016P022P018nsss(0) <='1';
          else
          cVar2S7S115P016P022P018nsss(0) <='0';
          end if;
        if(cVar1S8S115N044P042P023N008(0)='1' AND  A(21)='0' AND B(27)='1' AND D(22)='1' )then
          cVar2S8S115N016P022P043nsss(0) <='1';
          else
          cVar2S8S115N016P022P043nsss(0) <='0';
          end if;
        if(cVar1S9S115N044P042P023P024(0)='1' AND  A(26)='1' )then
          cVar2S9S115P006nsss(0) <='1';
          else
          cVar2S9S115P006nsss(0) <='0';
          end if;
        if(cVar1S10S115N044P042P023P024(0)='1' AND  A(26)='0' AND E(22)='1' )then
          cVar2S10S115N006P045nsss(0) <='1';
          else
          cVar2S10S115N006P045nsss(0) <='0';
          end if;
        if(cVar1S11S115N044P042P023P024(0)='1' AND  A(26)='0' AND E(22)='0' AND E( 9)='1' )then
          cVar2S11S115N006N045P064nsss(0) <='1';
          else
          cVar2S11S115N006N045P064nsss(0) <='0';
          end if;
        if(cVar1S13S115N044P042P024N005(0)='1' AND  A(15)='0' AND D( 9)='0' AND A(27)='1' )then
          cVar2S13S115P009P062P004nsss(0) <='1';
          else
          cVar2S13S115P009P062P004nsss(0) <='0';
          end if;
        if(cVar1S2S116P016P044N023N025(0)='1' AND  B(25)='0' AND E(13)='0' )then
          cVar2S2S116P026P048nsss(0) <='1';
          else
          cVar2S2S116P026P048nsss(0) <='0';
          end if;
        if(cVar1S4S116P016N044P041N020(0)='1' AND  D( 9)='0' AND E(18)='0' )then
          cVar2S4S116P062P061nsss(0) <='1';
          else
          cVar2S4S116P062P061nsss(0) <='0';
          end if;
        if(cVar1S5S116P016N044N041P004(0)='1' AND  A(24)='1' AND B(24)='1' AND A(22)='0' )then
          cVar2S5S116P010P028P014nsss(0) <='1';
          else
          cVar2S5S116P010P028P014nsss(0) <='0';
          end if;
        if(cVar1S6S116P016N044N041P004(0)='1' AND  A(24)='1' AND B(24)='0' AND D(23)='0' )then
          cVar2S6S116P010N028P039nsss(0) <='1';
          else
          cVar2S6S116P010N028P039nsss(0) <='0';
          end if;
        if(cVar1S7S116P016N044N041P004(0)='1' AND  A(24)='0' AND B(15)='1' AND A(22)='0' )then
          cVar2S7S116N010P027P014nsss(0) <='1';
          else
          cVar2S7S116N010P027P014nsss(0) <='0';
          end if;
        if(cVar1S8S116P016N044N041P004(0)='1' AND  A(24)='0' AND B(15)='0' AND B(28)='0' )then
          cVar2S8S116N010N027P020nsss(0) <='1';
          else
          cVar2S8S116N010N027P020nsss(0) <='0';
          end if;
        if(cVar1S9S116P016N044N041P004(0)='1' AND  A(18)='0' AND E(15)='1' )then
          cVar2S9S116P003P040nsss(0) <='1';
          else
          cVar2S9S116P003P040nsss(0) <='0';
          end if;
        if(cVar1S10S116P016P039P041P022(0)='1' AND  A(28)='0' AND A(12)='0' AND A(13)='1' )then
          cVar2S10S116P002P015P013nsss(0) <='1';
          else
          cVar2S10S116P002P015P013nsss(0) <='0';
          end if;
        if(cVar1S11S116P016P039P041P022(0)='1' AND  A(28)='1' AND D( 8)='1' AND D(16)='0' )then
          cVar2S11S116P002P066P067nsss(0) <='1';
          else
          cVar2S11S116P002P066P067nsss(0) <='0';
          end if;
        if(cVar1S12S116P016P039P041P022(0)='1' AND  A(28)='1' AND D( 8)='0' AND A(27)='1' )then
          cVar2S12S116P002N066P004nsss(0) <='1';
          else
          cVar2S12S116P002N066P004nsss(0) <='0';
          end if;
        if(cVar1S13S116P016P039P041P022(0)='1' AND  A(10)='1' AND A(14)='1' )then
          cVar2S13S116P019P011nsss(0) <='1';
          else
          cVar2S13S116P019P011nsss(0) <='0';
          end if;
        if(cVar1S14S116P016P039P041P069(0)='1' AND  A(24)='0' AND A(23)='1' )then
          cVar2S14S116P010P012nsss(0) <='1';
          else
          cVar2S14S116P010P012nsss(0) <='0';
          end if;
        if(cVar1S16S116P016P039N005P069(0)='1' AND  B(21)='1' )then
          cVar2S16S116P034nsss(0) <='1';
          else
          cVar2S16S116P034nsss(0) <='0';
          end if;
        if(cVar1S2S117P044N025N023P032(0)='1' AND  A(29)='0' AND E(11)='0' AND D(16)='1' )then
          cVar2S2S117P000P056P067nsss(0) <='1';
          else
          cVar2S2S117P000P056P067nsss(0) <='0';
          end if;
        if(cVar1S3S117N044P023P042P002(0)='1' AND  A(17)='0' AND D(23)='0' AND B(14)='1' )then
          cVar2S3S117P005P039P029nsss(0) <='1';
          else
          cVar2S3S117P005P039P029nsss(0) <='0';
          end if;
        if(cVar1S4S117N044P023P042P002(0)='1' AND  A(17)='0' AND D(23)='1' AND A(18)='1' )then
          cVar2S4S117P005P039P003nsss(0) <='1';
          else
          cVar2S4S117P005P039P003nsss(0) <='0';
          end if;
        if(cVar1S5S117N044P023P042P002(0)='1' AND  A(17)='1' AND B(13)='0' AND B(28)='1' )then
          cVar2S5S117P005P031P020nsss(0) <='1';
          else
          cVar2S5S117P005P031P020nsss(0) <='0';
          end if;
        if(cVar1S6S117N044P023P042P002(0)='1' AND  D(15)='1' )then
          cVar2S6S117P038nsss(0) <='1';
          else
          cVar2S6S117P038nsss(0) <='0';
          end if;
        if(cVar1S7S117N044P023P042P002(0)='1' AND  D(15)='0' AND D(11)='0' AND B(23)='1' )then
          cVar2S7S117N038P054P030nsss(0) <='1';
          else
          cVar2S7S117N038P054P030nsss(0) <='0';
          end if;
        if(cVar1S8S117N044P023P042P024(0)='1' AND  A(28)='1' )then
          cVar2S8S117P002nsss(0) <='1';
          else
          cVar2S8S117P002nsss(0) <='0';
          end if;
        if(cVar1S9S117N044P023P042P024(0)='1' AND  A(28)='0' AND E(16)='1' )then
          cVar2S9S117N002P069nsss(0) <='1';
          else
          cVar2S9S117N002P069nsss(0) <='0';
          end if;
        if(cVar1S10S117N044P023P042P024(0)='1' AND  A(28)='0' AND E(16)='0' AND E( 9)='1' )then
          cVar2S10S117N002N069P064nsss(0) <='1';
          else
          cVar2S10S117N002N069P064nsss(0) <='0';
          end if;
        if(cVar1S12S117N044P023P024N005(0)='1' AND  E( 8)='1' )then
          cVar2S12S117P068nsss(0) <='1';
          else
          cVar2S12S117P068nsss(0) <='0';
          end if;
        if(cVar1S2S118P044N025N023P032(0)='1' AND  A(29)='0' AND E(11)='0' )then
          cVar2S2S118P000P056nsss(0) <='1';
          else
          cVar2S2S118P000P056nsss(0) <='0';
          end if;
        if(cVar1S3S118N044P023P042P002(0)='1' AND  A(17)='0' AND D(23)='0' )then
          cVar2S3S118P005P039nsss(0) <='1';
          else
          cVar2S3S118P005P039nsss(0) <='0';
          end if;
        if(cVar1S4S118N044P023P042P002(0)='1' AND  A(17)='0' AND D(23)='1' AND A(18)='1' )then
          cVar2S4S118P005P039P003nsss(0) <='1';
          else
          cVar2S4S118P005P039P003nsss(0) <='0';
          end if;
        if(cVar1S5S118N044P023P042P002(0)='1' AND  A(17)='1' AND B(13)='0' AND E(23)='1' )then
          cVar2S5S118P005P031P041nsss(0) <='1';
          else
          cVar2S5S118P005P031P041nsss(0) <='0';
          end if;
        if(cVar1S6S118N044P023P042P002(0)='1' AND  D(15)='1' )then
          cVar2S6S118P038nsss(0) <='1';
          else
          cVar2S6S118P038nsss(0) <='0';
          end if;
        if(cVar1S7S118N044P023P042P024(0)='1' AND  A(28)='1' )then
          cVar2S7S118P002nsss(0) <='1';
          else
          cVar2S7S118P002nsss(0) <='0';
          end if;
        if(cVar1S8S118N044P023P042P024(0)='1' AND  A(28)='0' AND E(16)='1' )then
          cVar2S8S118N002P069nsss(0) <='1';
          else
          cVar2S8S118N002P069nsss(0) <='0';
          end if;
        if(cVar1S9S118N044P023P042P024(0)='1' AND  A(28)='0' AND E(16)='0' AND A(18)='1' )then
          cVar2S9S118N002N069P003nsss(0) <='1';
          else
          cVar2S9S118N002N069P003nsss(0) <='0';
          end if;
        if(cVar1S11S118N044P023P024N005(0)='1' AND  E( 8)='1' )then
          cVar2S11S118P068nsss(0) <='1';
          else
          cVar2S11S118P068nsss(0) <='0';
          end if;
        if(cVar1S2S119P044N025N023P000(0)='1' AND  B(22)='0' AND A(13)='0' AND D(10)='1' )then
          cVar2S2S119P032P013P058nsss(0) <='1';
          else
          cVar2S2S119P032P013P058nsss(0) <='0';
          end if;
        if(cVar1S3S119N044P023P042P053(0)='1' AND  A(27)='0' AND D(20)='1' )then
          cVar2S3S119P004P051nsss(0) <='1';
          else
          cVar2S3S119P004P051nsss(0) <='0';
          end if;
        if(cVar1S4S119N044P023P042N053(0)='1' AND  D(20)='0' AND E(23)='1' AND B(28)='1' )then
          cVar2S4S119P051P041P020nsss(0) <='1';
          else
          cVar2S4S119P051P041P020nsss(0) <='0';
          end if;
        if(cVar1S5S119N044P023P042P024(0)='1' AND  A(28)='1' )then
          cVar2S5S119P002nsss(0) <='1';
          else
          cVar2S5S119P002nsss(0) <='0';
          end if;
        if(cVar1S6S119N044P023P042P024(0)='1' AND  A(28)='0' AND D(17)='1' )then
          cVar2S6S119N002P063nsss(0) <='1';
          else
          cVar2S6S119N002P063nsss(0) <='0';
          end if;
        if(cVar1S7S119N044P023P042P024(0)='1' AND  A(28)='0' AND D(17)='0' AND E(16)='1' )then
          cVar2S7S119N002N063P069nsss(0) <='1';
          else
          cVar2S7S119N002N063P069nsss(0) <='0';
          end if;
        if(cVar1S9S119N044P023P024N008(0)='1' AND  E(16)='0' AND B(20)='1' )then
          cVar2S9S119P069P036nsss(0) <='1';
          else
          cVar2S9S119P069P036nsss(0) <='0';
          end if;
        if(cVar1S10S119N044P023P024N008(0)='1' AND  E(16)='0' AND B(20)='0' AND E( 8)='1' )then
          cVar2S10S119P069N036P068nsss(0) <='1';
          else
          cVar2S10S119P069N036P068nsss(0) <='0';
          end if;
        if(cVar1S2S120P044N025N023P000(0)='1' AND  B(22)='0' AND A(13)='0' )then
          cVar2S2S120P032P013nsss(0) <='1';
          else
          cVar2S2S120P032P013nsss(0) <='0';
          end if;
        if(cVar1S3S120N044P023P042P054(0)='1' AND  E(11)='0' AND B(23)='0' AND E(19)='0' )then
          cVar2S3S120P056P030P057nsss(0) <='1';
          else
          cVar2S3S120P056P030P057nsss(0) <='0';
          end if;
        if(cVar1S4S120N044P023P042P054(0)='1' AND  E(11)='1' AND D(10)='1' )then
          cVar2S4S120P056P058nsss(0) <='1';
          else
          cVar2S4S120P056P058nsss(0) <='0';
          end if;
        if(cVar1S5S120N044P023P042P054(0)='1' AND  E(11)='1' AND A(27)='0' )then
          cVar2S5S120P056P004nsss(0) <='1';
          else
          cVar2S5S120P056P004nsss(0) <='0';
          end if;
        if(cVar1S6S120N044P023P042P024(0)='1' AND  D( 9)='0' AND E(17)='1' )then
          cVar2S6S120P062P065nsss(0) <='1';
          else
          cVar2S6S120P062P065nsss(0) <='0';
          end if;
        if(cVar1S7S120N044P023P042P024(0)='1' AND  D( 9)='0' AND E(17)='0' AND E( 8)='1' )then
          cVar2S7S120P062N065P068nsss(0) <='1';
          else
          cVar2S7S120P062N065P068nsss(0) <='0';
          end if;
        if(cVar1S9S120N044P023P024N005(0)='1' AND  E( 8)='1' )then
          cVar2S9S120P068nsss(0) <='1';
          else
          cVar2S9S120P068nsss(0) <='0';
          end if;
        if(cVar1S3S121P042N023N002N055(0)='1' AND  A(26)='1' AND E(14)='1' )then
          cVar2S3S121P006P044nsss(0) <='1';
          else
          cVar2S3S121P006P044nsss(0) <='0';
          end if;
        if(cVar1S4S121P042N023N002N055(0)='1' AND  A(26)='0' AND B(26)='0' AND E(17)='1' )then
          cVar2S4S121N006P024P065nsss(0) <='1';
          else
          cVar2S4S121N006P024P065nsss(0) <='0';
          end if;
        if(cVar1S5S121N042P023P052P065(0)='1' AND  B(20)='0' )then
          cVar2S5S121P036nsss(0) <='1';
          else
          cVar2S5S121P036nsss(0) <='0';
          end if;
        if(cVar1S6S121N042P023P052N065(0)='1' AND  D( 9)='1' )then
          cVar2S6S121P062nsss(0) <='1';
          else
          cVar2S6S121P062nsss(0) <='0';
          end if;
        if(cVar1S7S121N042P023P052N065(0)='1' AND  D( 9)='0' AND D(12)='1' AND A(13)='0' )then
          cVar2S7S121N062P050P013nsss(0) <='1';
          else
          cVar2S7S121N062P050P013nsss(0) <='0';
          end if;
        if(cVar1S8S121N042P023P052N065(0)='1' AND  D( 9)='0' AND D(12)='0' AND E(20)='1' )then
          cVar2S8S121N062N050P053nsss(0) <='1';
          else
          cVar2S8S121N062N050P053nsss(0) <='0';
          end if;
        if(cVar1S9S121N042P023N052P050(0)='1' AND  D(13)='1' AND B(16)='1' )then
          cVar2S9S121P046P025nsss(0) <='1';
          else
          cVar2S9S121P046P025nsss(0) <='0';
          end if;
        if(cVar1S10S121N042P023N052P050(0)='1' AND  D(13)='0' AND B(16)='1' AND E(22)='1' )then
          cVar2S10S121N046P025P045nsss(0) <='1';
          else
          cVar2S10S121N046P025P045nsss(0) <='0';
          end if;
        if(cVar1S11S121N042P023N052P050(0)='1' AND  A(27)='0' AND D(17)='0' AND E(13)='1' )then
          cVar2S11S121P004P063P048nsss(0) <='1';
          else
          cVar2S11S121P004P063P048nsss(0) <='0';
          end if;
        if(cVar1S13S121N042P023P024N008(0)='1' AND  E(16)='0' AND B(20)='1' )then
          cVar2S13S121P069P036nsss(0) <='1';
          else
          cVar2S13S121P069P036nsss(0) <='0';
          end if;
        if(cVar1S14S121N042P023P024N008(0)='1' AND  E(16)='0' AND B(20)='0' AND E( 8)='1' )then
          cVar2S14S121P069N036P068nsss(0) <='1';
          else
          cVar2S14S121P069N036P068nsss(0) <='0';
          end if;
        if(cVar1S1S122P044P026N025P000(0)='1' AND  B(17)='1' )then
          cVar2S1S122P023nsss(0) <='1';
          else
          cVar2S1S122P023nsss(0) <='0';
          end if;
        if(cVar1S2S122P044P026N025P000(0)='1' AND  B(17)='0' AND B(22)='0' AND D(16)='1' )then
          cVar2S2S122N023P032P067nsss(0) <='1';
          else
          cVar2S2S122N023P032P067nsss(0) <='0';
          end if;
        if(cVar1S3S122N044P023P042P020(0)='1' AND  D(23)='1' )then
          cVar2S3S122P039nsss(0) <='1';
          else
          cVar2S3S122P039nsss(0) <='0';
          end if;
        if(cVar1S4S122N044P023P042P020(0)='1' AND  D(23)='0' AND D( 9)='0' AND A(25)='0' )then
          cVar2S4S122N039P062P008nsss(0) <='1';
          else
          cVar2S4S122N039P062P008nsss(0) <='0';
          end if;
        if(cVar1S5S122N044P023P042P020(0)='1' AND  D(23)='0' AND D( 9)='1' AND A(22)='1' )then
          cVar2S5S122N039P062P014nsss(0) <='1';
          else
          cVar2S5S122N039P062P014nsss(0) <='0';
          end if;
        if(cVar1S6S122N044P023P042N020(0)='1' AND  D(23)='0' AND D(18)='1' AND A(27)='0' )then
          cVar2S6S122P039P059P004nsss(0) <='1';
          else
          cVar2S6S122P039P059P004nsss(0) <='0';
          end if;
        if(cVar1S7S122N044P023P042N020(0)='1' AND  D(23)='0' AND D(18)='0' AND E(18)='0' )then
          cVar2S7S122P039N059P061nsss(0) <='1';
          else
          cVar2S7S122P039N059P061nsss(0) <='0';
          end if;
        if(cVar1S8S122N044P023P042N020(0)='1' AND  D(23)='1' AND A(23)='0' AND D(12)='0' )then
          cVar2S8S122P039P012P050nsss(0) <='1';
          else
          cVar2S8S122P039P012P050nsss(0) <='0';
          end if;
        if(cVar1S9S122N044P023P042P024(0)='1' AND  D( 9)='0' AND D(17)='1' )then
          cVar2S9S122P062P063nsss(0) <='1';
          else
          cVar2S9S122P062P063nsss(0) <='0';
          end if;
        if(cVar1S10S122N044P023P042P024(0)='1' AND  D( 9)='0' AND D(17)='0' AND A(18)='1' )then
          cVar2S10S122P062N063P003nsss(0) <='1';
          else
          cVar2S10S122P062N063P003nsss(0) <='0';
          end if;
        if(cVar1S12S122N044P023P024N006(0)='1' AND  E(22)='1' )then
          cVar2S12S122P045nsss(0) <='1';
          else
          cVar2S12S122P045nsss(0) <='0';
          end if;
        if(cVar1S13S122N044P023P024N006(0)='1' AND  E(22)='0' AND E(16)='0' AND A(22)='1' )then
          cVar2S13S122N045P069P014nsss(0) <='1';
          else
          cVar2S13S122N045P069P014nsss(0) <='0';
          end if;
        if(cVar1S3S123P042N023N002N055(0)='1' AND  A(26)='1' AND E(14)='1' )then
          cVar2S3S123P006P044nsss(0) <='1';
          else
          cVar2S3S123P006P044nsss(0) <='0';
          end if;
        if(cVar1S4S123P042N023N002N055(0)='1' AND  A(26)='0' AND B(26)='0' AND E(17)='1' )then
          cVar2S4S123N006P024P065nsss(0) <='1';
          else
          cVar2S4S123N006P024P065nsss(0) <='0';
          end if;
        if(cVar1S5S123N042P023P019P006(0)='1' AND  D(16)='0' AND E(16)='0' )then
          cVar2S5S123P067P069nsss(0) <='1';
          else
          cVar2S5S123P067P069nsss(0) <='0';
          end if;
        if(cVar1S6S123N042P023P019P006(0)='1' AND  D(16)='0' AND E(16)='1' AND A(22)='0' )then
          cVar2S6S123P067P069P014nsss(0) <='1';
          else
          cVar2S6S123P067P069P014nsss(0) <='0';
          end if;
        if(cVar1S7S123N042P023P019P006(0)='1' AND  D(16)='1' AND B(26)='0' AND D(19)='1' )then
          cVar2S7S123P067P024P055nsss(0) <='1';
          else
          cVar2S7S123P067P024P055nsss(0) <='0';
          end if;
        if(cVar1S8S123N042P023P019P006(0)='1' AND  D(13)='1' )then
          cVar2S8S123P046nsss(0) <='1';
          else
          cVar2S8S123P046nsss(0) <='0';
          end if;
        if(cVar1S9S123N042P023N019P069(0)='1' AND  E(22)='0' AND B(14)='1' )then
          cVar2S9S123P045P029nsss(0) <='1';
          else
          cVar2S9S123P045P029nsss(0) <='0';
          end if;
        if(cVar1S10S123N042P023N019P069(0)='1' AND  E(22)='0' AND B(14)='0' AND A(15)='0' )then
          cVar2S10S123P045N029P009nsss(0) <='1';
          else
          cVar2S10S123P045N029P009nsss(0) <='0';
          end if;
        if(cVar1S11S123N042P023N019N069(0)='1' AND  D(20)='1' AND A(14)='1' )then
          cVar2S11S123P051P011nsss(0) <='1';
          else
          cVar2S11S123P051P011nsss(0) <='0';
          end if;
        if(cVar1S12S123N042P023N019N069(0)='1' AND  D(20)='1' AND A(14)='0' AND A(24)='1' )then
          cVar2S12S123P051N011P010nsss(0) <='1';
          else
          cVar2S12S123P051N011P010nsss(0) <='0';
          end if;
        if(cVar1S13S123N042P023N019N069(0)='1' AND  D(20)='0' AND D(15)='1' AND E(15)='1' )then
          cVar2S13S123N051P038P040nsss(0) <='1';
          else
          cVar2S13S123N051P038P040nsss(0) <='0';
          end if;
        if(cVar1S15S123N042P023P024N007(0)='1' AND  A(17)='1' )then
          cVar2S15S123P005nsss(0) <='1';
          else
          cVar2S15S123P005nsss(0) <='0';
          end if;
        if(cVar1S0S124P019P018P067P039(0)='1' AND  A(18)='1' )then
          cVar2S0S124P003nsss(0) <='1';
          else
          cVar2S0S124P003nsss(0) <='0';
          end if;
        if(cVar1S1S124P019P018P067P039(0)='1' AND  A(18)='0' AND B(28)='1' )then
          cVar2S1S124N003P020nsss(0) <='1';
          else
          cVar2S1S124N003P020nsss(0) <='0';
          end if;
        if(cVar1S2S124P019P018P067P039(0)='1' AND  A(18)='0' AND B(28)='0' AND A(13)='1' )then
          cVar2S2S124N003N020P013nsss(0) <='1';
          else
          cVar2S2S124N003N020P013nsss(0) <='0';
          end if;
        if(cVar1S3S124P019P018P067N039(0)='1' AND  D(17)='1' AND D(10)='1' )then
          cVar2S3S124P063P058nsss(0) <='1';
          else
          cVar2S3S124P063P058nsss(0) <='0';
          end if;
        if(cVar1S4S124P019P018P067N039(0)='1' AND  D(17)='1' AND D(10)='0' AND A(19)='0' )then
          cVar2S4S124P063N058P001nsss(0) <='1';
          else
          cVar2S4S124P063N058P001nsss(0) <='0';
          end if;
        if(cVar1S5S124P019P018P067N039(0)='1' AND  D(17)='0' AND E(17)='0' )then
          cVar2S5S124N063P065nsss(0) <='1';
          else
          cVar2S5S124N063P065nsss(0) <='0';
          end if;
        if(cVar1S6S124P019P018P067P028(0)='1' AND  A(26)='0' AND B(18)='0' AND E(14)='1' )then
          cVar2S6S124P006P021P044nsss(0) <='1';
          else
          cVar2S6S124P006P021P044nsss(0) <='0';
          end if;
        if(cVar1S7S124P019P018P067P028(0)='1' AND  A(26)='1' AND A(23)='0' AND A(22)='1' )then
          cVar2S7S124P006P012P014nsss(0) <='1';
          else
          cVar2S7S124P006P012P014nsss(0) <='0';
          end if;
        if(cVar1S8S124P019P018P039P033(0)='1' AND  A(16)='0' AND A(12)='0' )then
          cVar2S8S124P007P015nsss(0) <='1';
          else
          cVar2S8S124P007P015nsss(0) <='0';
          end if;
        if(cVar1S9S124P019P018P039P033(0)='1' AND  A(16)='0' AND A(12)='1' AND A(22)='0' )then
          cVar2S9S124P007P015P014nsss(0) <='1';
          else
          cVar2S9S124P007P015P014nsss(0) <='0';
          end if;
        if(cVar1S10S124P019P018P039N033(0)='1' AND  A(26)='1' AND D( 8)='0' )then
          cVar2S10S124P006P066nsss(0) <='1';
          else
          cVar2S10S124P006P066nsss(0) <='0';
          end if;
        if(cVar1S11S124P019P018P039N033(0)='1' AND  A(26)='0' AND A(15)='1' AND E(17)='0' )then
          cVar2S11S124N006P009P065nsss(0) <='1';
          else
          cVar2S11S124N006P009P065nsss(0) <='0';
          end if;
        if(cVar1S12S124P019P018P039P017(0)='1' AND  A(21)='0' )then
          cVar2S12S124P016nsss(0) <='1';
          else
          cVar2S12S124P016nsss(0) <='0';
          end if;
        if(cVar1S14S124P019P051P042N067(0)='1' AND  B(10)='1' )then
          cVar2S14S124P037nsss(0) <='1';
          else
          cVar2S14S124P037nsss(0) <='0';
          end if;
        if(cVar1S15S124P019P051P042N067(0)='1' AND  B(10)='0' AND A(12)='1' )then
          cVar2S15S124N037P015nsss(0) <='1';
          else
          cVar2S15S124N037P015nsss(0) <='0';
          end if;
        if(cVar1S16S124P019P051N042P029(0)='1' AND  A(13)='0' AND E(13)='0' AND A(17)='1' )then
          cVar2S16S124P013P048P005nsss(0) <='1';
          else
          cVar2S16S124P013P048P005nsss(0) <='0';
          end if;
        if(cVar1S17S124P019P051N042P029(0)='1' AND  A(13)='0' AND E(13)='1' AND A(21)='0' )then
          cVar2S17S124P013P048P016nsss(0) <='1';
          else
          cVar2S17S124P013P048P016nsss(0) <='0';
          end if;
        if(cVar1S18S124P019P051N042P029(0)='1' AND  A(24)='1' )then
          cVar2S18S124P010nsss(0) <='1';
          else
          cVar2S18S124P010nsss(0) <='0';
          end if;
        if(cVar1S19S124P019P051N042P029(0)='1' AND  A(24)='0' AND D(16)='0' AND A(13)='1' )then
          cVar2S19S124N010P067P013nsss(0) <='1';
          else
          cVar2S19S124N010P067P013nsss(0) <='0';
          end if;
        if(cVar1S20S124P019P051P037P024(0)='1' AND  E(18)='1' )then
          cVar2S20S124P061nsss(0) <='1';
          else
          cVar2S20S124P061nsss(0) <='0';
          end if;
        if(cVar1S21S124P019P051P037P024(0)='1' AND  E(18)='0' AND A(11)='1' AND A(22)='0' )then
          cVar2S21S124N061P017P014nsss(0) <='1';
          else
          cVar2S21S124N061P017P014nsss(0) <='0';
          end if;
        if(cVar1S22S124P019P051N037P000(0)='1' AND  B(25)='1' )then
          cVar2S22S124P026nsss(0) <='1';
          else
          cVar2S22S124P026nsss(0) <='0';
          end if;
        if(cVar1S23S124P019P051N037P000(0)='1' AND  B(25)='0' AND A(11)='0' AND A(22)='1' )then
          cVar2S23S124N026P017P014nsss(0) <='1';
          else
          cVar2S23S124N026P017P014nsss(0) <='0';
          end if;
        if(cVar1S0S125P018P050P029P032(0)='1' AND  E(18)='1' AND B(12)='1' )then
          cVar2S0S125P061P033nsss(0) <='1';
          else
          cVar2S0S125P061P033nsss(0) <='0';
          end if;
        if(cVar1S1S125P018P050P029P032(0)='1' AND  E(18)='1' AND B(12)='0' AND E( 9)='0' )then
          cVar2S1S125P061N033P064nsss(0) <='1';
          else
          cVar2S1S125P061N033P064nsss(0) <='0';
          end if;
        if(cVar1S2S125P018P050P029P032(0)='1' AND  E(18)='0' AND D(18)='0' )then
          cVar2S2S125N061P059nsss(0) <='1';
          else
          cVar2S2S125N061P059nsss(0) <='0';
          end if;
        if(cVar1S3S125P018P050P029P032(0)='1' AND  A(13)='1' AND A(22)='0' )then
          cVar2S3S125P013P014nsss(0) <='1';
          else
          cVar2S3S125P013P014nsss(0) <='0';
          end if;
        if(cVar1S4S125P018P050P029P032(0)='1' AND  A(13)='1' AND A(22)='1' AND A(21)='1' )then
          cVar2S4S125P013P014P016nsss(0) <='1';
          else
          cVar2S4S125P013P014P016nsss(0) <='0';
          end if;
        if(cVar1S5S125P018P050P029P011(0)='1' AND  A(21)='0' )then
          cVar2S5S125P016nsss(0) <='1';
          else
          cVar2S5S125P016nsss(0) <='0';
          end if;
        if(cVar1S6S125P018P050P029N011(0)='1' AND  A(13)='1' )then
          cVar2S6S125P013nsss(0) <='1';
          else
          cVar2S6S125P013nsss(0) <='0';
          end if;
        if(cVar1S7S125P018P050P004P012(0)='1' AND  E(11)='0' AND B(21)='1' )then
          cVar2S7S125P056P034nsss(0) <='1';
          else
          cVar2S7S125P056P034nsss(0) <='0';
          end if;
        if(cVar1S8S125P018P050P004P012(0)='1' AND  E(11)='0' AND B(21)='0' AND A(21)='0' )then
          cVar2S8S125P056N034P016nsss(0) <='1';
          else
          cVar2S8S125P056N034P016nsss(0) <='0';
          end if;
        if(cVar1S9S125P018P050P004P012(0)='1' AND  A(21)='1' AND A(24)='1' )then
          cVar2S9S125P016P010nsss(0) <='1';
          else
          cVar2S9S125P016P010nsss(0) <='0';
          end if;
        if(cVar1S10S125N018P039P054P034(0)='1' AND  B(28)='1' )then
          cVar2S10S125P020nsss(0) <='1';
          else
          cVar2S10S125P020nsss(0) <='0';
          end if;
        if(cVar1S11S125N018P039P054P034(0)='1' AND  B(28)='0' AND A(23)='0' )then
          cVar2S11S125N020P012nsss(0) <='1';
          else
          cVar2S11S125N020P012nsss(0) <='0';
          end if;
        if(cVar1S12S125N018N039P014P060(0)='1' AND  B(22)='1' )then
          cVar2S12S125P032nsss(0) <='1';
          else
          cVar2S12S125P032nsss(0) <='0';
          end if;
        if(cVar1S13S125N018N039P014P060(0)='1' AND  B(22)='0' AND B(21)='1' )then
          cVar2S13S125N032P034nsss(0) <='1';
          else
          cVar2S13S125N032P034nsss(0) <='0';
          end if;
        if(cVar1S14S125N018N039P014P060(0)='1' AND  B(22)='0' AND B(21)='0' AND A(21)='0' )then
          cVar2S14S125N032N034P016nsss(0) <='1';
          else
          cVar2S14S125N032N034P016nsss(0) <='0';
          end if;
        if(cVar1S15S125N018N039P014N060(0)='1' AND  E(14)='0' AND D(11)='0' AND B(13)='0' )then
          cVar2S15S125P044P054P031nsss(0) <='1';
          else
          cVar2S15S125P044P054P031nsss(0) <='0';
          end if;
        if(cVar1S16S125N018N039P014N060(0)='1' AND  E(14)='0' AND D(11)='1' AND E(17)='1' )then
          cVar2S16S125P044P054P065nsss(0) <='1';
          else
          cVar2S16S125P044P054P065nsss(0) <='0';
          end if;
        if(cVar1S17S125N018N039N014P044(0)='1' AND  D( 9)='0' )then
          cVar2S17S125P062nsss(0) <='1';
          else
          cVar2S17S125P062nsss(0) <='0';
          end if;
        if(cVar1S18S125N018N039N014N044(0)='1' AND  D(14)='0' AND B(23)='1' AND A(23)='1' )then
          cVar2S18S125P042P030P012nsss(0) <='1';
          else
          cVar2S18S125P042P030P012nsss(0) <='0';
          end if;
        if(cVar1S19S125N018N039N014N044(0)='1' AND  D(14)='0' AND B(23)='0' AND B(24)='1' )then
          cVar2S19S125P042N030P028nsss(0) <='1';
          else
          cVar2S19S125P042N030P028nsss(0) <='0';
          end if;
        if(cVar1S20S125N018N039N014N044(0)='1' AND  D(14)='1' AND E(15)='1' )then
          cVar2S20S125P042P040nsss(0) <='1';
          else
          cVar2S20S125P042P040nsss(0) <='0';
          end if;
        if(cVar1S0S126P018P014P037P004(0)='1' AND  D(14)='1' )then
          cVar2S0S126P042nsss(0) <='1';
          else
          cVar2S0S126P042nsss(0) <='0';
          end if;
        if(cVar1S1S126P018P014P037P004(0)='1' AND  D(14)='0' AND A(13)='1' AND A(14)='0' )then
          cVar2S1S126N042P013P011nsss(0) <='1';
          else
          cVar2S1S126N042P013P011nsss(0) <='0';
          end if;
        if(cVar1S2S126P018P014P037P004(0)='1' AND  D(14)='0' AND A(13)='0' AND A(12)='0' )then
          cVar2S2S126N042N013P015nsss(0) <='1';
          else
          cVar2S2S126N042N013P015nsss(0) <='0';
          end if;
        if(cVar1S3S126P018P014P037N004(0)='1' AND  B(23)='1' AND D(18)='1' )then
          cVar2S3S126P030P059nsss(0) <='1';
          else
          cVar2S3S126P030P059nsss(0) <='0';
          end if;
        if(cVar1S4S126P018P014P037N004(0)='1' AND  B(23)='1' AND D(18)='0' AND B(13)='0' )then
          cVar2S4S126P030N059P031nsss(0) <='1';
          else
          cVar2S4S126P030N059P031nsss(0) <='0';
          end if;
        if(cVar1S5S126P018P014P037N004(0)='1' AND  B(23)='0' AND D(19)='0' AND A(11)='0' )then
          cVar2S5S126N030P055P017nsss(0) <='1';
          else
          cVar2S5S126N030P055P017nsss(0) <='0';
          end if;
        if(cVar1S6S126P018P014P037N004(0)='1' AND  B(23)='0' AND D(19)='1' AND D(17)='1' )then
          cVar2S6S126N030P055P063nsss(0) <='1';
          else
          cVar2S6S126N030P055P063nsss(0) <='0';
          end if;
        if(cVar1S7S126P018P014P037P016(0)='1' AND  A(26)='0' AND D( 9)='1' AND E( 9)='1' )then
          cVar2S7S126P006P062P064nsss(0) <='1';
          else
          cVar2S7S126P006P062P064nsss(0) <='0';
          end if;
        if(cVar1S8S126P018P014P037P016(0)='1' AND  A(26)='0' AND D( 9)='0' )then
          cVar2S8S126P006N062psss(0) <='1';
          else
          cVar2S8S126P006N062psss(0) <='0';
          end if;
        if(cVar1S9S126P018P014P037N016(0)='1' AND  B(20)='0' AND A(26)='1' AND A(10)='1' )then
          cVar2S9S126P036P006P019nsss(0) <='1';
          else
          cVar2S9S126P036P006P019nsss(0) <='0';
          end if;
        if(cVar1S10S126P018P014P037N016(0)='1' AND  B(20)='0' AND A(26)='0' AND D(19)='1' )then
          cVar2S10S126P036N006P055nsss(0) <='1';
          else
          cVar2S10S126P036N006P055nsss(0) <='0';
          end if;
        if(cVar1S12S126P018P014P060N032(0)='1' AND  B(21)='1' )then
          cVar2S12S126P034nsss(0) <='1';
          else
          cVar2S12S126P034nsss(0) <='0';
          end if;
        if(cVar1S13S126P018P014P060N032(0)='1' AND  B(21)='0' AND A(21)='0' AND D(16)='0' )then
          cVar2S13S126N034P016P067nsss(0) <='1';
          else
          cVar2S13S126N034P016P067nsss(0) <='0';
          end if;
        if(cVar1S14S126P018P014P060N032(0)='1' AND  B(21)='0' AND A(21)='1' AND A(11)='1' )then
          cVar2S14S126N034P016P017nsss(0) <='1';
          else
          cVar2S14S126N034P016P017nsss(0) <='0';
          end if;
        if(cVar1S15S126P018P014N060P044(0)='1' AND  D(13)='0' AND B(15)='0' AND A(11)='1' )then
          cVar2S15S126P046P027P017nsss(0) <='1';
          else
          cVar2S15S126P046P027P017nsss(0) <='0';
          end if;
        if(cVar1S17S126P018P061N033P048(0)='1' AND  A(14)='1' AND D(16)='0' )then
          cVar2S17S126P011P067nsss(0) <='1';
          else
          cVar2S17S126P011P067nsss(0) <='0';
          end if;
        if(cVar1S18S126P018P061N033P048(0)='1' AND  A(14)='0' AND B(11)='1' AND D( 9)='0' )then
          cVar2S18S126N011P035P062nsss(0) <='1';
          else
          cVar2S18S126N011P035P062nsss(0) <='0';
          end if;
        if(cVar1S19S126P018P061N033P048(0)='1' AND  A(14)='0' AND B(11)='0' AND B(20)='1' )then
          cVar2S19S126N011N035P036nsss(0) <='1';
          else
          cVar2S19S126N011N035P036nsss(0) <='0';
          end if;
        if(cVar1S21S126P018N061P042N063(0)='1' AND  A(24)='0' AND A(21)='0' AND A(22)='0' )then
          cVar2S21S126P010P016P014nsss(0) <='1';
          else
          cVar2S21S126P010P016P014nsss(0) <='0';
          end if;
        if(cVar1S22S126P018N061P042N063(0)='1' AND  A(24)='0' AND A(21)='1' AND A(12)='0' )then
          cVar2S22S126P010P016P015nsss(0) <='1';
          else
          cVar2S22S126P010P016P015nsss(0) <='0';
          end if;
        if(cVar1S23S126P018N061N042P050(0)='1' AND  A(19)='1' AND A(15)='0' )then
          cVar2S23S126P001P009nsss(0) <='1';
          else
          cVar2S23S126P001P009nsss(0) <='0';
          end if;
        if(cVar1S24S126P018N061N042P050(0)='1' AND  A(19)='0' AND B(17)='0' AND A(18)='1' )then
          cVar2S24S126N001P023P003nsss(0) <='1';
          else
          cVar2S24S126N001P023P003nsss(0) <='0';
          end if;
        if(cVar1S25S126P018N061N042P050(0)='1' AND  A(29)='0' AND E(21)='1' )then
          cVar2S25S126P000P049nsss(0) <='1';
          else
          cVar2S25S126P000P049nsss(0) <='0';
          end if;
        if(cVar1S0S127P017P015P014P010(0)='1' AND  B(20)='1' )then
          cVar2S0S127P036nsss(0) <='1';
          else
          cVar2S0S127P036nsss(0) <='0';
          end if;
        if(cVar1S1S127P017P015P014P010(0)='1' AND  B(20)='0' AND B(24)='1' )then
          cVar2S1S127N036P028nsss(0) <='1';
          else
          cVar2S1S127N036P028nsss(0) <='0';
          end if;
        if(cVar1S2S127P017P015P014P010(0)='1' AND  B(20)='0' AND B(24)='0' AND B(11)='0' )then
          cVar2S2S127N036N028P035nsss(0) <='1';
          else
          cVar2S2S127N036N028P035nsss(0) <='0';
          end if;
        if(cVar1S3S127P017P015P014N010(0)='1' AND  B(22)='1' AND A(10)='0' )then
          cVar2S3S127P032P019nsss(0) <='1';
          else
          cVar2S3S127P032P019nsss(0) <='0';
          end if;
        if(cVar1S4S127P017P015P014N010(0)='1' AND  B(22)='1' AND A(10)='1' AND A(21)='1' )then
          cVar2S4S127P032P019P016nsss(0) <='1';
          else
          cVar2S4S127P032P019P016nsss(0) <='0';
          end if;
        if(cVar1S5S127P017P015P014N010(0)='1' AND  B(22)='0' AND B(17)='0' )then
          cVar2S5S127N032P023nsss(0) <='1';
          else
          cVar2S5S127N032P023nsss(0) <='0';
          end if;
        if(cVar1S6S127P017P015P014P066(0)='1' AND  A(24)='0' AND B(22)='0' AND E(11)='0' )then
          cVar2S6S127P010P032P056nsss(0) <='1';
          else
          cVar2S6S127P010P032P056nsss(0) <='0';
          end if;
        if(cVar1S7S127P017P015P014P066(0)='1' AND  A(24)='0' AND B(22)='1' AND D(18)='1' )then
          cVar2S7S127P010P032P059nsss(0) <='1';
          else
          cVar2S7S127P010P032P059nsss(0) <='0';
          end if;
        if(cVar1S8S127P017P015P014P066(0)='1' AND  A(24)='1' AND A(26)='0' AND A(10)='0' )then
          cVar2S8S127P010P006P019nsss(0) <='1';
          else
          cVar2S8S127P010P006P019nsss(0) <='0';
          end if;
        if(cVar1S9S127P017P015P014P066(0)='1' AND  E( 8)='1' AND A(13)='1' AND A(20)='1' )then
          cVar2S9S127P068P013P018nsss(0) <='1';
          else
          cVar2S9S127P068P013P018nsss(0) <='0';
          end if;
        if(cVar1S10S127P017P015P014P066(0)='1' AND  E( 8)='1' AND A(13)='0' AND A(23)='1' )then
          cVar2S10S127P068N013P012nsss(0) <='1';
          else
          cVar2S10S127P068N013P012nsss(0) <='0';
          end if;
        if(cVar1S11S127P017P015P000P019(0)='1' AND  B(24)='0' AND A(21)='0' )then
          cVar2S11S127P028P016nsss(0) <='1';
          else
          cVar2S11S127P028P016nsss(0) <='0';
          end if;
        if(cVar1S12S127P017P015P000P019(0)='1' AND  B(24)='0' AND A(21)='1' AND E(15)='1' )then
          cVar2S12S127P028P016P040nsss(0) <='1';
          else
          cVar2S12S127P028P016P040nsss(0) <='0';
          end if;
        if(cVar1S13S127P017P015P000N019(0)='1' AND  E(18)='0' AND B(28)='1' )then
          cVar2S13S127P061P020nsss(0) <='1';
          else
          cVar2S13S127P061P020nsss(0) <='0';
          end if;
        if(cVar1S14S127P017P015P000N019(0)='1' AND  E(18)='1' AND A(13)='0' AND A(21)='1' )then
          cVar2S14S127P061P013P016nsss(0) <='1';
          else
          cVar2S14S127P061P013P016nsss(0) <='0';
          end if;
        if(cVar1S15S127P017P015P000P008(0)='1' AND  D(17)='1' )then
          cVar2S15S127P063nsss(0) <='1';
          else
          cVar2S15S127P063nsss(0) <='0';
          end if;
        if(cVar1S16S127P017P015P000P008(0)='1' AND  D(17)='0' AND A(24)='0' AND A(21)='1' )then
          cVar2S16S127N063P010P016nsss(0) <='1';
          else
          cVar2S16S127N063P010P016nsss(0) <='0';
          end if;
        if(cVar1S18S127N017P018N027P002(0)='1' AND  A(27)='1' )then
          cVar2S18S127P004nsss(0) <='1';
          else
          cVar2S18S127P004nsss(0) <='0';
          end if;
        if(cVar1S19S127N017P018N027P002(0)='1' AND  A(27)='0' AND A(21)='0' AND A(22)='1' )then
          cVar2S19S127N004P016P014nsss(0) <='1';
          else
          cVar2S19S127N004P016P014nsss(0) <='0';
          end if;
        if(cVar1S20S127N017P018N027N002(0)='1' AND  D(12)='0' AND E(14)='1' )then
          cVar2S20S127P050P044nsss(0) <='1';
          else
          cVar2S20S127P050P044nsss(0) <='0';
          end if;
        if(cVar1S21S127N017P018N027N002(0)='1' AND  D(12)='0' AND E(14)='0' AND B(16)='0' )then
          cVar2S21S127P050N044P025nsss(0) <='1';
          else
          cVar2S21S127P050N044P025nsss(0) <='0';
          end if;
        if(cVar1S22S127N017P018N027N002(0)='1' AND  D(12)='1' AND B(14)='1' )then
          cVar2S22S127P050P029nsss(0) <='1';
          else
          cVar2S22S127P050P029nsss(0) <='0';
          end if;
        if(cVar1S23S127N017N018P067P045(0)='1' AND  B(20)='0' AND B(11)='0' AND D(23)='0' )then
          cVar2S23S127P036P035P039nsss(0) <='1';
          else
          cVar2S23S127P036P035P039nsss(0) <='0';
          end if;
        if(cVar1S24S127N017N018P067P045(0)='1' AND  B(20)='0' AND B(11)='1' AND A(22)='1' )then
          cVar2S24S127P036P035P014nsss(0) <='1';
          else
          cVar2S24S127P036P035P014nsss(0) <='0';
          end if;
        if(cVar1S25S127N017N018P067P045(0)='1' AND  B(20)='1' AND A(21)='1' AND A(14)='0' )then
          cVar2S25S127P036P016P011nsss(0) <='1';
          else
          cVar2S25S127P036P016P011nsss(0) <='0';
          end if;
        if(cVar1S26S127N017N018N067P009(0)='1' AND  A(14)='1' AND D(19)='1' )then
          cVar2S26S127P011P055nsss(0) <='1';
          else
          cVar2S26S127P011P055nsss(0) <='0';
          end if;
        if(cVar1S27S127N017N018N067P009(0)='1' AND  A(14)='1' AND D(19)='0' AND A(29)='0' )then
          cVar2S27S127P011N055P000nsss(0) <='1';
          else
          cVar2S27S127P011N055P000nsss(0) <='0';
          end if;
        if(cVar1S28S127N017N018N067P009(0)='1' AND  A(14)='0' AND B(20)='1' AND B(25)='0' )then
          cVar2S28S127N011P036P026nsss(0) <='1';
          else
          cVar2S28S127N011P036P026nsss(0) <='0';
          end if;
        if(cVar1S29S127N017N018N067P009(0)='1' AND  B(15)='1' )then
          cVar2S29S127P027nsss(0) <='1';
          else
          cVar2S29S127P027nsss(0) <='0';
          end if;
        if(cVar1S30S127N017N018N067P009(0)='1' AND  B(15)='0' AND A(16)='1' AND A(14)='0' )then
          cVar2S30S127N027P007P011nsss(0) <='1';
          else
          cVar2S30S127N027P007P011nsss(0) <='0';
          end if;
        if(cVar1S31S127N017N018N067P009(0)='1' AND  B(15)='0' AND A(16)='0' AND E(17)='1' )then
          cVar2S31S127N027N007P065nsss(0) <='1';
          else
          cVar2S31S127N027N007P065nsss(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV3 : process(c1)
begin
 if c1'event and c1='1' then
        if(cVar2S0S0P014P067nsss(0)='1'  OR cVar2S1S0P014P013P015nsss(0)='1'  OR cVar2S2S0P063P008nsss(0)='1'  OR cVar2S3S0P030nsss(0)='1'  )then
          oVar1S0(0) <='1';
          else
          oVar1S0(0) <='0';
          end if;
        if(cVar2S4S0N030P057P018nsss(0)='1'  OR cVar2S5S0P061P032nsss(0)='1'  OR cVar2S6S0P012nsss(0)='1'  OR cVar2S7S0P067P014P017nsss(0)='1'  )then
          oVar1S1(0) <='1';
          else
          oVar1S1(0) <='0';
          end if;
        if(cVar2S8S0N067P061nsss(0)='1'  OR cVar2S9S0N067N061P051nsss(0)='1'  OR cVar2S10S0P037P059nsss(0)='1'  OR cVar2S11S0N037P034P016nsss(0)='1'  )then
          oVar1S2(0) <='1';
          else
          oVar1S2(0) <='0';
          end if;
        if(cVar2S12S0P069P056P031nsss(0)='1'  OR cVar2S13S0P060P033nsss(0)='1'  OR cVar2S14S0P032P061nsss(0)='1'  OR cVar2S15S0N032P033P060nsss(0)='1'  )then
          oVar1S3(0) <='1';
          else
          oVar1S3(0) <='0';
          end if;
        if(cVar2S16S0P065P063P060nsss(0)='1'  OR cVar2S17S0N065P056P031nsss(0)='1'  )then
          oVar1S4(0) <='1';
          else
          oVar1S4(0) <='0';
          end if;
        if(cVar2S0S1P014nsss(0)='1'  OR cVar2S1S1P014P024P012nsss(0)='1'  OR cVar2S2S1P014P017P036nsss(0)='1'  OR cVar2S3S1P014P017P008nsss(0)='1'  )then
          oVar1S5(0) <='1';
          else
          oVar1S5(0) <='0';
          end if;
        if(cVar2S4S1P009nsss(0)='1'  OR cVar2S5S1P008P016nsss(0)='1'  OR cVar2S6S1N008P069nsss(0)='1'  OR cVar1S7S1P067P010P024P028nsss(0)='1'  )then
          oVar1S6(0) <='1';
          else
          oVar1S6(0) <='0';
          end if;
        if(cVar2S8S1P002P000P011nsss(0)='1'  OR cVar2S9S1P032nsss(0)='1'  OR cVar2S10S1P069nsss(0)='1'  OR cVar2S11S1N069P012nsss(0)='1'  )then
          oVar1S7(0) <='1';
          else
          oVar1S7(0) <='0';
          end if;
        if(cVar2S12S1N069N012P065nsss(0)='1'  OR cVar2S13S1P060nsss(0)='1'  OR cVar2S14S1N060P037nsss(0)='1'  OR cVar2S15S1N060N037P015nsss(0)='1'  )then
          oVar1S8(0) <='1';
          else
          oVar1S8(0) <='0';
          end if;
        if(cVar2S16S1P036P017P012nsss(0)='1'  OR cVar1S17S1N067N068P055P030nsss(0)='1'  OR cVar2S18S1P028nsss(0)='1'  OR cVar2S19S1N028P031nsss(0)='1'  )then
          oVar1S9(0) <='1';
          else
          oVar1S9(0) <='0';
          end if;
        if(cVar2S20S1N028N031P029nsss(0)='1'  OR cVar2S21S1P029nsss(0)='1'  OR cVar2S22S1N029P027nsss(0)='1'  OR cVar2S23S1N029N027P026nsss(0)='1'  )then
          oVar1S10(0) <='1';
          else
          oVar1S10(0) <='0';
          end if;
        if(cVar2S24S1P042nsss(0)='1'  OR cVar2S25S1N042P064nsss(0)='1'  OR cVar2S26S1N042N064P065nsss(0)='1'  )then
          oVar1S11(0) <='1';
          else
          oVar1S11(0) <='0';
          end if;
        if(cVar1S0S2P016P047P000P049nsss(0)='1'  OR cVar2S1S2P036P045nsss(0)='1'  OR cVar2S2S2P036N045P015nsss(0)='1'  OR cVar1S3S2P016N047P052P029nsss(0)='1'  )then
          oVar1S12(0) <='1';
          else
          oVar1S12(0) <='0';
          end if;
        if(cVar2S4S2P060nsss(0)='1'  OR cVar2S5S2P065P033P058nsss(0)='1'  OR cVar2S6S2P065N033psss(0)='1'  OR cVar2S7S2P065P064nsss(0)='1'  )then
          oVar1S13(0) <='1';
          else
          oVar1S13(0) <='0';
          end if;
        if(cVar2S8S2P046nsss(0)='1'  OR cVar2S9S2N046P040nsss(0)='1'  OR cVar2S10S2N046N040P015nsss(0)='1'  OR cVar2S11S2P034P008nsss(0)='1'  )then
          oVar1S14(0) <='1';
          else
          oVar1S14(0) <='0';
          end if;
        if(cVar2S12S2N034P036nsss(0)='1'  OR cVar2S13S2P019P067nsss(0)='1'  OR cVar2S14S2P019N067P062nsss(0)='1'  OR cVar2S15S2P019P015P066nsss(0)='1'  )then
          oVar1S15(0) <='1';
          else
          oVar1S15(0) <='0';
          end if;
        if(cVar2S16S2P011P058nsss(0)='1'  OR cVar2S17S2P011N058P062nsss(0)='1'  OR cVar2S18S2P065P062P012nsss(0)='1'  OR cVar2S19S2P065N062P027nsss(0)='1'  )then
          oVar1S16(0) <='1';
          else
          oVar1S16(0) <='0';
          end if;
        if(cVar2S20S2P067P062nsss(0)='1'  OR cVar2S21S2N067P060P012nsss(0)='1'  OR cVar2S22S2N067N060P029nsss(0)='1'  OR cVar2S23S2P044P028nsss(0)='1'  )then
          oVar1S17(0) <='1';
          else
          oVar1S17(0) <='0';
          end if;
        if(cVar2S24S2P026nsss(0)='1'  )then
          oVar1S18(0) <='1';
          else
          oVar1S18(0) <='0';
          end if;
        if(cVar1S0S3P047P049P064P014nsss(0)='1'  OR cVar2S1S3P012nsss(0)='1'  OR cVar1S2S3P047P049P064psss(0)='1'  OR cVar1S3S3P047N049P034P063nsss(0)='1'  )then
          oVar1S19(0) <='1';
          else
          oVar1S19(0) <='0';
          end if;
        if(cVar1S4S3N047P052P029nsss(0)='1'  OR cVar1S5S3N047P052N029P027nsss(0)='1'  OR cVar2S6S3P028nsss(0)='1'  OR cVar2S7S3N028P026P008nsss(0)='1'  )then
          oVar1S20(0) <='1';
          else
          oVar1S20(0) <='0';
          end if;
        if(cVar2S8S3N028N026P050nsss(0)='1'  OR cVar2S9S3P033P010nsss(0)='1'  OR cVar2S10S3N033psss(0)='1'  OR cVar2S11S3P010P059nsss(0)='1'  )then
          oVar1S21(0) <='1';
          else
          oVar1S21(0) <='0';
          end if;
        if(cVar2S12S3P046P025nsss(0)='1'  OR cVar2S13S3P046N025P027nsss(0)='1'  OR cVar2S14S3N046P028nsss(0)='1'  OR cVar2S15S3N046N028P040nsss(0)='1'  )then
          oVar1S22(0) <='1';
          else
          oVar1S22(0) <='0';
          end if;
        if(cVar2S16S3P024P067P010nsss(0)='1'  OR cVar2S17S3P024N067P005nsss(0)='1'  OR cVar2S18S3P024P045nsss(0)='1'  )then
          oVar1S23(0) <='1';
          else
          oVar1S23(0) <='0';
          end if;
        if(cVar2S0S4P004nsss(0)='1'  OR cVar2S1S4P004P018nsss(0)='1'  OR cVar2S2S4P062P052nsss(0)='1'  OR cVar2S3S4P062N052P016nsss(0)='1'  )then
          oVar1S24(0) <='1';
          else
          oVar1S24(0) <='0';
          end if;
        if(cVar2S4S4P066P012nsss(0)='1'  OR cVar2S5S4P028nsss(0)='1'  OR cVar2S6S4N028P064nsss(0)='1'  OR cVar2S7S4P059P068nsss(0)='1'  )then
          oVar1S25(0) <='1';
          else
          oVar1S25(0) <='0';
          end if;
        if(cVar2S8S4P043nsss(0)='1'  OR cVar2S9S4N043P024nsss(0)='1'  OR cVar2S10S4N043N024P068nsss(0)='1'  OR cVar2S11S4P027nsss(0)='1'  )then
          oVar1S26(0) <='1';
          else
          oVar1S26(0) <='0';
          end if;
        if(cVar2S12S4N027P056P004nsss(0)='1'  OR cVar2S13S4N027N056psss(0)='1'  OR cVar2S14S4P018P009nsss(0)='1'  OR cVar2S15S4P018P012nsss(0)='1'  )then
          oVar1S27(0) <='1';
          else
          oVar1S27(0) <='0';
          end if;
        if(cVar2S16S4P015nsss(0)='1'  OR cVar2S17S4P053nsss(0)='1'  OR cVar2S18S4N053P035nsss(0)='1'  OR cVar2S19S4N053N035P017nsss(0)='1'  )then
          oVar1S28(0) <='1';
          else
          oVar1S28(0) <='0';
          end if;
        if(cVar2S20S4P010P035P006nsss(0)='1'  OR cVar2S21S4P010N035P025nsss(0)='1'  OR cVar2S22S4P010P036P003nsss(0)='1'  OR cVar1S23S4P014P024P047nsss(0)='1'  )then
          oVar1S29(0) <='1';
          else
          oVar1S29(0) <='0';
          end if;
        if(cVar1S24S4P014P024N047P045nsss(0)='1'  )then
          oVar1S30(0) <='1';
          else
          oVar1S30(0) <='0';
          end if;
        if(cVar1S0S5P053P051P024P028nsss(0)='1'  OR cVar2S1S5P029nsss(0)='1'  OR cVar2S2S5N029P026nsss(0)='1'  OR cVar2S3S5N029N026P027nsss(0)='1'  )then
          oVar1S31(0) <='1';
          else
          oVar1S31(0) <='0';
          end if;
        if(cVar1S4S5P053N051P010P047nsss(0)='1'  OR cVar2S5S5P052nsss(0)='1'  OR cVar2S6S5N052P015P011nsss(0)='1'  OR cVar2S7S5N052N015P068nsss(0)='1'  )then
          oVar1S32(0) <='1';
          else
          oVar1S32(0) <='0';
          end if;
        if(cVar1S8S5P053N051P010P055nsss(0)='1'  OR cVar2S9S5P004P055P065nsss(0)='1'  OR cVar2S10S5P004N055psss(0)='1'  OR cVar2S11S5P004P066P067nsss(0)='1'  )then
          oVar1S33(0) <='1';
          else
          oVar1S33(0) <='0';
          end if;
        if(cVar2S12S5P057nsss(0)='1'  OR cVar2S13S5N057P052nsss(0)='1'  OR cVar2S14S5P043nsss(0)='1'  OR cVar2S15S5N043P047P016nsss(0)='1'  )then
          oVar1S34(0) <='1';
          else
          oVar1S34(0) <='0';
          end if;
        if(cVar2S16S5P048nsss(0)='1'  OR cVar2S17S5N048P056P054nsss(0)='1'  OR cVar2S18S5N048N056P038nsss(0)='1'  OR cVar2S19S5P062P017nsss(0)='1'  )then
          oVar1S35(0) <='1';
          else
          oVar1S35(0) <='0';
          end if;
        if(cVar2S20S5P069P045nsss(0)='1'  )then
          oVar1S36(0) <='1';
          else
          oVar1S36(0) <='0';
          end if;
        if(cVar1S0S6P047P049P064P012nsss(0)='1'  OR cVar2S1S6P016nsss(0)='1'  OR cVar2S2S6P009nsss(0)='1'  OR cVar2S3S6N009P068nsss(0)='1'  )then
          oVar1S37(0) <='1';
          else
          oVar1S37(0) <='0';
          end if;
        if(cVar2S4S6P057nsss(0)='1'  OR cVar2S5S6P026P031nsss(0)='1'  OR cVar2S6S6P026N031P004nsss(0)='1'  OR cVar2S7S6P051nsss(0)='1'  )then
          oVar1S38(0) <='1';
          else
          oVar1S38(0) <='0';
          end if;
        if(cVar2S8S6N051P010P052nsss(0)='1'  OR cVar2S9S6P051nsss(0)='1'  OR cVar2S10S6P043nsss(0)='1'  OR cVar2S11S6P012P015P014nsss(0)='1'  )then
          oVar1S39(0) <='1';
          else
          oVar1S39(0) <='0';
          end if;
        if(cVar2S12S6P012N015P046nsss(0)='1'  )then
          oVar1S40(0) <='1';
          else
          oVar1S40(0) <='0';
          end if;
        if(cVar1S0S7P053P006P028nsss(0)='1'  OR cVar1S1S7P053P006N028P029nsss(0)='1'  OR cVar2S2S7P026P008nsss(0)='1'  OR cVar2S3S7P026N008P019nsss(0)='1'  )then
          oVar1S41(0) <='1';
          else
          oVar1S41(0) <='0';
          end if;
        if(cVar2S4S7N026P027nsss(0)='1'  OR cVar2S5S7P019nsss(0)='1'  OR cVar2S6S7P068nsss(0)='1'  OR cVar2S7S7P068P017P037nsss(0)='1'  )then
          oVar1S42(0) <='1';
          else
          oVar1S42(0) <='0';
          end if;
        if(cVar2S8S7P002P057nsss(0)='1'  OR cVar2S9S7P002N057P013nsss(0)='1'  OR cVar2S10S7P018P057nsss(0)='1'  OR cVar1S11S7N053N055P047P049nsss(0)='1'  )then
          oVar1S43(0) <='1';
          else
          oVar1S43(0) <='0';
          end if;
        if(cVar2S12S7P024nsss(0)='1'  OR cVar2S13S7N024P019P017nsss(0)='1'  OR cVar2S14S7P058P059nsss(0)='1'  OR cVar2S15S7P058P059P015nsss(0)='1'  )then
          oVar1S44(0) <='1';
          else
          oVar1S44(0) <='0';
          end if;
        if(cVar2S16S7N058P061P032nsss(0)='1'  OR cVar2S17S7P023P042nsss(0)='1'  OR cVar2S18S7P023N042P045nsss(0)='1'  OR cVar2S19S7N023P022nsss(0)='1'  )then
          oVar1S45(0) <='1';
          else
          oVar1S45(0) <='0';
          end if;
        if(cVar1S0S8P036P053P000P028nsss(0)='1'  OR cVar2S1S8P026nsss(0)='1'  OR cVar2S2S8N026P029nsss(0)='1'  OR cVar2S3S8N026N029P041nsss(0)='1'  )then
          oVar1S47(0) <='1';
          else
          oVar1S47(0) <='0';
          end if;
        if(cVar1S4S8P036N053P046P025nsss(0)='1'  OR cVar2S5S8P027nsss(0)='1'  OR cVar2S6S8N027P024nsss(0)='1'  OR cVar2S7S8N027N024P015nsss(0)='1'  )then
          oVar1S48(0) <='1';
          else
          oVar1S48(0) <='0';
          end if;
        if(cVar2S8S8P015nsss(0)='1'  OR cVar2S9S8N015P041P039nsss(0)='1'  OR cVar2S10S8N015N041psss(0)='1'  OR cVar2S11S8P069P015P007nsss(0)='1'  )then
          oVar1S49(0) <='1';
          else
          oVar1S49(0) <='0';
          end if;
        if(cVar2S12S8P069P015P049nsss(0)='1'  OR cVar2S13S8P024P018P000nsss(0)='1'  OR cVar2S14S8P024P018P017nsss(0)='1'  OR cVar2S15S8P029nsss(0)='1'  )then
          oVar1S50(0) <='1';
          else
          oVar1S50(0) <='0';
          end if;
        if(cVar2S16S8N029P062P065nsss(0)='1'  OR cVar2S17S8N029N062psss(0)='1'  OR cVar2S18S8P017P066P035nsss(0)='1'  OR cVar2S19S8N017P019P012nsss(0)='1'  )then
          oVar1S51(0) <='1';
          else
          oVar1S51(0) <='0';
          end if;
        if(cVar2S20S8P018P014nsss(0)='1'  )then
          oVar1S52(0) <='1';
          else
          oVar1S52(0) <='0';
          end if;
        if(cVar1S0S9P052P029nsss(0)='1'  OR cVar1S1S9P052N029P027nsss(0)='1'  OR cVar1S2S9P052N029N027P028nsss(0)='1'  OR cVar2S3S9P026P008nsss(0)='1'  )then
          oVar1S53(0) <='1';
          else
          oVar1S53(0) <='0';
          end if;
        if(cVar2S4S9N026P062P035nsss(0)='1'  OR cVar1S5S9N052P046P025nsss(0)='1'  OR cVar2S6S9P027nsss(0)='1'  OR cVar2S7S9N027P024nsss(0)='1'  )then
          oVar1S54(0) <='1';
          else
          oVar1S54(0) <='0';
          end if;
        if(cVar2S8S9N027N024P033nsss(0)='1'  OR cVar2S9S9P020nsss(0)='1'  OR cVar2S10S9N020P021nsss(0)='1'  OR cVar2S11S9N020N021P012nsss(0)='1'  )then
          oVar1S55(0) <='1';
          else
          oVar1S55(0) <='0';
          end if;
        if(cVar2S12S9P065P043nsss(0)='1'  OR cVar2S13S9P053P028P012nsss(0)='1'  OR cVar2S14S9P053N028P026nsss(0)='1'  OR cVar2S15S9N053P015P051nsss(0)='1'  )then
          oVar1S56(0) <='1';
          else
          oVar1S56(0) <='0';
          end if;
        if(cVar2S16S9N053N015P023nsss(0)='1'  OR cVar2S17S9P012P069P014nsss(0)='1'  )then
          oVar1S57(0) <='1';
          else
          oVar1S57(0) <='0';
          end if;
        if(cVar1S0S10P012P053P063P028nsss(0)='1'  OR cVar2S1S10P029nsss(0)='1'  OR cVar2S2S10N029P026nsss(0)='1'  OR cVar2S3S10N029N026P065nsss(0)='1'  )then
          oVar1S58(0) <='1';
          else
          oVar1S58(0) <='0';
          end if;
        if(cVar2S4S10P014P051nsss(0)='1'  OR cVar2S5S10P020nsss(0)='1'  OR cVar2S6S10N020P021nsss(0)='1'  OR cVar2S7S10N020N021P018nsss(0)='1'  )then
          oVar1S59(0) <='1';
          else
          oVar1S59(0) <='0';
          end if;
        if(cVar2S8S10P069P016P043nsss(0)='1'  OR cVar2S9S10P046nsss(0)='1'  OR cVar2S10S10N046P002P020nsss(0)='1'  OR cVar2S11S10N046P002P040nsss(0)='1'  )then
          oVar1S60(0) <='1';
          else
          oVar1S60(0) <='0';
          end if;
        if(cVar2S12S10P050P008P034nsss(0)='1'  OR cVar2S13S10P056nsss(0)='1'  OR cVar2S14S10N056P057nsss(0)='1'  OR cVar2S15S10N056N057P013nsss(0)='1'  )then
          oVar1S61(0) <='1';
          else
          oVar1S61(0) <='0';
          end if;
        if(cVar2S16S10P017P015nsss(0)='1'  OR cVar2S17S10P063nsss(0)='1'  OR cVar2S18S10N063P066nsss(0)='1'  OR cVar2S19S10N063N066P015nsss(0)='1'  )then
          oVar1S62(0) <='1';
          else
          oVar1S62(0) <='0';
          end if;
        if(cVar2S20S10P014P015P025nsss(0)='1'  OR cVar2S21S10P014P015P032nsss(0)='1'  OR cVar2S22S10N014P066P019nsss(0)='1'  OR cVar2S23S10P057P026nsss(0)='1'  )then
          oVar1S63(0) <='1';
          else
          oVar1S63(0) <='0';
          end if;
        if(cVar1S0S11P053P006P028nsss(0)='1'  OR cVar1S1S11P053P006N028P029nsss(0)='1'  OR cVar2S2S11P026P008nsss(0)='1'  OR cVar2S3S11P026N008P019nsss(0)='1'  )then
          oVar1S65(0) <='1';
          else
          oVar1S65(0) <='0';
          end if;
        if(cVar2S4S11N026P009P010nsss(0)='1'  OR cVar2S5S11P019nsss(0)='1'  OR cVar1S6S11N053P041P020nsss(0)='1'  OR cVar1S7S11N053P041N020P021nsss(0)='1'  )then
          oVar1S66(0) <='1';
          else
          oVar1S66(0) <='0';
          end if;
        if(cVar2S8S11P008P065P069nsss(0)='1'  OR cVar2S9S11P025nsss(0)='1'  OR cVar2S10S11N025P027nsss(0)='1'  OR cVar2S11S11N025N027P024nsss(0)='1'  )then
          oVar1S67(0) <='1';
          else
          oVar1S67(0) <='0';
          end if;
        if(cVar2S12S11P030P057nsss(0)='1'  OR cVar2S13S11P030N057P054nsss(0)='1'  OR cVar2S14S11N030P052P050nsss(0)='1'  OR cVar2S15S11N030N052P045nsss(0)='1'  )then
          oVar1S68(0) <='1';
          else
          oVar1S68(0) <='0';
          end if;
        if(cVar2S16S11P007P012P009nsss(0)='1'  )then
          oVar1S69(0) <='1';
          else
          oVar1S69(0) <='0';
          end if;
        if(cVar2S0S12P024P068nsss(0)='1'  OR cVar2S1S12P024N068P008nsss(0)='1'  OR cVar2S2S12P018nsss(0)='1'  OR cVar2S3S12P034nsss(0)='1'  )then
          oVar1S70(0) <='1';
          else
          oVar1S70(0) <='0';
          end if;
        if(cVar2S4S12N034P036P014nsss(0)='1'  OR cVar2S5S12P065P034nsss(0)='1'  OR cVar2S6S12P065P067P069nsss(0)='1'  OR cVar2S7S12P020nsss(0)='1'  )then
          oVar1S71(0) <='1';
          else
          oVar1S71(0) <='0';
          end if;
        if(cVar2S8S12N020P012nsss(0)='1'  OR cVar2S9S12P027nsss(0)='1'  OR cVar2S10S12N027P034nsss(0)='1'  OR cVar2S11S12N027P034P061nsss(0)='1'  )then
          oVar1S72(0) <='1';
          else
          oVar1S72(0) <='0';
          end if;
        if(cVar2S12S12P034P014P062nsss(0)='1'  OR cVar2S13S12P034N014P017nsss(0)='1'  OR cVar2S14S12N034P017P011nsss(0)='1'  OR cVar2S15S12P061nsss(0)='1'  )then
          oVar1S73(0) <='1';
          else
          oVar1S73(0) <='0';
          end if;
        if(cVar2S16S12N061P007nsss(0)='1'  OR cVar2S17S12P051P011nsss(0)='1'  OR cVar2S18S12P051P011P013nsss(0)='1'  OR cVar2S19S12P060P053nsss(0)='1'  )then
          oVar1S74(0) <='1';
          else
          oVar1S74(0) <='0';
          end if;
        if(cVar2S20S12P060N053P014nsss(0)='1'  OR cVar2S21S12P058nsss(0)='1'  OR cVar2S22S12N058P057nsss(0)='1'  OR cVar2S23S12P017P058P054nsss(0)='1'  )then
          oVar1S75(0) <='1';
          else
          oVar1S75(0) <='0';
          end if;
        if(cVar2S0S13P064P062nsss(0)='1'  OR cVar2S1S13P064N062P014nsss(0)='1'  OR cVar2S2S13N064P003P017nsss(0)='1'  OR cVar2S3S13P008P060P062nsss(0)='1'  )then
          oVar1S77(0) <='1';
          else
          oVar1S77(0) <='0';
          end if;
        if(cVar2S4S13P018P067P008nsss(0)='1'  OR cVar2S5S13P018N067P068nsss(0)='1'  OR cVar2S6S13N018P019P059nsss(0)='1'  OR cVar2S7S13P050nsss(0)='1'  )then
          oVar1S78(0) <='1';
          else
          oVar1S78(0) <='0';
          end if;
        if(cVar2S8S13N050P019nsss(0)='1'  OR cVar2S9S13P048nsss(0)='1'  OR cVar2S10S13N048P054P050nsss(0)='1'  OR cVar2S11S13P029nsss(0)='1'  )then
          oVar1S79(0) <='1';
          else
          oVar1S79(0) <='0';
          end if;
        if(cVar2S12S13N029P028nsss(0)='1'  OR cVar2S13S13N029N028P026nsss(0)='1'  OR cVar2S14S13P055P030nsss(0)='1'  OR cVar2S15S13P055N030P032nsss(0)='1'  )then
          oVar1S80(0) <='1';
          else
          oVar1S80(0) <='0';
          end if;
        if(cVar2S16S13N055P041P039nsss(0)='1'  OR cVar2S17S13N055N041P015nsss(0)='1'  OR cVar2S18S13P018P009P019nsss(0)='1'  OR cVar2S19S13N018P003P012nsss(0)='1'  )then
          oVar1S81(0) <='1';
          else
          oVar1S81(0) <='0';
          end if;
        if(cVar1S0S14P015P016P034P063nsss(0)='1'  OR cVar2S1S14P011P065nsss(0)='1'  OR cVar2S2S14P050P018nsss(0)='1'  OR cVar2S3S14P050P018P035nsss(0)='1'  )then
          oVar1S83(0) <='1';
          else
          oVar1S83(0) <='0';
          end if;
        if(cVar2S4S14P003P066nsss(0)='1'  OR cVar2S5S14N003P009P024nsss(0)='1'  OR cVar2S6S14N003N009P059nsss(0)='1'  OR cVar1S7S14P015N016P046P025nsss(0)='1'  )then
          oVar1S84(0) <='1';
          else
          oVar1S84(0) <='0';
          end if;
        if(cVar2S8S14P003P009nsss(0)='1'  OR cVar2S9S14P003N009P024nsss(0)='1'  OR cVar2S10S14P043nsss(0)='1'  OR cVar2S11S14N043P042nsss(0)='1'  )then
          oVar1S85(0) <='1';
          else
          oVar1S85(0) <='0';
          end if;
        if(cVar2S12S14N043N042P017nsss(0)='1'  OR cVar2S13S14P056P029nsss(0)='1'  OR cVar2S14S14P056N029P012nsss(0)='1'  OR cVar2S15S14N056P047P049nsss(0)='1'  )then
          oVar1S86(0) <='1';
          else
          oVar1S86(0) <='0';
          end if;
        if(cVar2S16S14N056N047P065nsss(0)='1'  OR cVar2S17S14P061nsss(0)='1'  OR cVar2S18S14N061P036nsss(0)='1'  OR cVar2S19S14P050P035P034nsss(0)='1'  )then
          oVar1S87(0) <='1';
          else
          oVar1S87(0) <='0';
          end if;
        if(cVar2S20S14P050N035P060nsss(0)='1'  OR cVar2S21S14P033P061nsss(0)='1'  OR cVar2S22S14P033N061P060nsss(0)='1'  OR cVar2S23S14N033P035P018nsss(0)='1'  )then
          oVar1S88(0) <='1';
          else
          oVar1S88(0) <='0';
          end if;
        if(cVar2S24S14P068P062nsss(0)='1'  OR cVar2S25S14N068P017P000nsss(0)='1'  OR cVar1S26S14P015P009P027nsss(0)='1'  )then
          oVar1S89(0) <='1';
          else
          oVar1S89(0) <='0';
          end if;
        if(cVar1S0S15P046P025nsss(0)='1'  OR cVar2S1S15P047nsss(0)='1'  OR cVar2S2S15N047P016nsss(0)='1'  OR cVar2S3S15N047P016P012nsss(0)='1'  )then
          oVar1S90(0) <='1';
          else
          oVar1S90(0) <='0';
          end if;
        if(cVar2S4S15P035P013P015nsss(0)='1'  OR cVar2S5S15P000P063P008nsss(0)='1'  OR cVar2S6S15P000N063P011nsss(0)='1'  OR cVar2S7S15P035P051P062nsss(0)='1'  )then
          oVar1S91(0) <='1';
          else
          oVar1S91(0) <='0';
          end if;
        if(cVar2S8S15N035P036P024nsss(0)='1'  OR cVar2S9S15N035N036P065nsss(0)='1'  OR cVar2S10S15P022P008P041nsss(0)='1'  OR cVar2S11S15P022P008P037nsss(0)='1'  )then
          oVar1S92(0) <='1';
          else
          oVar1S92(0) <='0';
          end if;
        if(cVar2S12S15P057P068P034nsss(0)='1'  OR cVar1S13S15N046N016P056P057nsss(0)='1'  OR cVar2S14S15P029nsss(0)='1'  OR cVar2S15S15N029P012nsss(0)='1'  )then
          oVar1S93(0) <='1';
          else
          oVar1S93(0) <='0';
          end if;
        if(cVar2S16S15P047P049nsss(0)='1'  OR cVar2S17S15N047P041P020nsss(0)='1'  OR cVar2S18S15N047N041P038nsss(0)='1'  OR cVar2S19S15P029nsss(0)='1'  )then
          oVar1S94(0) <='1';
          else
          oVar1S94(0) <='0';
          end if;
        if(cVar1S0S16P016P000P023P042nsss(0)='1'  OR cVar2S1S16P045nsss(0)='1'  OR cVar2S2S16P043nsss(0)='1'  OR cVar2S3S16N043P014P042nsss(0)='1'  )then
          oVar1S96(0) <='1';
          else
          oVar1S96(0) <='0';
          end if;
        if(cVar2S4S16P042nsss(0)='1'  OR cVar2S5S16P042N040P069nsss(0)='1'  OR cVar2S6S16P060P056P002nsss(0)='1'  OR cVar2S7S16P011P018nsss(0)='1'  )then
          oVar1S97(0) <='1';
          else
          oVar1S97(0) <='0';
          end if;
        if(cVar2S8S16P011P018P017nsss(0)='1'  OR cVar2S9S16P011P017nsss(0)='1'  OR cVar2S10S16P000P065P068nsss(0)='1'  OR cVar2S11S16P050nsss(0)='1'  )then
          oVar1S98(0) <='1';
          else
          oVar1S98(0) <='0';
          end if;
        if(cVar2S12S16P003P066P013nsss(0)='1'  OR cVar2S13S16N003P009P066nsss(0)='1'  OR cVar2S14S16N003N009P036nsss(0)='1'  OR cVar2S15S16P045P035nsss(0)='1'  )then
          oVar1S99(0) <='1';
          else
          oVar1S99(0) <='0';
          end if;
        if(cVar2S16S16P045N035P061nsss(0)='1'  OR cVar2S17S16P024P057P068nsss(0)='1'  OR cVar2S18S16P036P012P017nsss(0)='1'  )then
          oVar1S100(0) <='1';
          else
          oVar1S100(0) <='0';
          end if;
        if(cVar1S0S17P023P042nsss(0)='1'  OR cVar1S1S17P023N042P005nsss(0)='1'  OR cVar2S2S17P062P022P066nsss(0)='1'  OR cVar2S3S17P024P028nsss(0)='1'  )then
          oVar1S101(0) <='1';
          else
          oVar1S101(0) <='0';
          end if;
        if(cVar2S4S17P024N028P039nsss(0)='1'  OR cVar2S5S17P062P017P012nsss(0)='1'  OR cVar2S6S17P011P033P019nsss(0)='1'  OR cVar2S7S17P011N033P032nsss(0)='1'  )then
          oVar1S102(0) <='1';
          else
          oVar1S102(0) <='0';
          end if;
        if(cVar2S8S17P011P013P015nsss(0)='1'  OR cVar2S9S17P022P004nsss(0)='1'  OR cVar2S10S17P022N004P035nsss(0)='1'  OR cVar2S11S17N022P043P034nsss(0)='1'  )then
          oVar1S103(0) <='1';
          else
          oVar1S103(0) <='0';
          end if;
        if(cVar2S12S17N022P043P024nsss(0)='1'  OR cVar1S13S17N023P005P006P041nsss(0)='1'  OR cVar2S14S17P047nsss(0)='1'  OR cVar2S15S17N047P043nsss(0)='1'  )then
          oVar1S104(0) <='1';
          else
          oVar1S104(0) <='0';
          end if;
        if(cVar2S0S18P032nsss(0)='1'  OR cVar2S1S18N032P033nsss(0)='1'  OR cVar2S2S18N032N033P035nsss(0)='1'  OR cVar2S3S18P016nsss(0)='1'  )then
          oVar1S106(0) <='1';
          else
          oVar1S106(0) <='0';
          end if;
        if(cVar1S4S18P011N058P046P025nsss(0)='1'  OR cVar2S5S18P047nsss(0)='1'  OR cVar2S6S18N047P014nsss(0)='1'  OR cVar2S7S18P040nsss(0)='1'  )then
          oVar1S107(0) <='1';
          else
          oVar1S107(0) <='0';
          end if;
        if(cVar2S8S18N040P039nsss(0)='1'  OR cVar2S9S18P020P039nsss(0)='1'  OR cVar2S10S18P020N039P040nsss(0)='1'  OR cVar2S11S18N020P039P038nsss(0)='1'  )then
          oVar1S108(0) <='1';
          else
          oVar1S108(0) <='0';
          end if;
        if(cVar1S12S18P011P029P066P054nsss(0)='1'  OR cVar2S13S18P051nsss(0)='1'  OR cVar2S14S18N051P052nsss(0)='1'  OR cVar2S15S18N051N052P014nsss(0)='1'  )then
          oVar1S109(0) <='1';
          else
          oVar1S109(0) <='0';
          end if;
        if(cVar2S16S18P003P028nsss(0)='1'  OR cVar2S17S18P003N028P027nsss(0)='1'  OR cVar2S18S18P003P015P018nsss(0)='1'  OR cVar2S19S18P008P015P012nsss(0)='1'  )then
          oVar1S110(0) <='1';
          else
          oVar1S110(0) <='0';
          end if;
        if(cVar1S0S19P021P040nsss(0)='1'  OR cVar1S1S19P021N040P041nsss(0)='1'  OR cVar2S2S19P067P006nsss(0)='1'  OR cVar2S3S19P067N006P011nsss(0)='1'  )then
          oVar1S112(0) <='1';
          else
          oVar1S112(0) <='0';
          end if;
        if(cVar2S4S19P011P013nsss(0)='1'  OR cVar2S5S19P011N013P026nsss(0)='1'  OR cVar2S6S19P039nsss(0)='1'  OR cVar2S7S19N039P040nsss(0)='1'  )then
          oVar1S113(0) <='1';
          else
          oVar1S113(0) <='0';
          end if;
        if(cVar2S8S19N039N040P064nsss(0)='1'  OR cVar2S9S19P039P046nsss(0)='1'  OR cVar2S10S19P060P018P035nsss(0)='1'  )then
          oVar1S114(0) <='1';
          else
          oVar1S114(0) <='0';
          end if;
        if(cVar1S0S20P032P023P042nsss(0)='1'  OR cVar1S1S20P032P023N042P005nsss(0)='1'  OR cVar2S2S20P067P043nsss(0)='1'  OR cVar2S3S20P000P039nsss(0)='1'  )then
          oVar1S115(0) <='1';
          else
          oVar1S115(0) <='0';
          end if;
        if(cVar2S4S20P054P035P045nsss(0)='1'  OR cVar2S5S20P054N035psss(0)='1'  OR cVar2S6S20P054P052P010nsss(0)='1'  OR cVar2S7S20P006P039nsss(0)='1'  )then
          oVar1S116(0) <='1';
          else
          oVar1S116(0) <='0';
          end if;
        if(cVar2S8S20P006N039P043nsss(0)='1'  OR cVar2S9S20P060nsss(0)='1'  OR cVar2S10S20N060P034P063nsss(0)='1'  OR cVar2S11S20P064nsss(0)='1'  )then
          oVar1S117(0) <='1';
          else
          oVar1S117(0) <='0';
          end if;
        if(cVar2S12S20N064P036P066nsss(0)='1'  OR cVar2S13S20P059P069P016nsss(0)='1'  OR cVar2S14S20P059P015nsss(0)='1'  OR cVar2S15S20P017nsss(0)='1'  )then
          oVar1S118(0) <='1';
          else
          oVar1S118(0) <='0';
          end if;
        if(cVar1S0S21P023P042nsss(0)='1'  OR cVar1S1S21P023N042P024P005nsss(0)='1'  OR cVar2S2S21P067P015P068nsss(0)='1'  OR cVar2S3S21P010nsss(0)='1'  )then
          oVar1S120(0) <='1';
          else
          oVar1S120(0) <='0';
          end if;
        if(cVar2S4S21P026nsss(0)='1'  OR cVar2S5S21N026P025nsss(0)='1'  OR cVar2S6S21N026N025P027nsss(0)='1'  OR cVar2S7S21P056P039P004nsss(0)='1'  )then
          oVar1S121(0) <='1';
          else
          oVar1S121(0) <='0';
          end if;
        if(cVar2S8S21N056P052P029nsss(0)='1'  OR cVar2S9S21P032P043P015nsss(0)='1'  OR cVar2S10S21P051P018P009nsss(0)='1'  )then
          oVar1S122(0) <='1';
          else
          oVar1S122(0) <='0';
          end if;
        if(cVar2S0S22P050nsss(0)='1'  OR cVar2S1S22N050P009P014nsss(0)='1'  OR cVar2S2S22P050nsss(0)='1'  OR cVar2S3S22P050P029nsss(0)='1'  )then
          oVar1S123(0) <='1';
          else
          oVar1S123(0) <='0';
          end if;
        if(cVar2S4S22P050N029P026nsss(0)='1'  OR cVar2S5S22P011P066nsss(0)='1'  OR cVar2S6S22N011P008nsss(0)='1'  OR cVar1S7S22P001P010P028P034nsss(0)='1'  )then
          oVar1S124(0) <='1';
          else
          oVar1S124(0) <='0';
          end if;
        if(cVar2S8S22P024P029nsss(0)='1'  OR cVar2S9S22P024N029P058nsss(0)='1'  OR cVar2S10S22P034P012nsss(0)='1'  OR cVar2S11S22P016P035nsss(0)='1'  )then
          oVar1S125(0) <='1';
          else
          oVar1S125(0) <='0';
          end if;
        if(cVar2S12S22P016N035P019nsss(0)='1'  )then
          oVar1S126(0) <='1';
          else
          oVar1S126(0) <='0';
          end if;
        if(cVar1S0S23P027P000P048nsss(0)='1'  OR cVar2S1S23P062P009nsss(0)='1'  OR cVar2S2S23P062N009P014nsss(0)='1'  OR cVar1S3S23N027P009P023P042nsss(0)='1'  )then
          oVar1S127(0) <='1';
          else
          oVar1S127(0) <='0';
          end if;
        if(cVar2S4S23P045nsss(0)='1'  OR cVar2S5S23N045P069P036nsss(0)='1'  OR cVar2S6S23P062P051nsss(0)='1'  OR cVar2S7S23N062P063P065nsss(0)='1'  )then
          oVar1S128(0) <='1';
          else
          oVar1S128(0) <='0';
          end if;
        if(cVar2S8S23P022P043nsss(0)='1'  OR cVar2S9S23P022N043P014nsss(0)='1'  OR cVar2S10S23N022P043P021nsss(0)='1'  OR cVar2S11S23P066P036P019nsss(0)='1'  )then
          oVar1S129(0) <='1';
          else
          oVar1S129(0) <='0';
          end if;
        if(cVar2S12S23P066N036P047nsss(0)='1'  OR cVar2S13S23P014P064P019nsss(0)='1'  OR cVar2S14S23P066P059nsss(0)='1'  )then
          oVar1S130(0) <='1';
          else
          oVar1S130(0) <='0';
          end if;
        if(cVar2S0S24P030nsss(0)='1'  OR cVar2S1S24N030P031nsss(0)='1'  OR cVar2S2S24N030N031P068nsss(0)='1'  OR cVar2S3S24P013P016nsss(0)='1'  )then
          oVar1S131(0) <='1';
          else
          oVar1S131(0) <='0';
          end if;
        if(cVar2S4S24P013N016P014nsss(0)='1'  OR cVar2S5S24P020nsss(0)='1'  OR cVar2S6S24N020P021nsss(0)='1'  OR cVar2S7S24N020N021P004nsss(0)='1'  )then
          oVar1S132(0) <='1';
          else
          oVar1S132(0) <='0';
          end if;
        if(cVar2S8S24P039nsss(0)='1'  OR cVar1S9S24P008P026P045P047nsss(0)='1'  OR cVar2S10S24P055P004P010nsss(0)='1'  OR cVar1S11S24P008P026P004P051nsss(0)='1'  )then
          oVar1S133(0) <='1';
          else
          oVar1S133(0) <='0';
          end if;
        if(cVar2S12S24P050nsss(0)='1'  OR cVar2S13S24N050P062P067nsss(0)='1'  OR cVar2S14S24P068P065P063nsss(0)='1'  OR cVar2S15S24P068N065P067nsss(0)='1'  )then
          oVar1S134(0) <='1';
          else
          oVar1S134(0) <='0';
          end if;
        if(cVar2S16S24N068P036P028nsss(0)='1'  OR cVar2S17S24N068P036P033nsss(0)='1'  )then
          oVar1S135(0) <='1';
          else
          oVar1S135(0) <='0';
          end if;
        if(cVar2S0S25P014nsss(0)='1'  OR cVar2S1S25P014P019nsss(0)='1'  OR cVar2S2S25P013nsss(0)='1'  OR cVar2S3S25P004P010P069nsss(0)='1'  )then
          oVar1S136(0) <='1';
          else
          oVar1S136(0) <='0';
          end if;
        if(cVar2S4S25P004N010P032nsss(0)='1'  OR cVar1S5S25N055P057P041P020nsss(0)='1'  OR cVar2S6S25P021nsss(0)='1'  OR cVar2S7S25N021P008P035nsss(0)='1'  )then
          oVar1S137(0) <='1';
          else
          oVar1S137(0) <='0';
          end if;
        if(cVar2S8S25P028P012nsss(0)='1'  OR cVar2S9S25N028P029nsss(0)='1'  OR cVar2S10S25N028N029P069nsss(0)='1'  OR cVar2S11S25P040P021nsss(0)='1'  )then
          oVar1S138(0) <='1';
          else
          oVar1S138(0) <='0';
          end if;
        if(cVar2S12S25P040N021P020nsss(0)='1'  OR cVar2S13S25P061P069P059nsss(0)='1'  )then
          oVar1S139(0) <='1';
          else
          oVar1S139(0) <='0';
          end if;
        if(cVar2S0S26P062P064nsss(0)='1'  OR cVar2S1S26P062N064P066nsss(0)='1'  OR cVar2S2S26N062P067nsss(0)='1'  OR cVar2S3S26N062N067P064nsss(0)='1'  )then
          oVar1S140(0) <='1';
          else
          oVar1S140(0) <='0';
          end if;
        if(cVar2S4S26P066nsss(0)='1'  OR cVar2S5S26P067P015P011nsss(0)='1'  OR cVar2S6S26N067P026nsss(0)='1'  OR cVar2S7S26N067N026P036nsss(0)='1'  )then
          oVar1S141(0) <='1';
          else
          oVar1S141(0) <='0';
          end if;
        if(cVar2S8S26P024P020P034nsss(0)='1'  OR cVar2S9S26P024P008nsss(0)='1'  OR cVar1S10S26P017N019P037P064nsss(0)='1'  OR cVar2S11S26P035P015nsss(0)='1'  )then
          oVar1S142(0) <='1';
          else
          oVar1S142(0) <='0';
          end if;
        if(cVar2S12S26N035P066P013nsss(0)='1'  OR cVar2S13S26N035N066P058nsss(0)='1'  OR cVar2S14S26P018P015P066nsss(0)='1'  OR cVar2S15S26P018N015P013nsss(0)='1'  )then
          oVar1S143(0) <='1';
          else
          oVar1S143(0) <='0';
          end if;
        if(cVar2S16S26N018P016P015nsss(0)='1'  OR cVar2S17S26P018nsss(0)='1'  OR cVar2S18S26N018P015nsss(0)='1'  OR cVar2S19S26P006P003nsss(0)='1'  )then
          oVar1S144(0) <='1';
          else
          oVar1S144(0) <='0';
          end if;
        if(cVar2S20S26P009P055nsss(0)='1'  OR cVar2S21S26P009N055P066nsss(0)='1'  OR cVar2S22S26P009P036nsss(0)='1'  OR cVar2S23S26P062P035nsss(0)='1'  )then
          oVar1S145(0) <='1';
          else
          oVar1S145(0) <='0';
          end if;
        if(cVar2S24S26P062N035P015nsss(0)='1'  OR cVar2S25S26P015P066nsss(0)='1'  OR cVar2S26S26P015P066P068nsss(0)='1'  OR cVar2S27S26P015P016nsss(0)='1'  )then
          oVar1S146(0) <='1';
          else
          oVar1S146(0) <='0';
          end if;
        if(cVar2S28S26P051P002P054nsss(0)='1'  OR cVar2S29S26P003P068P008nsss(0)='1'  OR cVar2S30S26P011P018nsss(0)='1'  OR cVar2S31S26N011P069P068nsss(0)='1'  )then
          oVar1S147(0) <='1';
          else
          oVar1S147(0) <='0';
          end if;
        if(cVar2S0S27P045P022nsss(0)='1'  OR cVar1S1S27P017P051P048P026nsss(0)='1'  OR cVar2S2S27P019P018P015nsss(0)='1'  OR cVar2S3S27P019N018P053nsss(0)='1'  )then
          oVar1S149(0) <='1';
          else
          oVar1S149(0) <='0';
          end if;
        if(cVar2S4S27P019P014P037nsss(0)='1'  OR cVar2S5S27P000P007nsss(0)='1'  OR cVar2S6S27P000P007P012nsss(0)='1'  OR cVar2S7S27P062P015nsss(0)='1'  )then
          oVar1S150(0) <='1';
          else
          oVar1S150(0) <='0';
          end if;
        if(cVar2S8S27P062P015P066nsss(0)='1'  OR cVar2S9S27N062P007nsss(0)='1'  OR cVar2S10S27N062N007P064nsss(0)='1'  OR cVar2S11S27P008P032nsss(0)='1'  )then
          oVar1S151(0) <='1';
          else
          oVar1S151(0) <='0';
          end if;
        if(cVar2S12S27P048nsss(0)='1'  OR cVar2S13S27N048P009nsss(0)='1'  OR cVar2S14S27N048N009P026nsss(0)='1'  OR cVar2S15S27P029P011nsss(0)='1'  )then
          oVar1S152(0) <='1';
          else
          oVar1S152(0) <='0';
          end if;
        if(cVar2S16S27P029N011P009nsss(0)='1'  OR cVar2S17S27N029P023nsss(0)='1'  OR cVar2S18S27N029N023P025nsss(0)='1'  OR cVar2S19S27P055P065P003nsss(0)='1'  )then
          oVar1S153(0) <='1';
          else
          oVar1S153(0) <='0';
          end if;
        if(cVar2S20S27P067P020P057nsss(0)='1'  )then
          oVar1S154(0) <='1';
          else
          oVar1S154(0) <='0';
          end if;
        if(cVar2S0S28P023nsss(0)='1'  OR cVar2S1S28N023P022nsss(0)='1'  OR cVar2S2S28N023N022P007nsss(0)='1'  OR cVar2S3S28P042nsss(0)='1'  )then
          oVar1S155(0) <='1';
          else
          oVar1S155(0) <='0';
          end if;
        if(cVar2S4S28P042P040nsss(0)='1'  OR cVar1S5S28P017P068P064P055nsss(0)='1'  OR cVar2S6S28P067P065P014nsss(0)='1'  OR cVar2S7S28N067P062P058nsss(0)='1'  )then
          oVar1S156(0) <='1';
          else
          oVar1S156(0) <='0';
          end if;
        if(cVar2S8S28P009P034nsss(0)='1'  OR cVar2S9S28P009N034P013nsss(0)='1'  OR cVar2S10S28P035P002nsss(0)='1'  OR cVar2S11S28P063P037P012nsss(0)='1'  )then
          oVar1S157(0) <='1';
          else
          oVar1S157(0) <='0';
          end if;
        if(cVar2S12S28P063P037P016nsss(0)='1'  OR cVar2S13S28P063P015nsss(0)='1'  OR cVar2S14S28P044P012P004nsss(0)='1'  OR cVar2S15S28P044N012P065nsss(0)='1'  )then
          oVar1S158(0) <='1';
          else
          oVar1S158(0) <='0';
          end if;
        if(cVar2S16S28P065nsss(0)='1'  OR cVar2S17S28N065P037P018nsss(0)='1'  OR cVar2S18S28P000P009nsss(0)='1'  OR cVar2S19S28P013P063P064nsss(0)='1'  )then
          oVar1S159(0) <='1';
          else
          oVar1S159(0) <='0';
          end if;
        if(cVar2S20S28P013N063P062nsss(0)='1'  OR cVar2S21S28P013P065P014nsss(0)='1'  OR cVar2S22S28P014P051P069nsss(0)='1'  OR cVar2S23S28P014P018P015nsss(0)='1'  )then
          oVar1S160(0) <='1';
          else
          oVar1S160(0) <='0';
          end if;
        if(cVar2S24S28P065nsss(0)='1'  OR cVar2S25S28N065P069P012nsss(0)='1'  OR cVar2S26S28P011P036nsss(0)='1'  OR cVar2S27S28P011N036P016nsss(0)='1'  )then
          oVar1S161(0) <='1';
          else
          oVar1S161(0) <='0';
          end if;
        if(cVar2S0S29P034P020nsss(0)='1'  OR cVar2S1S29P034P015P019nsss(0)='1'  OR cVar2S2S29P063P034P060nsss(0)='1'  OR cVar2S3S29P063N034P030nsss(0)='1'  )then
          oVar1S163(0) <='1';
          else
          oVar1S163(0) <='0';
          end if;
        if(cVar2S4S29N063P065P031nsss(0)='1'  OR cVar2S5S29P010nsss(0)='1'  OR cVar2S6S29P020P016P024nsss(0)='1'  OR cVar2S7S29P018P069P012nsss(0)='1'  )then
          oVar1S164(0) <='1';
          else
          oVar1S164(0) <='0';
          end if;
        if(cVar1S8S29N017P044P023nsss(0)='1'  OR cVar1S9S29N017P044N023P025nsss(0)='1'  OR cVar2S10S29P007P022nsss(0)='1'  OR cVar2S11S29P030P068nsss(0)='1'  )then
          oVar1S165(0) <='1';
          else
          oVar1S165(0) <='0';
          end if;
        if(cVar2S12S29P030P068P037nsss(0)='1'  OR cVar2S13S29N030P031nsss(0)='1'  OR cVar2S14S29N030N031P032nsss(0)='1'  OR cVar2S15S29P065nsss(0)='1'  )then
          oVar1S166(0) <='1';
          else
          oVar1S166(0) <='0';
          end if;
        if(cVar2S16S29P020nsss(0)='1'  OR cVar2S17S29N020P061P021nsss(0)='1'  OR cVar2S18S29P036P047nsss(0)='1'  OR cVar2S19S29P036P016P002nsss(0)='1'  )then
          oVar1S167(0) <='1';
          else
          oVar1S167(0) <='0';
          end if;
        if(cVar2S0S30P023nsss(0)='1'  OR cVar2S1S30N023P022nsss(0)='1'  OR cVar2S2S30N023N022P062nsss(0)='1'  OR cVar2S3S30P020nsss(0)='1'  )then
          oVar1S169(0) <='1';
          else
          oVar1S169(0) <='0';
          end if;
        if(cVar2S4S30N020P059P016nsss(0)='1'  OR cVar2S5S30P064P062nsss(0)='1'  OR cVar2S6S30P064N062P066nsss(0)='1'  OR cVar2S7S30N064P062nsss(0)='1'  )then
          oVar1S170(0) <='1';
          else
          oVar1S170(0) <='0';
          end if;
        if(cVar2S8S30P031nsss(0)='1'  OR cVar2S9S30N031P062P033nsss(0)='1'  OR cVar2S10S30P052P050nsss(0)='1'  OR cVar2S11S30N052P062P009nsss(0)='1'  )then
          oVar1S171(0) <='1';
          else
          oVar1S171(0) <='0';
          end if;
        if(cVar2S12S30P014P067nsss(0)='1'  OR cVar2S13S30P005P011P004nsss(0)='1'  OR cVar2S14S30P005P011P012nsss(0)='1'  OR cVar2S15S30P011P002P035nsss(0)='1'  )then
          oVar1S172(0) <='1';
          else
          oVar1S172(0) <='0';
          end if;
        if(cVar2S16S30N011P026P068nsss(0)='1'  OR cVar2S17S30N011N026P058nsss(0)='1'  OR cVar2S18S30P034P008P062nsss(0)='1'  OR cVar2S19S30P046P015nsss(0)='1'  )then
          oVar1S173(0) <='1';
          else
          oVar1S173(0) <='0';
          end if;
        if(cVar2S0S31P014P059nsss(0)='1'  OR cVar2S1S31P034P004nsss(0)='1'  OR cVar2S2S31P067P015nsss(0)='1'  OR cVar2S3S31P009nsss(0)='1'  )then
          oVar1S175(0) <='1';
          else
          oVar1S175(0) <='0';
          end if;
        if(cVar2S4S31P052nsss(0)='1'  OR cVar2S5S31N052P008nsss(0)='1'  OR cVar2S6S31N052N008P010nsss(0)='1'  OR cVar2S7S31P021nsss(0)='1'  )then
          oVar1S176(0) <='1';
          else
          oVar1S176(0) <='0';
          end if;
        if(cVar2S8S31N021P002nsss(0)='1'  OR cVar2S9S31N021N002P004nsss(0)='1'  OR cVar2S10S31P038P044P042nsss(0)='1'  OR cVar2S11S31P038P010nsss(0)='1'  )then
          oVar1S177(0) <='1';
          else
          oVar1S177(0) <='0';
          end if;
        if(cVar2S12S31P064nsss(0)='1'  OR cVar2S13S31P064P063nsss(0)='1'  OR cVar2S14S31P069nsss(0)='1'  OR cVar2S15S31N069P064P017nsss(0)='1'  )then
          oVar1S178(0) <='1';
          else
          oVar1S178(0) <='0';
          end if;
        if(cVar2S16S31P034P008P015nsss(0)='1'  OR cVar2S17S31P063P014P069nsss(0)='1'  )then
          oVar1S179(0) <='1';
          else
          oVar1S179(0) <='0';
          end if;
        if(cVar2S0S32P068P005nsss(0)='1'  OR cVar2S1S32N068P055nsss(0)='1'  OR cVar2S2S32N068N055P054nsss(0)='1'  OR cVar2S3S32P062P041P039nsss(0)='1'  )then
          oVar1S180(0) <='1';
          else
          oVar1S180(0) <='0';
          end if;
        if(cVar2S4S32P062N041psss(0)='1'  OR cVar1S5S32P061P033P060P032nsss(0)='1'  OR cVar2S6S32P035P034P013nsss(0)='1'  OR cVar2S7S32N035P065P066nsss(0)='1'  )then
          oVar1S181(0) <='1';
          else
          oVar1S181(0) <='0';
          end if;
        if(cVar2S8S32P013P017nsss(0)='1'  OR cVar2S9S32N013P067P014nsss(0)='1'  OR cVar2S10S32P034P039nsss(0)='1'  OR cVar2S11S32P016P034nsss(0)='1'  )then
          oVar1S182(0) <='1';
          else
          oVar1S182(0) <='0';
          end if;
        if(cVar2S12S32P033P058nsss(0)='1'  OR cVar2S13S32N033P034nsss(0)='1'  OR cVar2S14S32N033N034P035nsss(0)='1'  OR cVar2S15S32P013P063nsss(0)='1'  )then
          oVar1S183(0) <='1';
          else
          oVar1S183(0) <='0';
          end if;
        if(cVar2S16S32P034nsss(0)='1'  OR cVar2S17S32P064nsss(0)='1'  OR cVar2S18S32N064P068P019nsss(0)='1'  OR cVar2S19S32P008P015P014nsss(0)='1'  )then
          oVar1S184(0) <='1';
          else
          oVar1S184(0) <='0';
          end if;
        if(cVar2S20S32P008N015P014nsss(0)='1'  OR cVar2S21S32P011P014P016nsss(0)='1'  )then
          oVar1S185(0) <='1';
          else
          oVar1S185(0) <='0';
          end if;
        if(cVar2S0S33P005P050nsss(0)='1'  OR cVar2S1S33P035P009nsss(0)='1'  OR cVar2S2S33N035P001P053nsss(0)='1'  OR cVar2S3S33P015P017nsss(0)='1'  )then
          oVar1S186(0) <='1';
          else
          oVar1S186(0) <='0';
          end if;
        if(cVar2S4S33P030P019P068nsss(0)='1'  OR cVar2S5S33P030P019P064nsss(0)='1'  OR cVar2S6S33P006P010P019nsss(0)='1'  OR cVar1S7S33N062P041P020nsss(0)='1'  )then
          oVar1S187(0) <='1';
          else
          oVar1S187(0) <='0';
          end if;
        if(cVar2S8S33P051P021nsss(0)='1'  OR cVar2S9S33P051N021P008nsss(0)='1'  OR cVar2S10S33P032P015nsss(0)='1'  OR cVar2S11S33P032N015P013nsss(0)='1'  )then
          oVar1S188(0) <='1';
          else
          oVar1S188(0) <='0';
          end if;
        if(cVar2S12S33P063P034P056nsss(0)='1'  OR cVar2S13S33P063P034P013nsss(0)='1'  OR cVar2S14S33P063P067nsss(0)='1'  OR cVar2S15S33P011P029nsss(0)='1'  )then
          oVar1S189(0) <='1';
          else
          oVar1S189(0) <='0';
          end if;
        if(cVar2S16S33P011N029P069nsss(0)='1'  OR cVar2S17S33N011P044nsss(0)='1'  OR cVar2S18S33P008P012P014nsss(0)='1'  )then
          oVar1S190(0) <='1';
          else
          oVar1S190(0) <='0';
          end if;
        if(cVar2S0S34P005nsss(0)='1'  OR cVar2S1S34P005P017nsss(0)='1'  OR cVar2S2S34P016P018nsss(0)='1'  OR cVar2S3S34P069P051nsss(0)='1'  )then
          oVar1S191(0) <='1';
          else
          oVar1S191(0) <='0';
          end if;
        if(cVar2S4S34N069P032P061nsss(0)='1'  OR cVar2S5S34N069P032P061nsss(0)='1'  OR cVar2S6S34P061P004nsss(0)='1'  OR cVar2S7S34P061N004P015nsss(0)='1'  )then
          oVar1S192(0) <='1';
          else
          oVar1S192(0) <='0';
          end if;
        if(cVar2S8S34P061P018P063nsss(0)='1'  OR cVar1S9S34P011P029P052nsss(0)='1'  OR cVar2S10S34P033P010P019nsss(0)='1'  OR cVar2S11S34P033N010P008nsss(0)='1'  )then
          oVar1S193(0) <='1';
          else
          oVar1S193(0) <='0';
          end if;
        if(cVar2S12S34P019nsss(0)='1'  OR cVar2S13S34P003P015P006nsss(0)='1'  OR cVar2S14S34P003N015P031nsss(0)='1'  OR cVar2S15S34P003P015P018nsss(0)='1'  )then
          oVar1S194(0) <='1';
          else
          oVar1S194(0) <='0';
          end if;
        if(cVar2S16S34P021P007P016nsss(0)='1'  OR cVar2S17S34P069P006P065nsss(0)='1'  )then
          oVar1S195(0) <='1';
          else
          oVar1S195(0) <='0';
          end if;
        if(cVar2S0S35P063P066nsss(0)='1'  OR cVar2S1S35P063N066P065nsss(0)='1'  OR cVar2S2S35P063P035P067nsss(0)='1'  OR cVar2S3S35P002P056P036nsss(0)='1'  )then
          oVar1S196(0) <='1';
          else
          oVar1S196(0) <='0';
          end if;
        if(cVar2S4S35P043P063P019nsss(0)='1'  OR cVar1S5S35P015P022P012P014nsss(0)='1'  OR cVar2S6S35P068P024nsss(0)='1'  OR cVar2S7S35N068P055nsss(0)='1'  )then
          oVar1S197(0) <='1';
          else
          oVar1S197(0) <='0';
          end if;
        if(cVar2S8S35N068N055P014nsss(0)='1'  OR cVar2S9S35P060nsss(0)='1'  OR cVar2S10S35P063P012nsss(0)='1'  OR cVar2S11S35P063P012P014nsss(0)='1'  )then
          oVar1S198(0) <='1';
          else
          oVar1S198(0) <='0';
          end if;
        if(cVar2S12S35N063P065P035nsss(0)='1'  OR cVar2S13S35P020P039nsss(0)='1'  OR cVar2S14S35P020N039P035nsss(0)='1'  OR cVar2S15S35N020P011nsss(0)='1'  )then
          oVar1S199(0) <='1';
          else
          oVar1S199(0) <='0';
          end if;
        if(cVar2S16S35N020N011P006nsss(0)='1'  OR cVar2S17S35P008P012nsss(0)='1'  OR cVar2S18S35N008P062P043nsss(0)='1'  OR cVar2S19S35N008P062P060nsss(0)='1'  )then
          oVar1S200(0) <='1';
          else
          oVar1S200(0) <='0';
          end if;
        if(cVar2S20S35P065P035nsss(0)='1'  )then
          oVar1S201(0) <='1';
          else
          oVar1S201(0) <='0';
          end if;
        if(cVar2S0S36P060P066nsss(0)='1'  OR cVar2S1S36P060P066P012nsss(0)='1'  OR cVar2S2S36P060P014nsss(0)='1'  OR cVar2S3S36P016P067nsss(0)='1'  )then
          oVar1S202(0) <='1';
          else
          oVar1S202(0) <='0';
          end if;
        if(cVar2S4S36P016N067P068nsss(0)='1'  OR cVar2S5S36P016P066nsss(0)='1'  OR cVar2S6S36P034P029nsss(0)='1'  OR cVar2S7S36P034P029P052nsss(0)='1'  )then
          oVar1S203(0) <='1';
          else
          oVar1S203(0) <='0';
          end if;
        if(cVar2S8S36P034P029nsss(0)='1'  OR cVar2S9S36P034N029P061nsss(0)='1'  OR cVar2S10S36P064P066nsss(0)='1'  OR cVar2S11S36N064P013P019nsss(0)='1'  )then
          oVar1S204(0) <='1';
          else
          oVar1S204(0) <='0';
          end if;
        if(cVar2S12S36P004P024P012nsss(0)='1'  OR cVar2S13S36P013P041P062nsss(0)='1'  OR cVar2S14S36N013P031P041nsss(0)='1'  OR cVar2S15S36N013P031P066nsss(0)='1'  )then
          oVar1S205(0) <='1';
          else
          oVar1S205(0) <='0';
          end if;
        if(cVar1S16S36P011P004P029P054nsss(0)='1'  OR cVar2S17S36P051nsss(0)='1'  OR cVar2S18S36N051P052nsss(0)='1'  OR cVar2S19S36P021P039P028nsss(0)='1'  )then
          oVar1S206(0) <='1';
          else
          oVar1S206(0) <='0';
          end if;
        if(cVar2S20S36P000P065P015nsss(0)='1'  OR cVar2S21S36P003P008P064nsss(0)='1'  )then
          oVar1S207(0) <='1';
          else
          oVar1S207(0) <='0';
          end if;
        if(cVar2S0S37P045P053P000nsss(0)='1'  OR cVar2S1S37P045N053P051nsss(0)='1'  OR cVar2S2S37P045P068nsss(0)='1'  OR cVar2S3S37P036P054P016nsss(0)='1'  )then
          oVar1S208(0) <='1';
          else
          oVar1S208(0) <='0';
          end if;
        if(cVar1S4S37P015P031P022P012nsss(0)='1'  OR cVar2S5S37P010nsss(0)='1'  OR cVar2S6S37N010P059nsss(0)='1'  OR cVar1S7S37N015P065P007P052nsss(0)='1'  )then
          oVar1S209(0) <='1';
          else
          oVar1S209(0) <='0';
          end if;
        if(cVar2S8S37P050P060P063nsss(0)='1'  OR cVar2S9S37P050P060P062nsss(0)='1'  OR cVar2S10S37P010P018nsss(0)='1'  OR cVar1S11S37N015N065P022P043nsss(0)='1'  )then
          oVar1S210(0) <='1';
          else
          oVar1S210(0) <='0';
          end if;
        if(cVar2S12S37P024P069P004nsss(0)='1'  OR cVar2S13S37P062P052nsss(0)='1'  OR cVar2S14S37P062N052P061nsss(0)='1'  OR cVar2S15S37N062P063P010nsss(0)='1'  )then
          oVar1S211(0) <='1';
          else
          oVar1S211(0) <='0';
          end if;
        if(cVar2S16S37P045P005nsss(0)='1'  OR cVar2S17S37P045N005P014nsss(0)='1'  OR cVar2S18S37N045P009nsss(0)='1'  )then
          oVar1S212(0) <='1';
          else
          oVar1S212(0) <='0';
          end if;
        if(cVar2S0S38P069P060P016nsss(0)='1'  OR cVar2S1S38P069N060psss(0)='1'  OR cVar2S2S38P069P067P032nsss(0)='1'  OR cVar2S3S38P067P035nsss(0)='1'  )then
          oVar1S213(0) <='1';
          else
          oVar1S213(0) <='0';
          end if;
        if(cVar2S4S38P067P035P063nsss(0)='1'  OR cVar2S5S38N067P032nsss(0)='1'  OR cVar2S6S38N067P032P012nsss(0)='1'  OR cVar2S7S38P000P034nsss(0)='1'  )then
          oVar1S214(0) <='1';
          else
          oVar1S214(0) <='0';
          end if;
        if(cVar2S8S38P051P066nsss(0)='1'  OR cVar2S9S38P051P014P049nsss(0)='1'  OR cVar1S10S38P006P024P014P047nsss(0)='1'  OR cVar2S11S38P049P000nsss(0)='1'  )then
          oVar1S215(0) <='1';
          else
          oVar1S215(0) <='0';
          end if;
        if(cVar2S12S38P049N000P017nsss(0)='1'  OR cVar2S13S38P026P015P066nsss(0)='1'  OR cVar2S14S38P011P013nsss(0)='1'  OR cVar2S15S38P005P000P067nsss(0)='1'  )then
          oVar1S216(0) <='1';
          else
          oVar1S216(0) <='0';
          end if;
        if(cVar2S16S38P005P010nsss(0)='1'  OR cVar2S17S38P017P010P063nsss(0)='1'  OR cVar2S18S38P068P065nsss(0)='1'  )then
          oVar1S217(0) <='1';
          else
          oVar1S217(0) <='0';
          end if;
        if(cVar2S0S39P065P068P062nsss(0)='1'  OR cVar2S1S39P065P068P012nsss(0)='1'  OR cVar2S2S39N065P063nsss(0)='1'  OR cVar2S3S39N065P063P064nsss(0)='1'  )then
          oVar1S218(0) <='1';
          else
          oVar1S218(0) <='0';
          end if;
        if(cVar2S4S39P045nsss(0)='1'  OR cVar2S5S39P035P008P015nsss(0)='1'  OR cVar2S6S39P022P068P031nsss(0)='1'  OR cVar2S7S39P022P068P061nsss(0)='1'  )then
          oVar1S219(0) <='1';
          else
          oVar1S219(0) <='0';
          end if;
        if(cVar2S8S39P022P014P018nsss(0)='1'  OR cVar2S9S39P036nsss(0)='1'  OR cVar2S10S39P069P060P036nsss(0)='1'  OR cVar2S11S39P069N060psss(0)='1'  )then
          oVar1S220(0) <='1';
          else
          oVar1S220(0) <='0';
          end if;
        if(cVar2S12S39P032P037P041nsss(0)='1'  OR cVar2S13S39P032P012P018nsss(0)='1'  OR cVar2S14S39P047nsss(0)='1'  OR cVar2S15S39N047P013P015nsss(0)='1'  )then
          oVar1S221(0) <='1';
          else
          oVar1S221(0) <='0';
          end if;
        if(cVar2S16S39P021nsss(0)='1'  OR cVar2S17S39P014P013P018nsss(0)='1'  OR cVar2S18S39P053nsss(0)='1'  )then
          oVar1S222(0) <='1';
          else
          oVar1S222(0) <='0';
          end if;
        if(cVar2S0S40P056nsss(0)='1'  OR cVar2S1S40N056P018nsss(0)='1'  OR cVar2S2S40N056P018P015nsss(0)='1'  OR cVar2S3S40P010nsss(0)='1'  )then
          oVar1S223(0) <='1';
          else
          oVar1S223(0) <='0';
          end if;
        if(cVar2S4S40N010P057nsss(0)='1'  OR cVar2S5S40N010N057P016nsss(0)='1'  OR cVar2S6S40P055P027P009nsss(0)='1'  OR cVar2S7S40P055N027psss(0)='1'  )then
          oVar1S224(0) <='1';
          else
          oVar1S224(0) <='0';
          end if;
        if(cVar2S8S40P055P013P016nsss(0)='1'  OR cVar2S9S40P031P013nsss(0)='1'  OR cVar2S10S40N031P000P010nsss(0)='1'  OR cVar2S11S40P036P037nsss(0)='1'  )then
          oVar1S225(0) <='1';
          else
          oVar1S225(0) <='0';
          end if;
        if(cVar2S12S40P036N037P061nsss(0)='1'  OR cVar2S13S40P018P013nsss(0)='1'  OR cVar2S14S40P018N013P019nsss(0)='1'  OR cVar2S15S40P013nsss(0)='1'  )then
          oVar1S226(0) <='1';
          else
          oVar1S226(0) <='0';
          end if;
        if(cVar2S16S40P008P060nsss(0)='1'  OR cVar2S17S40P008N060P034nsss(0)='1'  OR cVar2S18S40P069P035P012nsss(0)='1'  OR cVar2S19S40P069P037P067nsss(0)='1'  )then
          oVar1S227(0) <='1';
          else
          oVar1S227(0) <='0';
          end if;
        if(cVar2S20S40P069N037P035nsss(0)='1'  OR cVar2S21S40P017P018nsss(0)='1'  OR cVar2S22S40P003P043nsss(0)='1'  )then
          oVar1S228(0) <='1';
          else
          oVar1S228(0) <='0';
          end if;
        if(cVar1S0S41P035P015P027P050nsss(0)='1'  OR cVar2S1S41P014P048nsss(0)='1'  OR cVar2S2S41P043nsss(0)='1'  OR cVar2S3S41N043P017P010nsss(0)='1'  )then
          oVar1S229(0) <='1';
          else
          oVar1S229(0) <='0';
          end if;
        if(cVar2S4S41P043P056P004nsss(0)='1'  OR cVar2S5S41P043N056P047nsss(0)='1'  OR cVar2S6S41P043P005nsss(0)='1'  OR cVar2S7S41P043N005P024nsss(0)='1'  )then
          oVar1S230(0) <='1';
          else
          oVar1S230(0) <='0';
          end if;
        if(cVar2S8S41P004P012nsss(0)='1'  OR cVar2S9S41P004P012P037nsss(0)='1'  OR cVar2S10S41P059P056nsss(0)='1'  OR cVar2S11S41P059N056P004nsss(0)='1'  )then
          oVar1S231(0) <='1';
          else
          oVar1S231(0) <='0';
          end if;
        if(cVar2S12S41N059P012P013nsss(0)='1'  OR cVar2S13S41N059N012P003nsss(0)='1'  OR cVar2S14S41P009P008P016nsss(0)='1'  OR cVar2S15S41P012P067nsss(0)='1'  )then
          oVar1S232(0) <='1';
          else
          oVar1S232(0) <='0';
          end if;
        if(cVar2S16S41N012P009P011nsss(0)='1'  OR cVar2S17S41P034P022P059nsss(0)='1'  OR cVar2S18S41P034P037P018nsss(0)='1'  OR cVar2S19S41P065P012P015nsss(0)='1'  )then
          oVar1S233(0) <='1';
          else
          oVar1S233(0) <='0';
          end if;
        if(cVar2S0S42P027P050nsss(0)='1'  OR cVar2S1S42P027N050P049nsss(0)='1'  OR cVar2S2S42N027P049P007nsss(0)='1'  OR cVar2S3S42N027P049P047nsss(0)='1'  )then
          oVar1S235(0) <='1';
          else
          oVar1S235(0) <='0';
          end if;
        if(cVar2S4S42P040nsss(0)='1'  OR cVar2S5S42N040P010P007nsss(0)='1'  OR cVar2S6S42P033P007P003nsss(0)='1'  OR cVar2S7S42P067P058P037nsss(0)='1'  )then
          oVar1S236(0) <='1';
          else
          oVar1S236(0) <='0';
          end if;
        if(cVar2S8S42P067P066P069nsss(0)='1'  OR cVar2S9S42P067P066P008nsss(0)='1'  OR cVar2S10S42P066P035nsss(0)='1'  OR cVar2S11S42P066N035P008nsss(0)='1'  )then
          oVar1S237(0) <='1';
          else
          oVar1S237(0) <='0';
          end if;
        if(cVar2S12S42P066P037nsss(0)='1'  OR cVar2S13S42P065P036P066nsss(0)='1'  OR cVar2S14S42P065P018P068nsss(0)='1'  OR cVar2S15S42P065N018P035nsss(0)='1'  )then
          oVar1S238(0) <='1';
          else
          oVar1S238(0) <='0';
          end if;
        if(cVar2S16S42P013P019P012nsss(0)='1'  OR cVar2S17S42P013P019P018nsss(0)='1'  OR cVar2S18S42P013P016P014nsss(0)='1'  OR cVar2S19S42P065P018P010nsss(0)='1'  )then
          oVar1S239(0) <='1';
          else
          oVar1S239(0) <='0';
          end if;
        if(cVar2S20S42P027nsss(0)='1'  )then
          oVar1S240(0) <='1';
          else
          oVar1S240(0) <='0';
          end if;
        if(cVar2S0S43P009P032P033nsss(0)='1'  OR cVar2S1S43P009N032psss(0)='1'  OR cVar2S2S43P009P004P067nsss(0)='1'  OR cVar2S3S43P008P002P050nsss(0)='1'  )then
          oVar1S241(0) <='1';
          else
          oVar1S241(0) <='0';
          end if;
        if(cVar2S4S43P008P018P059nsss(0)='1'  OR cVar2S5S43P016P019nsss(0)='1'  OR cVar2S6S43P057P063P006nsss(0)='1'  OR cVar1S7S43N015P027P048nsss(0)='1'  )then
          oVar1S242(0) <='1';
          else
          oVar1S242(0) <='0';
          end if;
        if(cVar2S8S43P049nsss(0)='1'  OR cVar2S9S43N049P035P003nsss(0)='1'  OR cVar2S10S43P018P011P010nsss(0)='1'  OR cVar2S11S43P010nsss(0)='1'  )then
          oVar1S243(0) <='1';
          else
          oVar1S243(0) <='0';
          end if;
        if(cVar2S12S43N010P057nsss(0)='1'  OR cVar2S13S43N010N057P016nsss(0)='1'  OR cVar2S14S43P021nsss(0)='1'  OR cVar2S15S43N021P020nsss(0)='1'  )then
          oVar1S244(0) <='1';
          else
          oVar1S244(0) <='0';
          end if;
        if(cVar2S16S43N021N020P018nsss(0)='1'  OR cVar2S17S43P038P002P029nsss(0)='1'  )then
          oVar1S245(0) <='1';
          else
          oVar1S245(0) <='0';
          end if;
        if(cVar1S0S44P015P027P000P048nsss(0)='1'  OR cVar2S1S44P005P035nsss(0)='1'  OR cVar2S2S44P014P066nsss(0)='1'  OR cVar2S3S44N014P032nsss(0)='1'  )then
          oVar1S246(0) <='1';
          else
          oVar1S246(0) <='0';
          end if;
        if(cVar2S4S44N014P032P012nsss(0)='1'  OR cVar2S5S44P067P032P037nsss(0)='1'  OR cVar2S6S44P067N032P051nsss(0)='1'  OR cVar2S7S44P067P012P019nsss(0)='1'  )then
          oVar1S247(0) <='1';
          else
          oVar1S247(0) <='0';
          end if;
        if(cVar2S8S44P031nsss(0)='1'  OR cVar2S9S44N031P061P063nsss(0)='1'  OR cVar2S10S44N031N061P011nsss(0)='1'  OR cVar2S11S44P000P036P069nsss(0)='1'  )then
          oVar1S248(0) <='1';
          else
          oVar1S248(0) <='0';
          end if;
        if(cVar2S12S44N000P068P055nsss(0)='1'  OR cVar2S13S44N000N068P011nsss(0)='1'  OR cVar2S14S44P031P065P047nsss(0)='1'  OR cVar2S15S44P031P065P019nsss(0)='1'  )then
          oVar1S249(0) <='1';
          else
          oVar1S249(0) <='0';
          end if;
        if(cVar2S16S44P031P034nsss(0)='1'  OR cVar2S17S44P008P004P037nsss(0)='1'  OR cVar2S18S44P057P000nsss(0)='1'  OR cVar2S19S44P063P016P009nsss(0)='1'  )then
          oVar1S250(0) <='1';
          else
          oVar1S250(0) <='0';
          end if;
        if(cVar2S20S44P063N016P014nsss(0)='1'  OR cVar2S21S44P006P035nsss(0)='1'  OR cVar2S22S44P012nsss(0)='1'  )then
          oVar1S251(0) <='1';
          else
          oVar1S251(0) <='0';
          end if;
        if(cVar2S0S45P000P016nsss(0)='1'  OR cVar2S1S45P000N016P067nsss(0)='1'  OR cVar2S2S45N000P069P032nsss(0)='1'  OR cVar2S3S45N000P069P067nsss(0)='1'  )then
          oVar1S252(0) <='1';
          else
          oVar1S252(0) <='0';
          end if;
        if(cVar2S4S45P064nsss(0)='1'  OR cVar2S5S45N064P069P013nsss(0)='1'  OR cVar1S6S45P015P018P030P069nsss(0)='1'  OR cVar2S7S45N057P016P014nsss(0)='1'  )then
          oVar1S253(0) <='1';
          else
          oVar1S253(0) <='0';
          end if;
        if(cVar2S8S45P034P064nsss(0)='1'  OR cVar2S9S45P034N064P066nsss(0)='1'  OR cVar2S10S45N034psss(0)='1'  OR cVar2S11S45P064P029P069nsss(0)='1'  )then
          oVar1S254(0) <='1';
          else
          oVar1S254(0) <='0';
          end if;
        if(cVar2S12S45P064P010nsss(0)='1'  OR cVar2S13S45P014P017P066nsss(0)='1'  OR cVar2S14S45P014N017P047nsss(0)='1'  OR cVar2S15S45N014P027nsss(0)='1'  )then
          oVar1S255(0) <='1';
          else
          oVar1S255(0) <='0';
          end if;
        if(cVar2S16S45N014N027P066nsss(0)='1'  OR cVar2S17S45P025P018nsss(0)='1'  OR cVar2S18S45P013P019nsss(0)='1'  OR cVar2S19S45P057P006nsss(0)='1'  )then
          oVar1S256(0) <='1';
          else
          oVar1S256(0) <='0';
          end if;
        if(cVar2S20S45P053P063P016nsss(0)='1'  OR cVar2S21S45P006P012P016nsss(0)='1'  OR cVar2S22S45P014nsss(0)='1'  )then
          oVar1S257(0) <='1';
          else
          oVar1S257(0) <='0';
          end if;
        if(cVar2S0S46P014nsss(0)='1'  OR cVar2S1S46P031P013nsss(0)='1'  OR cVar2S2S46N031P016P014nsss(0)='1'  OR cVar2S3S46P023nsss(0)='1'  )then
          oVar1S258(0) <='1';
          else
          oVar1S258(0) <='0';
          end if;
        if(cVar2S4S46N023P031nsss(0)='1'  OR cVar2S5S46P060P062nsss(0)='1'  OR cVar2S6S46P060N062P012nsss(0)='1'  OR cVar2S7S46N060P007P059nsss(0)='1'  )then
          oVar1S259(0) <='1';
          else
          oVar1S259(0) <='0';
          end if;
        if(cVar2S8S46N060N007P023nsss(0)='1'  OR cVar2S9S46P049P033P001nsss(0)='1'  OR cVar2S10S46P049P051P069nsss(0)='1'  OR cVar2S11S46P014P045nsss(0)='1'  )then
          oVar1S260(0) <='1';
          else
          oVar1S260(0) <='0';
          end if;
        if(cVar2S12S46P039P010P016nsss(0)='1'  OR cVar2S13S46P069P034nsss(0)='1'  OR cVar2S14S46P069N034P066nsss(0)='1'  OR cVar2S15S46P069P036nsss(0)='1'  )then
          oVar1S261(0) <='1';
          else
          oVar1S261(0) <='0';
          end if;
        if(cVar2S16S46P031nsss(0)='1'  OR cVar2S17S46N031P030nsss(0)='1'  OR cVar2S18S46P057P008P004nsss(0)='1'  OR cVar2S19S46P057P069nsss(0)='1'  )then
          oVar1S262(0) <='1';
          else
          oVar1S262(0) <='0';
          end if;
        if(cVar2S20S46P037P060P062nsss(0)='1'  OR cVar2S21S46N037P069P036nsss(0)='1'  )then
          oVar1S263(0) <='1';
          else
          oVar1S263(0) <='0';
          end if;
        if(cVar2S0S47P059P000P057nsss(0)='1'  OR cVar2S1S47N059P061nsss(0)='1'  OR cVar2S2S47P045P014nsss(0)='1'  OR cVar2S3S47P060P024nsss(0)='1'  )then
          oVar1S264(0) <='1';
          else
          oVar1S264(0) <='0';
          end if;
        if(cVar2S4S47P068P013nsss(0)='1'  OR cVar2S5S47P059nsss(0)='1'  OR cVar2S6S47N059P069P066nsss(0)='1'  OR cVar2S7S47P011nsss(0)='1'  )then
          oVar1S265(0) <='1';
          else
          oVar1S265(0) <='0';
          end if;
        if(cVar2S8S47P013P014nsss(0)='1'  OR cVar2S9S47P010P028nsss(0)='1'  OR cVar2S10S47P010N028P030nsss(0)='1'  OR cVar2S11S47N010P036P014nsss(0)='1'  )then
          oVar1S266(0) <='1';
          else
          oVar1S266(0) <='0';
          end if;
        if(cVar2S12S47N010N036P008nsss(0)='1'  OR cVar2S13S47P059P061P040nsss(0)='1'  OR cVar2S14S47P059P061P018nsss(0)='1'  OR cVar2S15S47P059P033P058nsss(0)='1'  )then
          oVar1S267(0) <='1';
          else
          oVar1S267(0) <='0';
          end if;
        if(cVar2S16S47P002nsss(0)='1'  OR cVar2S17S47N002P054nsss(0)='1'  OR cVar2S18S47N002N054P007nsss(0)='1'  OR cVar2S19S47P066nsss(0)='1'  )then
          oVar1S268(0) <='1';
          else
          oVar1S268(0) <='0';
          end if;
        if(cVar2S20S47P051P061P032nsss(0)='1'  OR cVar2S21S47P051P053P018nsss(0)='1'  )then
          oVar1S269(0) <='1';
          else
          oVar1S269(0) <='0';
          end if;
        if(cVar2S0S48P025nsss(0)='1'  OR cVar2S1S48N025P009P011nsss(0)='1'  OR cVar2S2S48N025N009P006nsss(0)='1'  OR cVar2S3S48P049P047nsss(0)='1'  )then
          oVar1S270(0) <='1';
          else
          oVar1S270(0) <='0';
          end if;
        if(cVar2S4S48P049P009nsss(0)='1'  OR cVar2S5S48P049N009P026nsss(0)='1'  OR cVar2S6S48P032nsss(0)='1'  OR cVar2S7S48P030nsss(0)='1'  )then
          oVar1S271(0) <='1';
          else
          oVar1S271(0) <='0';
          end if;
        if(cVar2S8S48N030P031nsss(0)='1'  OR cVar2S9S48P029P068nsss(0)='1'  OR cVar2S10S48N029P003P032nsss(0)='1'  OR cVar2S11S48P053P020nsss(0)='1'  )then
          oVar1S272(0) <='1';
          else
          oVar1S272(0) <='0';
          end if;
        if(cVar2S12S48P003P064P057nsss(0)='1'  OR cVar2S13S48N003P026P008nsss(0)='1'  OR cVar2S14S48P016P065P018nsss(0)='1'  OR cVar2S15S48P016P067P012nsss(0)='1'  )then
          oVar1S273(0) <='1';
          else
          oVar1S273(0) <='0';
          end if;
        if(cVar2S16S48P034P013nsss(0)='1'  OR cVar2S17S48P034N013P067nsss(0)='1'  )then
          oVar1S274(0) <='1';
          else
          oVar1S274(0) <='0';
          end if;
        if(cVar2S0S49P034P032P015nsss(0)='1'  OR cVar2S1S49N034P028P010nsss(0)='1'  OR cVar2S2S49N034N028psss(0)='1'  OR cVar2S3S49P039P062P061nsss(0)='1'  )then
          oVar1S275(0) <='1';
          else
          oVar1S275(0) <='0';
          end if;
        if(cVar2S4S49P068nsss(0)='1'  OR cVar2S5S49P034P053P018nsss(0)='1'  OR cVar2S6S49P017P037P035nsss(0)='1'  OR cVar2S7S49N017P066nsss(0)='1'  )then
          oVar1S276(0) <='1';
          else
          oVar1S276(0) <='0';
          end if;
        if(cVar2S8S49P066P014nsss(0)='1'  OR cVar2S9S49P013P014nsss(0)='1'  OR cVar1S10S49N019P007P025nsss(0)='1'  OR cVar2S11S49P054P065nsss(0)='1'  )then
          oVar1S277(0) <='1';
          else
          oVar1S277(0) <='0';
          end if;
        if(cVar2S12S49P054P065P034nsss(0)='1'  OR cVar2S13S49P001P033P037nsss(0)='1'  OR cVar2S14S49P001N033P032nsss(0)='1'  OR cVar2S15S49P010P028nsss(0)='1'  )then
          oVar1S278(0) <='1';
          else
          oVar1S278(0) <='0';
          end if;
        if(cVar2S16S49P010N028P030nsss(0)='1'  OR cVar2S17S49N010P036nsss(0)='1'  OR cVar2S18S49N010N036P032nsss(0)='1'  OR cVar2S19S49P030P013P031nsss(0)='1'  )then
          oVar1S279(0) <='1';
          else
          oVar1S279(0) <='0';
          end if;
        if(cVar2S20S49P030P012P014nsss(0)='1'  )then
          oVar1S280(0) <='1';
          else
          oVar1S280(0) <='0';
          end if;
        if(cVar1S0S50P019P014P027P009nsss(0)='1'  OR cVar2S1S50P037P026nsss(0)='1'  OR cVar2S2S50P036nsss(0)='1'  OR cVar2S3S50N036P013P031nsss(0)='1'  )then
          oVar1S281(0) <='1';
          else
          oVar1S281(0) <='0';
          end if;
        if(cVar2S4S50N036P013P010nsss(0)='1'  OR cVar2S5S50P004P029nsss(0)='1'  OR cVar2S6S50P011P006P002nsss(0)='1'  OR cVar2S7S50N011P054P036nsss(0)='1'  )then
          oVar1S282(0) <='1';
          else
          oVar1S282(0) <='0';
          end if;
        if(cVar2S8S50N011P054P018nsss(0)='1'  OR cVar2S9S50P065P006P037nsss(0)='1'  OR cVar1S10S50P019P014P030P035nsss(0)='1'  OR cVar2S11S50P062P039P043nsss(0)='1'  )then
          oVar1S283(0) <='1';
          else
          oVar1S283(0) <='0';
          end if;
        if(cVar2S12S50P062P064P008nsss(0)='1'  OR cVar2S13S50P034P032nsss(0)='1'  OR cVar2S14S50N034P069P012nsss(0)='1'  OR cVar2S15S50P012P068nsss(0)='1'  )then
          oVar1S284(0) <='1';
          else
          oVar1S284(0) <='0';
          end if;
        if(cVar2S16S50P036P010nsss(0)='1'  OR cVar2S17S50N036P008P015nsss(0)='1'  )then
          oVar1S285(0) <='1';
          else
          oVar1S285(0) <='0';
          end if;
        if(cVar2S0S51P040P038P021nsss(0)='1'  OR cVar2S1S51P040P066nsss(0)='1'  OR cVar2S2S51P012P013P016nsss(0)='1'  OR cVar2S3S51P012P068nsss(0)='1'  )then
          oVar1S286(0) <='1';
          else
          oVar1S286(0) <='0';
          end if;
        if(cVar2S4S51P036P010nsss(0)='1'  OR cVar2S5S51N036P008P016nsss(0)='1'  OR cVar2S6S51N036N008P066nsss(0)='1'  OR cVar2S7S51P012P050P004nsss(0)='1'  )then
          oVar1S287(0) <='1';
          else
          oVar1S287(0) <='0';
          end if;
        if(cVar2S8S51N012P050P014nsss(0)='1'  OR cVar2S9S51N012N050P061nsss(0)='1'  OR cVar2S10S51P061P033P002nsss(0)='1'  OR cVar1S11S51N019N017P005P023nsss(0)='1'  )then
          oVar1S288(0) <='1';
          else
          oVar1S288(0) <='0';
          end if;
        if(cVar2S12S51P021nsss(0)='1'  OR cVar2S13S51N021P006P054nsss(0)='1'  OR cVar2S14S51P030P046nsss(0)='1'  OR cVar2S15S51P030N046P031nsss(0)='1'  )then
          oVar1S289(0) <='1';
          else
          oVar1S289(0) <='0';
          end if;
        if(cVar2S16S51P030P057nsss(0)='1'  OR cVar2S17S51P030N057P015nsss(0)='1'  OR cVar2S18S51P057P010nsss(0)='1'  OR cVar2S19S51N057P000P037nsss(0)='1'  )then
          oVar1S290(0) <='1';
          else
          oVar1S290(0) <='0';
          end if;
        if(cVar2S20S51N057N000P013nsss(0)='1'  )then
          oVar1S291(0) <='1';
          else
          oVar1S291(0) <='0';
          end if;
        if(cVar2S0S52P004P048nsss(0)='1'  OR cVar2S1S52P004N048P052nsss(0)='1'  OR cVar2S2S52P048P027nsss(0)='1'  OR cVar2S3S52P048P027P009nsss(0)='1'  )then
          oVar1S292(0) <='1';
          else
          oVar1S292(0) <='0';
          end if;
        if(cVar2S4S52P048P025nsss(0)='1'  OR cVar2S5S52P048N025P046nsss(0)='1'  OR cVar2S6S52P014nsss(0)='1'  OR cVar2S7S52P016P017nsss(0)='1'  )then
          oVar1S293(0) <='1';
          else
          oVar1S293(0) <='0';
          end if;
        if(cVar2S8S52N016P057nsss(0)='1'  OR cVar2S9S52P058nsss(0)='1'  OR cVar2S10S52N058P014nsss(0)='1'  OR cVar2S11S52P030P014nsss(0)='1'  )then
          oVar1S294(0) <='1';
          else
          oVar1S294(0) <='0';
          end if;
        if(cVar2S12S52N030P000P036nsss(0)='1'  OR cVar2S13S52N030N000P002nsss(0)='1'  OR cVar2S14S52P050P059nsss(0)='1'  OR cVar2S15S52P010P012nsss(0)='1'  )then
          oVar1S295(0) <='1';
          else
          oVar1S295(0) <='0';
          end if;
        if(cVar2S16S52N010P009P011nsss(0)='1'  OR cVar2S17S52P016nsss(0)='1'  OR cVar2S18S52P017P037nsss(0)='1'  OR cVar2S19S52N017P012P066nsss(0)='1'  )then
          oVar1S296(0) <='1';
          else
          oVar1S296(0) <='0';
          end if;
        if(cVar2S20S52P017nsss(0)='1'  )then
          oVar1S297(0) <='1';
          else
          oVar1S297(0) <='0';
          end if;
        if(cVar2S0S53P010P046nsss(0)='1'  OR cVar2S1S53P010P012P028nsss(0)='1'  OR cVar2S2S53P026nsss(0)='1'  OR cVar2S3S53N026P037P014nsss(0)='1'  )then
          oVar1S298(0) <='1';
          else
          oVar1S298(0) <='0';
          end if;
        if(cVar2S4S53P008nsss(0)='1'  OR cVar2S5S53N008P047nsss(0)='1'  OR cVar2S6S53P060P015nsss(0)='1'  OR cVar2S7S53N060P064P017nsss(0)='1'  )then
          oVar1S299(0) <='1';
          else
          oVar1S299(0) <='0';
          end if;
        if(cVar2S8S53P066P014nsss(0)='1'  OR cVar1S9S53N019P050P021P027nsss(0)='1'  OR cVar2S10S53P039P007P032nsss(0)='1'  OR cVar2S11S53P060nsss(0)='1'  )then
          oVar1S300(0) <='1';
          else
          oVar1S300(0) <='0';
          end if;
        if(cVar2S12S53N060P069nsss(0)='1'  OR cVar2S13S53N060N069P016nsss(0)='1'  OR cVar2S14S53P042nsss(0)='1'  OR cVar2S15S53N042P045nsss(0)='1'  )then
          oVar1S301(0) <='1';
          else
          oVar1S301(0) <='0';
          end if;
        if(cVar2S16S53P042P044P046nsss(0)='1'  OR cVar2S17S53P042P065nsss(0)='1'  )then
          oVar1S302(0) <='1';
          else
          oVar1S302(0) <='0';
          end if;
        if(cVar2S0S54P050P004nsss(0)='1'  OR cVar2S1S54P042P065P064nsss(0)='1'  OR cVar2S2S54P042N065psss(0)='1'  OR cVar2S3S54P034P037nsss(0)='1'  )then
          oVar1S303(0) <='1';
          else
          oVar1S303(0) <='0';
          end if;
        if(cVar2S4S54P034P037P068nsss(0)='1'  OR cVar2S5S54P035P052nsss(0)='1'  OR cVar2S6S54P033nsss(0)='1'  OR cVar2S7S54N033P011P063nsss(0)='1'  )then
          oVar1S304(0) <='1';
          else
          oVar1S304(0) <='0';
          end if;
        if(cVar2S8S54P055nsss(0)='1'  OR cVar2S9S54N055P062P035nsss(0)='1'  OR cVar2S10S54N055N062P011nsss(0)='1'  OR cVar2S11S54P002P016P013nsss(0)='1'  )then
          oVar1S305(0) <='1';
          else
          oVar1S305(0) <='0';
          end if;
        if(cVar2S12S54P033nsss(0)='1'  OR cVar2S13S54P064P011nsss(0)='1'  OR cVar2S14S54P064P011P015nsss(0)='1'  OR cVar2S15S54P064P011P069nsss(0)='1'  )then
          oVar1S306(0) <='1';
          else
          oVar1S306(0) <='0';
          end if;
        if(cVar2S16S54P064P058P003nsss(0)='1'  OR cVar2S17S54N064P028nsss(0)='1'  OR cVar2S18S54N064N028P044nsss(0)='1'  OR cVar2S19S54P031nsss(0)='1'  )then
          oVar1S307(0) <='1';
          else
          oVar1S307(0) <='0';
          end if;
        if(cVar2S20S54N031P032nsss(0)='1'  OR cVar2S21S54P060nsss(0)='1'  OR cVar2S22S54N060P064P012nsss(0)='1'  OR cVar2S23S54P066P014nsss(0)='1'  )then
          oVar1S308(0) <='1';
          else
          oVar1S308(0) <='0';
          end if;
        if(cVar2S24S54P013P014nsss(0)='1'  )then
          oVar1S309(0) <='1';
          else
          oVar1S309(0) <='0';
          end if;
        if(cVar2S0S55P000P037nsss(0)='1'  OR cVar2S1S55P000N037P002nsss(0)='1'  OR cVar2S2S55N000P004P043nsss(0)='1'  OR cVar2S3S55N000P004P036nsss(0)='1'  )then
          oVar1S310(0) <='1';
          else
          oVar1S310(0) <='0';
          end if;
        if(cVar2S4S55P019P016nsss(0)='1'  OR cVar2S5S55P006P036nsss(0)='1'  OR cVar2S6S55P006N036P018nsss(0)='1'  OR cVar2S7S55P049P014nsss(0)='1'  )then
          oVar1S311(0) <='1';
          else
          oVar1S311(0) <='0';
          end if;
        if(cVar2S8S55P000P036P008nsss(0)='1'  OR cVar2S9S55P006P055P008nsss(0)='1'  OR cVar2S10S55P054P065nsss(0)='1'  OR cVar2S11S55P041P020nsss(0)='1'  )then
          oVar1S312(0) <='1';
          else
          oVar1S312(0) <='0';
          end if;
        if(cVar2S12S55P041P020P019nsss(0)='1'  OR cVar2S13S55P008nsss(0)='1'  OR cVar2S14S55N008P069P060nsss(0)='1'  OR cVar2S15S55P009P011P066nsss(0)='1'  )then
          oVar1S313(0) <='1';
          else
          oVar1S313(0) <='0';
          end if;
        if(cVar2S16S55P065P010P067nsss(0)='1'  OR cVar2S17S55N065P016nsss(0)='1'  OR cVar2S18S55N065P016P036nsss(0)='1'  OR cVar2S19S55P066P024P019nsss(0)='1'  )then
          oVar1S314(0) <='1';
          else
          oVar1S314(0) <='0';
          end if;
        if(cVar2S20S55P022nsss(0)='1'  OR cVar2S21S55N022P016P036nsss(0)='1'  OR cVar2S22S55P042P044P033nsss(0)='1'  OR cVar2S23S55P042P005nsss(0)='1'  )then
          oVar1S315(0) <='1';
          else
          oVar1S315(0) <='0';
          end if;
        if(cVar2S24S55P042N005P012nsss(0)='1'  )then
          oVar1S316(0) <='1';
          else
          oVar1S316(0) <='0';
          end if;
        if(cVar2S0S56P063P008nsss(0)='1'  OR cVar2S1S56N063P067P010nsss(0)='1'  OR cVar2S2S56N063N067P010nsss(0)='1'  OR cVar2S3S56P027P009nsss(0)='1'  )then
          oVar1S317(0) <='1';
          else
          oVar1S317(0) <='0';
          end if;
        if(cVar2S4S56P027N009P013nsss(0)='1'  OR cVar2S5S56N027P067nsss(0)='1'  OR cVar2S6S56N027P067P065nsss(0)='1'  OR cVar2S7S56P050P060nsss(0)='1'  )then
          oVar1S318(0) <='1';
          else
          oVar1S318(0) <='0';
          end if;
        if(cVar2S8S56P000P037nsss(0)='1'  OR cVar2S9S56P000N037P002nsss(0)='1'  OR cVar2S10S56N000P016P069nsss(0)='1'  OR cVar2S11S56P013P019nsss(0)='1'  )then
          oVar1S319(0) <='1';
          else
          oVar1S319(0) <='0';
          end if;
        if(cVar2S12S56P006P067nsss(0)='1'  OR cVar2S13S56P049P014nsss(0)='1'  OR cVar2S14S56P016P018nsss(0)='1'  OR cVar2S15S56P016psss(0)='1'  )then
          oVar1S320(0) <='1';
          else
          oVar1S320(0) <='0';
          end if;
        if(cVar2S16S56P064P051nsss(0)='1'  OR cVar2S17S56N064P034P056nsss(0)='1'  OR cVar1S18S56P068P009P024P006nsss(0)='1'  OR cVar2S19S56P016P014P018nsss(0)='1'  )then
          oVar1S321(0) <='1';
          else
          oVar1S321(0) <='0';
          end if;
        if(cVar2S20S56P050nsss(0)='1'  OR cVar2S21S56N050P000P011nsss(0)='1'  )then
          oVar1S322(0) <='1';
          else
          oVar1S322(0) <='0';
          end if;
        if(cVar2S0S57P067P013P063nsss(0)='1'  OR cVar2S1S57P067N013psss(0)='1'  OR cVar2S2S57P067P033P014nsss(0)='1'  OR cVar2S3S57P013P018P058nsss(0)='1'  )then
          oVar1S323(0) <='1';
          else
          oVar1S323(0) <='0';
          end if;
        if(cVar2S4S57P013N018P060nsss(0)='1'  OR cVar2S5S57P013P017P018nsss(0)='1'  OR cVar2S6S57P013P017P024nsss(0)='1'  OR cVar2S7S57P012P013P010nsss(0)='1'  )then
          oVar1S324(0) <='1';
          else
          oVar1S324(0) <='0';
          end if;
        if(cVar2S8S57P012P013P014nsss(0)='1'  OR cVar2S9S57P012P016P010nsss(0)='1'  OR cVar2S10S57P066P065nsss(0)='1'  OR cVar2S11S57P006P035nsss(0)='1'  )then
          oVar1S325(0) <='1';
          else
          oVar1S325(0) <='0';
          end if;
        if(cVar2S12S57P049nsss(0)='1'  OR cVar2S13S57P004nsss(0)='1'  OR cVar2S14S57P013P014P063nsss(0)='1'  OR cVar2S15S57P009nsss(0)='1'  )then
          oVar1S326(0) <='1';
          else
          oVar1S326(0) <='0';
          end if;
        if(cVar2S16S57N009P003nsss(0)='1'  OR cVar2S17S57P066P003nsss(0)='1'  OR cVar2S18S57N066P035nsss(0)='1'  OR cVar2S19S57N066N035P020nsss(0)='1'  )then
          oVar1S327(0) <='1';
          else
          oVar1S327(0) <='0';
          end if;
        if(cVar2S20S57P024P002P013nsss(0)='1'  )then
          oVar1S328(0) <='1';
          else
          oVar1S328(0) <='0';
          end if;
        if(cVar2S0S58P004P022nsss(0)='1'  OR cVar2S1S58P004N022P016nsss(0)='1'  OR cVar2S2S58N004P042nsss(0)='1'  OR cVar2S3S58N004P042P005nsss(0)='1'  )then
          oVar1S329(0) <='1';
          else
          oVar1S329(0) <='0';
          end if;
        if(cVar2S4S58P043P003P007nsss(0)='1'  OR cVar2S5S58P043N003P000nsss(0)='1'  OR cVar2S6S58P043P045nsss(0)='1'  OR cVar2S7S58P019P036nsss(0)='1'  )then
          oVar1S330(0) <='1';
          else
          oVar1S330(0) <='0';
          end if;
        if(cVar2S8S58P019N036P013nsss(0)='1'  OR cVar2S9S58P019P017P016nsss(0)='1'  OR cVar2S10S58P013P012nsss(0)='1'  OR cVar2S11S58P053P024P011nsss(0)='1'  )then
          oVar1S331(0) <='1';
          else
          oVar1S331(0) <='0';
          end if;
        if(cVar2S12S58N053P051P069nsss(0)='1'  OR cVar2S13S58N053P051P008nsss(0)='1'  OR cVar2S14S58P009P014P019nsss(0)='1'  OR cVar2S15S58P030nsss(0)='1'  )then
          oVar1S332(0) <='1';
          else
          oVar1S332(0) <='0';
          end if;
        if(cVar2S16S58P061P033nsss(0)='1'  OR cVar2S17S58P061N033P019nsss(0)='1'  OR cVar2S18S58P043nsss(0)='1'  OR cVar2S19S58P006nsss(0)='1'  )then
          oVar1S333(0) <='1';
          else
          oVar1S333(0) <='0';
          end if;
        if(cVar2S20S58P014P017nsss(0)='1'  OR cVar2S21S58N014P062nsss(0)='1'  OR cVar2S22S58P032nsss(0)='1'  )then
          oVar1S334(0) <='1';
          else
          oVar1S334(0) <='0';
          end if;
        if(cVar2S0S59P016nsss(0)='1'  OR cVar2S1S59P016P000nsss(0)='1'  OR cVar2S2S59P016N000P058nsss(0)='1'  OR cVar2S3S59P052P062P064nsss(0)='1'  )then
          oVar1S335(0) <='1';
          else
          oVar1S335(0) <='0';
          end if;
        if(cVar2S4S59P052P062P037nsss(0)='1'  OR cVar2S5S59P015nsss(0)='1'  OR cVar2S6S59P024P012P048nsss(0)='1'  OR cVar2S7S59P002P014nsss(0)='1'  )then
          oVar1S336(0) <='1';
          else
          oVar1S336(0) <='0';
          end if;
        if(cVar2S8S59P002P014P012nsss(0)='1'  OR cVar2S9S59P063P068nsss(0)='1'  OR cVar2S10S59N063P016P006nsss(0)='1'  OR cVar2S11S59P014nsss(0)='1'  )then
          oVar1S337(0) <='1';
          else
          oVar1S337(0) <='0';
          end if;
        if(cVar2S12S59P003P005P015nsss(0)='1'  OR cVar2S13S59P003P012P014nsss(0)='1'  OR cVar2S14S59P020nsss(0)='1'  OR cVar2S15S59N020P012P041nsss(0)='1'  )then
          oVar1S338(0) <='1';
          else
          oVar1S338(0) <='0';
          end if;
        if(cVar2S16S59P020P057P030nsss(0)='1'  OR cVar2S17S59P020P002nsss(0)='1'  OR cVar2S18S59P009P007nsss(0)='1'  OR cVar2S19S59P011P014P065nsss(0)='1'  )then
          oVar1S339(0) <='1';
          else
          oVar1S339(0) <='0';
          end if;
        if(cVar2S20S59P009nsss(0)='1'  )then
          oVar1S340(0) <='1';
          else
          oVar1S340(0) <='0';
          end if;
        if(cVar2S0S60P028nsss(0)='1'  OR cVar2S1S60N028P058nsss(0)='1'  OR cVar2S2S60N028N058P042nsss(0)='1'  OR cVar2S3S60P004nsss(0)='1'  )then
          oVar1S341(0) <='1';
          else
          oVar1S341(0) <='0';
          end if;
        if(cVar2S4S60N004P032nsss(0)='1'  OR cVar2S5S60N004N032P028nsss(0)='1'  OR cVar2S6S60P004P045nsss(0)='1'  OR cVar2S7S60P024P034P014nsss(0)='1'  )then
          oVar1S342(0) <='1';
          else
          oVar1S342(0) <='0';
          end if;
        if(cVar2S8S60P009P007P032nsss(0)='1'  OR cVar2S9S60P060nsss(0)='1'  OR cVar2S10S60N060P014P065nsss(0)='1'  OR cVar2S11S60P009nsss(0)='1'  )then
          oVar1S343(0) <='1';
          else
          oVar1S343(0) <='0';
          end if;
        if(cVar1S12S60P018P067P019P056nsss(0)='1'  OR cVar2S13S60P014nsss(0)='1'  OR cVar2S14S60P014P012P069nsss(0)='1'  OR cVar2S15S60P014N012P068nsss(0)='1'  )then
          oVar1S344(0) <='1';
          else
          oVar1S344(0) <='0';
          end if;
        if(cVar2S16S60P051P065P062nsss(0)='1'  OR cVar2S17S60P051N065P026nsss(0)='1'  OR cVar2S18S60P051P015nsss(0)='1'  OR cVar2S19S60P056P000P009nsss(0)='1'  )then
          oVar1S345(0) <='1';
          else
          oVar1S345(0) <='0';
          end if;
        if(cVar2S20S60P056P034P036nsss(0)='1'  OR cVar2S21S60P061P009P068nsss(0)='1'  OR cVar2S22S60P063nsss(0)='1'  )then
          oVar1S346(0) <='1';
          else
          oVar1S346(0) <='0';
          end if;
        if(cVar2S0S61P061P013nsss(0)='1'  OR cVar2S1S61P061N013P060nsss(0)='1'  OR cVar2S2S61N061P031nsss(0)='1'  OR cVar2S3S61N061N031P069nsss(0)='1'  )then
          oVar1S347(0) <='1';
          else
          oVar1S347(0) <='0';
          end if;
        if(cVar2S4S61P056P007P058nsss(0)='1'  OR cVar1S5S61P018P008P024P045nsss(0)='1'  OR cVar2S6S61P014P003nsss(0)='1'  OR cVar2S7S61P014P019P016nsss(0)='1'  )then
          oVar1S348(0) <='1';
          else
          oVar1S348(0) <='0';
          end if;
        if(cVar2S8S61P015P002nsss(0)='1'  OR cVar2S9S61P015P063P068nsss(0)='1'  OR cVar2S10S61P034P008P013nsss(0)='1'  OR cVar2S11S61P034N008psss(0)='1'  )then
          oVar1S349(0) <='1';
          else
          oVar1S349(0) <='0';
          end if;
        if(cVar2S12S61P022nsss(0)='1'  OR cVar2S13S61N022P040nsss(0)='1'  OR cVar2S14S61N022N040P016nsss(0)='1'  OR cVar2S15S61P022P028P010nsss(0)='1'  )then
          oVar1S350(0) <='1';
          else
          oVar1S350(0) <='0';
          end if;
        if(cVar2S16S61P022P043nsss(0)='1'  OR cVar2S17S61P007P069P063nsss(0)='1'  OR cVar2S18S61P007N069P036nsss(0)='1'  OR cVar2S19S61P011P014P017nsss(0)='1'  )then
          oVar1S351(0) <='1';
          else
          oVar1S351(0) <='0';
          end if;
        if(cVar2S20S61P009nsss(0)='1'  )then
          oVar1S352(0) <='1';
          else
          oVar1S352(0) <='0';
          end if;
        if(cVar2S0S62P010P014nsss(0)='1'  OR cVar2S1S62N010P030P053nsss(0)='1'  OR cVar2S2S62P026P054nsss(0)='1'  OR cVar2S3S62N026P053P051nsss(0)='1'  )then
          oVar1S353(0) <='1';
          else
          oVar1S353(0) <='0';
          end if;
        if(cVar2S4S62N026P053P011nsss(0)='1'  OR cVar2S5S62P069P051nsss(0)='1'  OR cVar2S6S62P063P060nsss(0)='1'  OR cVar2S7S62N063P036P009nsss(0)='1'  )then
          oVar1S354(0) <='1';
          else
          oVar1S354(0) <='0';
          end if;
        if(cVar2S8S62P045P061nsss(0)='1'  OR cVar2S9S62P045N061P008nsss(0)='1'  OR cVar2S10S62P045P066P036nsss(0)='1'  OR cVar2S11S62P015nsss(0)='1'  )then
          oVar1S355(0) <='1';
          else
          oVar1S355(0) <='0';
          end if;
        if(cVar2S12S62P057P031nsss(0)='1'  )then
          oVar1S356(0) <='1';
          else
          oVar1S356(0) <='0';
          end if;
        if(cVar2S0S63P014nsss(0)='1'  OR cVar2S1S63P030P006P019nsss(0)='1'  OR cVar2S2S63P012P014nsss(0)='1'  OR cVar2S3S63P012P014P015nsss(0)='1'  )then
          oVar1S357(0) <='1';
          else
          oVar1S357(0) <='0';
          end if;
        if(cVar2S4S63N012P058nsss(0)='1'  OR cVar2S5S63N012N058P016nsss(0)='1'  OR cVar2S6S63P057P054P026nsss(0)='1'  OR cVar2S7S63P057P054P013nsss(0)='1'  )then
          oVar1S358(0) <='1';
          else
          oVar1S358(0) <='0';
          end if;
        if(cVar2S8S63P057P062P054nsss(0)='1'  OR cVar2S9S63P062P069nsss(0)='1'  OR cVar2S10S63P062N069P066nsss(0)='1'  OR cVar2S11S63N062P001nsss(0)='1'  )then
          oVar1S359(0) <='1';
          else
          oVar1S359(0) <='0';
          end if;
        if(cVar2S12S63P016P014nsss(0)='1'  OR cVar2S13S63P030P056P061nsss(0)='1'  OR cVar2S14S63P030P069nsss(0)='1'  OR cVar2S15S63P068P017P055nsss(0)='1'  )then
          oVar1S360(0) <='1';
          else
          oVar1S360(0) <='0';
          end if;
        if(cVar2S16S63P068P017P059nsss(0)='1'  OR cVar2S17S63P059P057P024nsss(0)='1'  )then
          oVar1S361(0) <='1';
          else
          oVar1S361(0) <='0';
          end if;
        if(cVar2S0S64P010P067nsss(0)='1'  OR cVar2S1S64N010P006P053nsss(0)='1'  OR cVar2S2S64P041P020nsss(0)='1'  OR cVar2S3S64P041N020P021nsss(0)='1'  )then
          oVar1S362(0) <='1';
          else
          oVar1S362(0) <='0';
          end if;
        if(cVar2S4S64N041P020P002nsss(0)='1'  OR cVar2S5S64N041P020P040nsss(0)='1'  OR cVar2S6S64P036P010nsss(0)='1'  OR cVar2S7S64P009P012P013nsss(0)='1'  )then
          oVar1S363(0) <='1';
          else
          oVar1S363(0) <='0';
          end if;
        if(cVar2S8S64P009N012P064nsss(0)='1'  OR cVar2S9S64P009P034nsss(0)='1'  OR cVar2S10S64P011P014nsss(0)='1'  OR cVar2S11S64P036P009nsss(0)='1'  )then
          oVar1S364(0) <='1';
          else
          oVar1S364(0) <='0';
          end if;
        if(cVar2S12S64P064P016nsss(0)='1'  OR cVar2S13S64P064P016P017nsss(0)='1'  OR cVar2S14S64N064P062P006nsss(0)='1'  OR cVar2S15S64N064P062P013nsss(0)='1'  )then
          oVar1S365(0) <='1';
          else
          oVar1S365(0) <='0';
          end if;
        if(cVar2S16S64P048P019nsss(0)='1'  OR cVar2S17S64N048P029nsss(0)='1'  OR cVar2S18S64N048N029P009nsss(0)='1'  OR cVar1S19S64P018P034P039P068nsss(0)='1'  )then
          oVar1S366(0) <='1';
          else
          oVar1S366(0) <='0';
          end if;
        if(cVar2S20S64P055P009P013nsss(0)='1'  OR cVar2S21S64P055N009P037nsss(0)='1'  OR cVar2S22S64P065P012P036nsss(0)='1'  )then
          oVar1S367(0) <='1';
          else
          oVar1S367(0) <='0';
          end if;
        if(cVar2S0S65P065P006P016nsss(0)='1'  OR cVar2S1S65N065P036P062nsss(0)='1'  OR cVar2S2S65N065P036P064nsss(0)='1'  OR cVar2S3S65P016P041nsss(0)='1'  )then
          oVar1S368(0) <='1';
          else
          oVar1S368(0) <='0';
          end if;
        if(cVar2S4S65P016N041P014nsss(0)='1'  OR cVar2S5S65P019nsss(0)='1'  OR cVar2S6S65P029nsss(0)='1'  OR cVar2S7S65N029P005P009nsss(0)='1'  )then
          oVar1S369(0) <='1';
          else
          oVar1S369(0) <='0';
          end if;
        if(cVar2S8S65P055P060P012nsss(0)='1'  OR cVar2S9S65P065P012P015nsss(0)='1'  OR cVar2S10S65P057nsss(0)='1'  OR cVar2S11S65N057P052nsss(0)='1'  )then
          oVar1S370(0) <='1';
          else
          oVar1S370(0) <='0';
          end if;
        if(cVar2S12S65N057N052P051nsss(0)='1'  OR cVar2S13S65P006P067nsss(0)='1'  OR cVar2S14S65P020nsss(0)='1'  OR cVar2S15S65N020P012nsss(0)='1'  )then
          oVar1S371(0) <='1';
          else
          oVar1S371(0) <='0';
          end if;
        if(cVar2S16S65P036P008P013nsss(0)='1'  OR cVar2S17S65P020P033P016nsss(0)='1'  OR cVar2S18S65P020P040nsss(0)='1'  OR cVar2S19S65P020N040P007nsss(0)='1'  )then
          oVar1S372(0) <='1';
          else
          oVar1S372(0) <='0';
          end if;
        if(cVar2S20S65P010P012P016nsss(0)='1'  )then
          oVar1S373(0) <='1';
          else
          oVar1S373(0) <='0';
          end if;
        if(cVar1S0S66P016P000P002P040nsss(0)='1'  OR cVar2S1S66P041nsss(0)='1'  OR cVar2S2S66N041P032nsss(0)='1'  OR cVar2S3S66P032P014nsss(0)='1'  )then
          oVar1S374(0) <='1';
          else
          oVar1S374(0) <='0';
          end if;
        if(cVar2S4S66P032N014P013nsss(0)='1'  OR cVar2S5S66N032P014nsss(0)='1'  OR cVar2S6S66P014P032nsss(0)='1'  OR cVar2S7S66P027P034P066nsss(0)='1'  )then
          oVar1S375(0) <='1';
          else
          oVar1S375(0) <='0';
          end if;
        if(cVar2S8S66P043P063P065nsss(0)='1'  OR cVar2S9S66P069P010P015nsss(0)='1'  OR cVar2S10S66P011nsss(0)='1'  OR cVar1S11S66P016P039P007P005nsss(0)='1'  )then
          oVar1S376(0) <='1';
          else
          oVar1S376(0) <='0';
          end if;
        if(cVar2S12S66P069P051nsss(0)='1'  )then
          oVar1S377(0) <='1';
          else
          oVar1S377(0) <='0';
          end if;
        if(cVar2S0S67P037P039P057nsss(0)='1'  OR cVar2S1S67N037P069P035nsss(0)='1'  OR cVar2S2S67N037P069P032nsss(0)='1'  OR cVar2S3S67P065P017P018nsss(0)='1'  )then
          oVar1S378(0) <='1';
          else
          oVar1S378(0) <='0';
          end if;
        if(cVar1S4S67P014P024P027P009nsss(0)='1'  OR cVar1S5S67P014P024P031P043nsss(0)='1'  OR cVar1S6S67N014P027P009P050nsss(0)='1'  OR cVar2S7S67P017nsss(0)='1'  )then
          oVar1S379(0) <='1';
          else
          oVar1S379(0) <='0';
          end if;
        if(cVar2S8S67P053P011nsss(0)='1'  OR cVar2S9S67P047nsss(0)='1'  OR cVar2S10S67N047P043nsss(0)='1'  OR cVar2S11S67P047P048P025nsss(0)='1'  )then
          oVar1S380(0) <='1';
          else
          oVar1S380(0) <='0';
          end if;
        if(cVar2S12S67P047P026nsss(0)='1'  OR cVar2S13S67P008P026nsss(0)='1'  OR cVar2S14S67P008N026P017nsss(0)='1'  OR cVar2S15S67N008P010P052nsss(0)='1'  )then
          oVar1S381(0) <='1';
          else
          oVar1S381(0) <='0';
          end if;
        if(cVar2S0S68P055P065P034nsss(0)='1'  OR cVar2S1S68P055N065P069nsss(0)='1'  OR cVar2S2S68N055P057P047nsss(0)='1'  OR cVar2S3S68P048nsss(0)='1'  )then
          oVar1S383(0) <='1';
          else
          oVar1S383(0) <='0';
          end if;
        if(cVar1S4S68P006P024P049P026nsss(0)='1'  OR cVar2S5S68P027nsss(0)='1'  OR cVar2S6S68N027P046nsss(0)='1'  OR cVar1S7S68P006P024P010P047nsss(0)='1'  )then
          oVar1S384(0) <='1';
          else
          oVar1S384(0) <='0';
          end if;
        if(cVar2S8S68P000nsss(0)='1'  OR cVar2S9S68N000P051P004nsss(0)='1'  OR cVar2S10S68P036P066nsss(0)='1'  OR cVar2S11S68P047nsss(0)='1'  )then
          oVar1S385(0) <='1';
          else
          oVar1S385(0) <='0';
          end if;
        if(cVar2S12S68N047P013P015nsss(0)='1'  OR cVar2S13S68P005P000P002nsss(0)='1'  OR cVar2S14S68P005P010nsss(0)='1'  OR cVar2S15S68P036P011P015nsss(0)='1'  )then
          oVar1S386(0) <='1';
          else
          oVar1S386(0) <='0';
          end if;
        if(cVar2S16S68P014P067nsss(0)='1'  )then
          oVar1S387(0) <='1';
          else
          oVar1S387(0) <='0';
          end if;
        if(cVar2S0S69P012nsss(0)='1'  OR cVar2S1S69P012P014nsss(0)='1'  OR cVar2S2S69P012nsss(0)='1'  OR cVar1S3S69P055P026N010P065nsss(0)='1'  )then
          oVar1S388(0) <='1';
          else
          oVar1S388(0) <='0';
          end if;
        if(cVar2S4S69P006P069P057nsss(0)='1'  OR cVar2S5S69P006N069P011nsss(0)='1'  OR cVar2S6S69P008nsss(0)='1'  OR cVar2S7S69N008P056nsss(0)='1'  )then
          oVar1S389(0) <='1';
          else
          oVar1S389(0) <='0';
          end if;
        if(cVar2S8S69P024P010nsss(0)='1'  OR cVar2S9S69N024P047P027nsss(0)='1'  OR cVar1S10S69N055P030P063P002nsss(0)='1'  OR cVar2S11S69P056P012nsss(0)='1'  )then
          oVar1S390(0) <='1';
          else
          oVar1S390(0) <='0';
          end if;
        if(cVar2S12S69N056P059P012nsss(0)='1'  OR cVar2S13S69N056N059P035nsss(0)='1'  OR cVar2S14S69P018nsss(0)='1'  )then
          oVar1S391(0) <='1';
          else
          oVar1S391(0) <='0';
          end if;
        if(cVar2S0S70P046P021P040nsss(0)='1'  OR cVar2S1S70P046N021P040nsss(0)='1'  OR cVar2S2S70P046P018P019nsss(0)='1'  OR cVar2S3S70P045nsss(0)='1'  )then
          oVar1S392(0) <='1';
          else
          oVar1S392(0) <='0';
          end if;
        if(cVar2S4S70N045P024nsss(0)='1'  OR cVar2S5S70N045N024P007nsss(0)='1'  OR cVar1S6S70P050P027P048P025nsss(0)='1'  OR cVar2S7S70P047nsss(0)='1'  )then
          oVar1S393(0) <='1';
          else
          oVar1S393(0) <='0';
          end if;
        if(cVar2S8S70N047P012P036nsss(0)='1'  OR cVar2S9S70N047N012P069nsss(0)='1'  OR cVar2S10S70P032P003nsss(0)='1'  OR cVar2S11S70P032N003P051nsss(0)='1'  )then
          oVar1S394(0) <='1';
          else
          oVar1S394(0) <='0';
          end if;
        if(cVar1S12S70P050P043P027P009nsss(0)='1'  OR cVar2S13S70P052nsss(0)='1'  OR cVar2S14S70P031nsss(0)='1'  OR cVar2S15S70N031P052P010nsss(0)='1'  )then
          oVar1S395(0) <='1';
          else
          oVar1S395(0) <='0';
          end if;
        if(cVar1S0S71P021P040nsss(0)='1'  OR cVar1S1S71P021N040P048P039nsss(0)='1'  OR cVar2S2S71P060P064nsss(0)='1'  OR cVar2S3S71P030P006nsss(0)='1'  )then
          oVar1S397(0) <='1';
          else
          oVar1S397(0) <='0';
          end if;
        if(cVar2S4S71N030P041P031nsss(0)='1'  OR cVar2S5S71P030P016P002nsss(0)='1'  OR cVar2S6S71P030N016P032nsss(0)='1'  OR cVar2S7S71P030P055P054nsss(0)='1'  )then
          oVar1S398(0) <='1';
          else
          oVar1S398(0) <='0';
          end if;
        if(cVar2S8S71P002nsss(0)='1'  OR cVar2S9S71N002P018P015nsss(0)='1'  OR cVar2S10S71N002N018P037nsss(0)='1'  OR cVar1S11S71N021P038P040P015nsss(0)='1'  )then
          oVar1S399(0) <='1';
          else
          oVar1S399(0) <='0';
          end if;
        if(cVar2S12S71P018nsss(0)='1'  OR cVar1S13S71N021P038N040P010nsss(0)='1'  )then
          oVar1S400(0) <='1';
          else
          oVar1S400(0) <='0';
          end if;
        if(cVar1S0S72P016P021P038nsss(0)='1'  OR cVar2S1S72P019P013P017nsss(0)='1'  OR cVar2S2S72N019P010P068nsss(0)='1'  OR cVar2S3S72P044P023nsss(0)='1'  )then
          oVar1S401(0) <='1';
          else
          oVar1S401(0) <='0';
          end if;
        if(cVar2S4S72P044N023P013nsss(0)='1'  OR cVar2S5S72N044P042P005nsss(0)='1'  OR cVar2S6S72P010nsss(0)='1'  OR cVar1S7S72P016N021P040P002nsss(0)='1'  )then
          oVar1S402(0) <='1';
          else
          oVar1S402(0) <='0';
          end if;
        if(cVar2S8S72P065P069nsss(0)='1'  OR cVar2S9S72P043P037P006nsss(0)='1'  OR cVar2S10S72P043P065P019nsss(0)='1'  OR cVar2S11S72P019P011nsss(0)='1'  )then
          oVar1S403(0) <='1';
          else
          oVar1S403(0) <='0';
          end if;
        if(cVar2S12S72P010P015nsss(0)='1'  OR cVar1S13S72P016P039P054P005nsss(0)='1'  OR cVar2S14S72P061nsss(0)='1'  )then
          oVar1S404(0) <='1';
          else
          oVar1S404(0) <='0';
          end if;
        if(cVar1S0S73P021P040nsss(0)='1'  OR cVar2S1S73P011P020nsss(0)='1'  OR cVar2S2S73P011P013P016nsss(0)='1'  OR cVar2S3S73P041P030P014nsss(0)='1'  )then
          oVar1S405(0) <='1';
          else
          oVar1S405(0) <='0';
          end if;
        if(cVar2S4S73P041N030P031nsss(0)='1'  OR cVar2S5S73P030P051P028nsss(0)='1'  OR cVar2S6S73P030P055P054nsss(0)='1'  OR cVar2S7S73P002nsss(0)='1'  )then
          oVar1S406(0) <='1';
          else
          oVar1S406(0) <='0';
          end if;
        if(cVar2S8S73N002P018P012nsss(0)='1'  OR cVar2S9S73N002N018P037nsss(0)='1'  OR cVar1S10S73N021P038P020nsss(0)='1'  OR cVar2S11S73P012P016nsss(0)='1'  )then
          oVar1S407(0) <='1';
          else
          oVar1S407(0) <='0';
          end if;
        if(cVar2S12S73N012P018P019nsss(0)='1'  )then
          oVar1S408(0) <='1';
          else
          oVar1S408(0) <='0';
          end if;
        if(cVar1S0S74P014P027P002P009nsss(0)='1'  OR cVar2S1S74P010P008nsss(0)='1'  OR cVar2S2S74P010N008P012nsss(0)='1'  OR cVar2S3S74P066nsss(0)='1'  )then
          oVar1S409(0) <='1';
          else
          oVar1S409(0) <='0';
          end if;
        if(cVar2S4S74P066P037nsss(0)='1'  OR cVar2S5S74P013P039P053nsss(0)='1'  OR cVar2S6S74N013P032P031nsss(0)='1'  OR cVar2S7S74P047nsss(0)='1'  )then
          oVar1S410(0) <='1';
          else
          oVar1S410(0) <='0';
          end if;
        if(cVar2S8S74N047P054nsss(0)='1'  OR cVar2S9S74P047P048P025nsss(0)='1'  OR cVar2S10S74P047P048P025nsss(0)='1'  OR cVar2S11S74P047P026nsss(0)='1'  )then
          oVar1S411(0) <='1';
          else
          oVar1S411(0) <='0';
          end if;
        if(cVar2S12S74P047N026P011nsss(0)='1'  OR cVar2S13S74P030P048nsss(0)='1'  OR cVar2S14S74P048P062nsss(0)='1'  OR cVar2S15S74P048N062P017nsss(0)='1'  )then
          oVar1S412(0) <='1';
          else
          oVar1S412(0) <='0';
          end if;
        if(cVar2S16S74N048P027P021nsss(0)='1'  OR cVar2S17S74P018P017nsss(0)='1'  OR cVar1S18S74P014P024P031P045nsss(0)='1'  OR cVar2S19S74P012P003P064nsss(0)='1'  )then
          oVar1S413(0) <='1';
          else
          oVar1S413(0) <='0';
          end if;
        if(cVar2S20S74P012P000nsss(0)='1'  )then
          oVar1S414(0) <='1';
          else
          oVar1S414(0) <='0';
          end if;
        if(cVar2S0S75P034nsss(0)='1'  OR cVar2S1S75P031P014nsss(0)='1'  OR cVar2S2S75N031P029nsss(0)='1'  OR cVar2S3S75N031N029P058nsss(0)='1'  )then
          oVar1S415(0) <='1';
          else
          oVar1S415(0) <='0';
          end if;
        if(cVar2S4S75P018nsss(0)='1'  OR cVar2S5S75P036P034nsss(0)='1'  OR cVar2S6S75P036N034P017nsss(0)='1'  OR cVar2S7S75P060P034nsss(0)='1'  )then
          oVar1S416(0) <='1';
          else
          oVar1S416(0) <='0';
          end if;
        if(cVar2S8S75P060N034P036nsss(0)='1'  OR cVar2S9S75N060P031P058nsss(0)='1'  OR cVar2S10S75N060P031P067nsss(0)='1'  OR cVar2S11S75P013P031nsss(0)='1'  )then
          oVar1S417(0) <='1';
          else
          oVar1S417(0) <='0';
          end if;
        if(cVar2S12S75N013P012P019nsss(0)='1'  OR cVar2S13S75P068P026P067nsss(0)='1'  OR cVar1S14S75N010N014P027P050nsss(0)='1'  OR cVar2S15S75P046nsss(0)='1'  )then
          oVar1S418(0) <='1';
          else
          oVar1S418(0) <='0';
          end if;
        if(cVar2S16S75N046P049nsss(0)='1'  OR cVar2S17S75N046N049P069nsss(0)='1'  OR cVar2S18S75P047nsss(0)='1'  OR cVar2S19S75N047P054P043nsss(0)='1'  )then
          oVar1S419(0) <='1';
          else
          oVar1S419(0) <='0';
          end if;
        if(cVar2S20S75P047P044P023nsss(0)='1'  OR cVar2S21S75P047N044P041nsss(0)='1'  OR cVar2S22S75P047P026nsss(0)='1'  )then
          oVar1S420(0) <='1';
          else
          oVar1S420(0) <='0';
          end if;
        if(cVar2S0S76P028nsss(0)='1'  OR cVar2S1S76N028P024nsss(0)='1'  OR cVar2S2S76P013nsss(0)='1'  OR cVar1S3S76P014N010P027P050nsss(0)='1'  )then
          oVar1S421(0) <='1';
          else
          oVar1S421(0) <='0';
          end if;
        if(cVar2S4S76P046nsss(0)='1'  OR cVar2S5S76N046P049nsss(0)='1'  OR cVar2S6S76P052P024nsss(0)='1'  OR cVar2S7S76P052N024P047nsss(0)='1'  )then
          oVar1S422(0) <='1';
          else
          oVar1S422(0) <='0';
          end if;
        if(cVar2S8S76P052P062nsss(0)='1'  OR cVar2S9S76P052N062P068nsss(0)='1'  OR cVar2S10S76P004P008P026nsss(0)='1'  OR cVar2S11S76P004N008P058nsss(0)='1'  )then
          oVar1S423(0) <='1';
          else
          oVar1S423(0) <='0';
          end if;
        if(cVar2S12S76P043P022P067nsss(0)='1'  OR cVar2S13S76P043P036P066nsss(0)='1'  OR cVar2S14S76P036nsss(0)='1'  OR cVar2S15S76N036P019P018nsss(0)='1'  )then
          oVar1S424(0) <='1';
          else
          oVar1S424(0) <='0';
          end if;
        if(cVar2S16S76P017P019nsss(0)='1'  OR cVar1S17S76P014P024P031P045nsss(0)='1'  OR cVar2S18S76P012P003P049nsss(0)='1'  OR cVar2S19S76P012P000nsss(0)='1'  )then
          oVar1S425(0) <='1';
          else
          oVar1S425(0) <='0';
          end if;
        if(cVar2S0S77P057nsss(0)='1'  OR cVar2S1S77N057P053nsss(0)='1'  OR cVar2S2S77N057N053P013nsss(0)='1'  OR cVar2S3S77P031nsss(0)='1'  )then
          oVar1S427(0) <='1';
          else
          oVar1S427(0) <='0';
          end if;
        if(cVar2S4S77N031P025nsss(0)='1'  OR cVar2S5S77P018nsss(0)='1'  OR cVar2S6S77P036P034nsss(0)='1'  OR cVar2S7S77P036N034P017nsss(0)='1'  )then
          oVar1S428(0) <='1';
          else
          oVar1S428(0) <='0';
          end if;
        if(cVar1S8S77N010P025P046nsss(0)='1'  OR cVar1S9S77N010P025N046P007nsss(0)='1'  OR cVar2S10S77P024nsss(0)='1'  OR cVar2S11S77N024P017P014nsss(0)='1'  )then
          oVar1S429(0) <='1';
          else
          oVar1S429(0) <='0';
          end if;
        if(cVar2S12S77P040nsss(0)='1'  OR cVar2S13S77N040P011nsss(0)='1'  OR cVar2S14S77N040P011P006nsss(0)='1'  OR cVar2S15S77P020P039nsss(0)='1'  )then
          oVar1S430(0) <='1';
          else
          oVar1S430(0) <='0';
          end if;
        if(cVar1S16S77N010N025P046P047nsss(0)='1'  OR cVar2S17S77P067P018nsss(0)='1'  OR cVar2S18S77N067P009nsss(0)='1'  OR cVar2S19S77N067N009P008nsss(0)='1'  )then
          oVar1S431(0) <='1';
          else
          oVar1S431(0) <='0';
          end if;
        if(cVar2S0S78P043P021nsss(0)='1'  OR cVar2S1S78P021P040nsss(0)='1'  OR cVar2S2S78P021N040P006nsss(0)='1'  OR cVar2S3S78N021P038P040nsss(0)='1'  )then
          oVar1S433(0) <='1';
          else
          oVar1S433(0) <='0';
          end if;
        if(cVar1S4S78P039P041P020P040nsss(0)='1'  OR cVar2S5S78P022P064P007nsss(0)='1'  OR cVar2S6S78P022P064P014nsss(0)='1'  OR cVar1S7S78P039P041P033nsss(0)='1'  )then
          oVar1S434(0) <='1';
          else
          oVar1S434(0) <='0';
          end if;
        if(cVar1S8S78P039P020P041nsss(0)='1'  OR cVar2S9S78P021nsss(0)='1'  OR cVar2S10S78N021P008P009nsss(0)='1'  )then
          oVar1S435(0) <='1';
          else
          oVar1S435(0) <='0';
          end if;
        if(cVar1S0S79P021P040nsss(0)='1'  OR cVar2S1S79P057P020nsss(0)='1'  OR cVar2S2S79P043P048nsss(0)='1'  OR cVar2S3S79P043N048P052nsss(0)='1'  )then
          oVar1S436(0) <='1';
          else
          oVar1S436(0) <='0';
          end if;
        if(cVar2S4S79P047P024P016nsss(0)='1'  OR cVar2S5S79P047N024P056nsss(0)='1'  OR cVar2S6S79N047P049P058nsss(0)='1'  OR cVar2S7S79N047P049P018nsss(0)='1'  )then
          oVar1S437(0) <='1';
          else
          oVar1S437(0) <='0';
          end if;
        if(cVar2S8S79P018P042nsss(0)='1'  OR cVar2S9S79P018N042P015nsss(0)='1'  OR cVar2S10S79N018P037nsss(0)='1'  OR cVar1S11S79N021P038P065P020nsss(0)='1'  )then
          oVar1S438(0) <='1';
          else
          oVar1S438(0) <='0';
          end if;
        if(cVar2S12S79P036P018P015nsss(0)='1'  OR cVar2S13S79P036N018P012nsss(0)='1'  )then
          oVar1S439(0) <='1';
          else
          oVar1S439(0) <='0';
          end if;
        if(cVar1S0S80P037P048P025nsss(0)='1'  OR cVar1S1S80P037P048N025P027nsss(0)='1'  OR cVar2S2S80P062P019nsss(0)='1'  OR cVar2S3S80N062P047nsss(0)='1'  )then
          oVar1S440(0) <='1';
          else
          oVar1S440(0) <='0';
          end if;
        if(cVar2S4S80N062N047P018nsss(0)='1'  OR cVar2S5S80P019P067P065nsss(0)='1'  OR cVar2S6S80N019P057P053nsss(0)='1'  OR cVar2S7S80N019N057P031nsss(0)='1'  )then
          oVar1S441(0) <='1';
          else
          oVar1S441(0) <='0';
          end if;
        if(cVar2S8S80P017P067P065nsss(0)='1'  OR cVar2S9S80P017N067P066nsss(0)='1'  OR cVar2S10S80P017P035P063nsss(0)='1'  OR cVar2S11S80P044P017nsss(0)='1'  )then
          oVar1S442(0) <='1';
          else
          oVar1S442(0) <='0';
          end if;
        if(cVar2S12S80N044P017nsss(0)='1'  OR cVar2S13S80P003P058nsss(0)='1'  OR cVar2S14S80P003P058P060nsss(0)='1'  OR cVar2S15S80P041nsss(0)='1'  )then
          oVar1S443(0) <='1';
          else
          oVar1S443(0) <='0';
          end if;
        if(cVar2S16S80N041P039P008nsss(0)='1'  OR cVar2S17S80P046nsss(0)='1'  OR cVar2S18S80P014nsss(0)='1'  OR cVar2S19S80N014P019nsss(0)='1'  )then
          oVar1S444(0) <='1';
          else
          oVar1S444(0) <='0';
          end if;
        if(cVar2S20S80P014P008P017nsss(0)='1'  OR cVar2S21S80P014P019P069nsss(0)='1'  OR cVar1S22S80P037P013N018P031nsss(0)='1'  OR cVar2S23S80P012P051P010nsss(0)='1'  )then
          oVar1S445(0) <='1';
          else
          oVar1S445(0) <='0';
          end if;
        if(cVar2S24S80N012P069P008nsss(0)='1'  )then
          oVar1S446(0) <='1';
          else
          oVar1S446(0) <='0';
          end if;
        if(cVar2S0S81P061nsss(0)='1'  OR cVar2S1S81P053P014nsss(0)='1'  OR cVar2S2S81P053N014P012nsss(0)='1'  OR cVar2S3S81N053P035nsss(0)='1'  )then
          oVar1S447(0) <='1';
          else
          oVar1S447(0) <='0';
          end if;
        if(cVar2S4S81N053N035P015nsss(0)='1'  OR cVar2S5S81P016P059nsss(0)='1'  OR cVar2S6S81P063P056P065nsss(0)='1'  OR cVar2S7S81P063P056P066nsss(0)='1'  )then
          oVar1S448(0) <='1';
          else
          oVar1S448(0) <='0';
          end if;
        if(cVar2S8S81P063P024P003nsss(0)='1'  OR cVar2S9S81P012P018nsss(0)='1'  OR cVar2S10S81P036nsss(0)='1'  OR cVar2S11S81N036P018nsss(0)='1'  )then
          oVar1S449(0) <='1';
          else
          oVar1S449(0) <='0';
          end if;
        if(cVar2S12S81P062P063P018nsss(0)='1'  OR cVar2S13S81P031nsss(0)='1'  OR cVar2S14S81N031P013P060nsss(0)='1'  OR cVar2S15S81N031P013P067nsss(0)='1'  )then
          oVar1S450(0) <='1';
          else
          oVar1S450(0) <='0';
          end if;
        if(cVar2S16S81P005P067P066nsss(0)='1'  OR cVar2S17S81P005P067P062nsss(0)='1'  OR cVar1S18S81N019P037P003P034nsss(0)='1'  OR cVar2S19S81P036N016P013nsss(0)='1'  )then
          oVar1S451(0) <='1';
          else
          oVar1S451(0) <='0';
          end if;
        if(cVar1S20S81N019N037P048P062nsss(0)='1'  OR cVar2S21S81P027nsss(0)='1'  OR cVar2S22S81N027P025nsss(0)='1'  OR cVar2S23S81N027N025P054nsss(0)='1'  )then
          oVar1S452(0) <='1';
          else
          oVar1S452(0) <='0';
          end if;
        if(cVar2S24S81P013P012nsss(0)='1'  OR cVar2S25S81N013P011nsss(0)='1'  OR cVar2S26S81N013N011P015nsss(0)='1'  OR cVar2S27S81P015P004P035nsss(0)='1'  )then
          oVar1S453(0) <='1';
          else
          oVar1S453(0) <='0';
          end if;
        if(cVar2S28S81P015P004P013nsss(0)='1'  OR cVar2S29S81N015P051P011nsss(0)='1'  )then
          oVar1S454(0) <='1';
          else
          oVar1S454(0) <='0';
          end if;
        if(cVar1S0S82P019P030P040P021nsss(0)='1'  OR cVar2S1S82P002nsss(0)='1'  OR cVar2S2S82N002P066P018nsss(0)='1'  OR cVar2S3S82P021P050nsss(0)='1'  )then
          oVar1S455(0) <='1';
          else
          oVar1S455(0) <='0';
          end if;
        if(cVar2S4S82P021N050P055nsss(0)='1'  OR cVar2S5S82P021P006nsss(0)='1'  OR cVar1S6S82P019P030P045P056nsss(0)='1'  OR cVar2S7S82P002nsss(0)='1'  )then
          oVar1S456(0) <='1';
          else
          oVar1S456(0) <='0';
          end if;
        if(cVar2S8S82N002P057P014nsss(0)='1'  OR cVar2S9S82N002N057P007nsss(0)='1'  OR cVar1S10S82P019P017P055P065nsss(0)='1'  OR cVar2S11S82P059P053nsss(0)='1'  )then
          oVar1S457(0) <='1';
          else
          oVar1S457(0) <='0';
          end if;
        if(cVar2S12S82P053P014nsss(0)='1'  OR cVar2S13S82P053N014P016nsss(0)='1'  OR cVar2S14S82N053P061nsss(0)='1'  OR cVar2S15S82P016P059nsss(0)='1'  )then
          oVar1S458(0) <='1';
          else
          oVar1S458(0) <='0';
          end if;
        if(cVar2S16S82P031P008nsss(0)='1'  OR cVar2S17S82N031P024P016nsss(0)='1'  OR cVar2S18S82P014nsss(0)='1'  OR cVar2S19S82P008nsss(0)='1'  )then
          oVar1S459(0) <='1';
          else
          oVar1S459(0) <='0';
          end if;
        if(cVar2S0S83P003P034P024nsss(0)='1'  OR cVar2S1S83P003P018P016nsss(0)='1'  OR cVar2S2S83P061P033nsss(0)='1'  OR cVar2S3S83P061N033P018nsss(0)='1'  )then
          oVar1S461(0) <='1';
          else
          oVar1S461(0) <='0';
          end if;
        if(cVar2S4S83N061P032P011nsss(0)='1'  OR cVar2S5S83N061N032P034nsss(0)='1'  OR cVar2S6S83P033P009P065nsss(0)='1'  OR cVar2S7S83P033P037P068nsss(0)='1'  )then
          oVar1S462(0) <='1';
          else
          oVar1S462(0) <='0';
          end if;
        if(cVar2S8S83P060nsss(0)='1'  OR cVar2S9S83P036nsss(0)='1'  OR cVar2S10S83N036P069P011nsss(0)='1'  OR cVar2S11S83P035nsss(0)='1'  )then
          oVar1S463(0) <='1';
          else
          oVar1S463(0) <='0';
          end if;
        if(cVar1S12S83N015P021P038nsss(0)='1'  OR cVar2S13S83P013P012nsss(0)='1'  OR cVar2S14S83P013N012P019nsss(0)='1'  OR cVar2S15S83P026P035nsss(0)='1'  )then
          oVar1S464(0) <='1';
          else
          oVar1S464(0) <='0';
          end if;
        if(cVar2S16S83P026P035P014nsss(0)='1'  OR cVar2S17S83P026P068P018nsss(0)='1'  OR cVar2S18S83P051P011P066nsss(0)='1'  OR cVar2S19S83P051N011P008nsss(0)='1'  )then
          oVar1S465(0) <='1';
          else
          oVar1S465(0) <='0';
          end if;
        if(cVar2S20S83N051P053P047nsss(0)='1'  OR cVar2S21S83P014P012nsss(0)='1'  OR cVar2S22S83P014N012P040nsss(0)='1'  )then
          oVar1S466(0) <='1';
          else
          oVar1S466(0) <='0';
          end if;
        if(cVar1S0S84P067P037P021P040nsss(0)='1'  OR cVar2S1S84P064nsss(0)='1'  OR cVar2S2S84N064P011P066nsss(0)='1'  OR cVar2S3S84P031P011nsss(0)='1'  )then
          oVar1S467(0) <='1';
          else
          oVar1S467(0) <='0';
          end if;
        if(cVar2S4S84N031P029P015nsss(0)='1'  OR cVar2S5S84N031N029P056nsss(0)='1'  OR cVar2S6S84P031P032P058nsss(0)='1'  OR cVar2S7S84P031P032P059nsss(0)='1'  )then
          oVar1S468(0) <='1';
          else
          oVar1S468(0) <='0';
          end if;
        if(cVar2S8S84P031P012P014nsss(0)='1'  OR cVar1S9S84P067P037P028nsss(0)='1'  OR cVar2S10S84P048P000P017nsss(0)='1'  OR cVar2S11S84P048N000P051nsss(0)='1'  )then
          oVar1S469(0) <='1';
          else
          oVar1S469(0) <='0';
          end if;
        if(cVar2S12S84P048P046nsss(0)='1'  OR cVar2S13S84P018P004P009nsss(0)='1'  OR cVar2S14S84N018P031nsss(0)='1'  OR cVar2S15S84P068P032nsss(0)='1'  )then
          oVar1S470(0) <='1';
          else
          oVar1S470(0) <='0';
          end if;
        if(cVar2S16S84P068P012nsss(0)='1'  OR cVar2S17S84P015P018nsss(0)='1'  OR cVar2S18S84P058P009P012nsss(0)='1'  OR cVar2S19S84P052P011nsss(0)='1'  )then
          oVar1S471(0) <='1';
          else
          oVar1S471(0) <='0';
          end if;
        if(cVar2S20S84N052P063P059nsss(0)='1'  OR cVar2S21S84N052P063P024nsss(0)='1'  OR cVar2S22S84P000P028nsss(0)='1'  )then
          oVar1S472(0) <='1';
          else
          oVar1S472(0) <='0';
          end if;
        if(cVar2S0S85P019P014nsss(0)='1'  OR cVar2S1S85N019P012nsss(0)='1'  OR cVar2S2S85P057P035P030nsss(0)='1'  OR cVar2S3S85P057P035P062nsss(0)='1'  )then
          oVar1S473(0) <='1';
          else
          oVar1S473(0) <='0';
          end if;
        if(cVar2S4S85P057P018nsss(0)='1'  OR cVar2S5S85P046nsss(0)='1'  OR cVar2S6S85P017P066nsss(0)='1'  OR cVar2S7S85P017N066P036nsss(0)='1'  )then
          oVar1S474(0) <='1';
          else
          oVar1S474(0) <='0';
          end if;
        if(cVar2S8S85P017P015P019nsss(0)='1'  OR cVar2S9S85P017P015P035nsss(0)='1'  OR cVar2S10S85P031nsss(0)='1'  OR cVar2S11S85N031P012P066nsss(0)='1'  )then
          oVar1S475(0) <='1';
          else
          oVar1S475(0) <='0';
          end if;
        if(cVar1S12S85N037P058P011P031nsss(0)='1'  OR cVar2S13S85P033P062nsss(0)='1'  OR cVar2S14S85P033N062P012nsss(0)='1'  OR cVar2S15S85N033P010P016nsss(0)='1'  )then
          oVar1S476(0) <='1';
          else
          oVar1S476(0) <='0';
          end if;
        if(cVar2S16S85N033N010P035nsss(0)='1'  OR cVar2S17S85P013P017nsss(0)='1'  OR cVar2S18S85P013N017P014nsss(0)='1'  OR cVar1S19S85N037N058P021P040nsss(0)='1'  )then
          oVar1S477(0) <='1';
          else
          oVar1S477(0) <='0';
          end if;
        if(cVar2S20S85P061P064nsss(0)='1'  OR cVar2S21S85P061N064P011nsss(0)='1'  OR cVar2S22S85P025nsss(0)='1'  OR cVar2S23S85N025P027nsss(0)='1'  )then
          oVar1S478(0) <='1';
          else
          oVar1S478(0) <='0';
          end if;
        if(cVar2S24S85N025N027P026nsss(0)='1'  OR cVar2S25S85P046P020P039nsss(0)='1'  )then
          oVar1S479(0) <='1';
          else
          oVar1S479(0) <='0';
          end if;
        if(cVar1S0S86P037P048P025nsss(0)='1'  OR cVar2S1S86P027nsss(0)='1'  OR cVar2S2S86N027P012nsss(0)='1'  OR cVar2S3S86P047nsss(0)='1'  )then
          oVar1S480(0) <='1';
          else
          oVar1S480(0) <='0';
          end if;
        if(cVar2S4S86N047P062nsss(0)='1'  OR cVar2S5S86P032P056nsss(0)='1'  OR cVar2S6S86P032N056P001nsss(0)='1'  OR cVar2S7S86P032P069P015nsss(0)='1'  )then
          oVar1S481(0) <='1';
          else
          oVar1S481(0) <='0';
          end if;
        if(cVar2S8S86P009P019P044nsss(0)='1'  OR cVar2S9S86P009N019psss(0)='1'  OR cVar2S10S86P009P016P019nsss(0)='1'  OR cVar2S11S86P019P018nsss(0)='1'  )then
          oVar1S482(0) <='1';
          else
          oVar1S482(0) <='0';
          end if;
        if(cVar2S12S86P019N018P044nsss(0)='1'  OR cVar2S13S86P014nsss(0)='1'  OR cVar2S14S86P019P014nsss(0)='1'  OR cVar2S15S86N019P057nsss(0)='1'  )then
          oVar1S483(0) <='1';
          else
          oVar1S483(0) <='0';
          end if;
        if(cVar2S16S86P057P014nsss(0)='1'  OR cVar2S17S86P057N014P051nsss(0)='1'  OR cVar2S18S86P066P017nsss(0)='1'  OR cVar2S19S86P066P062P017nsss(0)='1'  )then
          oVar1S484(0) <='1';
          else
          oVar1S484(0) <='0';
          end if;
        if(cVar2S0S87P016P064nsss(0)='1'  OR cVar2S1S87P016N064P036nsss(0)='1'  OR cVar2S2S87N016P011nsss(0)='1'  OR cVar2S3S87N016N011P014nsss(0)='1'  )then
          oVar1S486(0) <='1';
          else
          oVar1S486(0) <='0';
          end if;
        if(cVar2S4S87P036P010P009nsss(0)='1'  OR cVar2S5S87N036P067P034nsss(0)='1'  OR cVar2S6S87N036N067P060nsss(0)='1'  OR cVar2S7S87P033P045P014nsss(0)='1'  )then
          oVar1S487(0) <='1';
          else
          oVar1S487(0) <='0';
          end if;
        if(cVar2S8S87P033N045P043nsss(0)='1'  OR cVar2S9S87P033P012P015nsss(0)='1'  OR cVar2S10S87P035P031P015nsss(0)='1'  OR cVar2S11S87P035P032P063nsss(0)='1'  )then
          oVar1S488(0) <='1';
          else
          oVar1S488(0) <='0';
          end if;
        if(cVar2S12S87P011nsss(0)='1'  OR cVar2S13S87P014nsss(0)='1'  OR cVar2S14S87P034P035nsss(0)='1'  OR cVar2S15S87N034P006P011nsss(0)='1'  )then
          oVar1S489(0) <='1';
          else
          oVar1S489(0) <='0';
          end if;
        if(cVar2S16S87N034N006P027nsss(0)='1'  OR cVar1S17S87N019P009P068P053nsss(0)='1'  OR cVar1S18S87N019N009P040P021nsss(0)='1'  OR cVar2S19S87P020nsss(0)='1'  )then
          oVar1S490(0) <='1';
          else
          oVar1S490(0) <='0';
          end if;
        if(cVar2S20S87N020P017P018nsss(0)='1'  OR cVar2S21S87N020N017P018nsss(0)='1'  OR cVar2S22S87P021P068P047nsss(0)='1'  OR cVar2S23S87P021N068P060nsss(0)='1'  )then
          oVar1S491(0) <='1';
          else
          oVar1S491(0) <='0';
          end if;
        if(cVar2S24S87P021P039nsss(0)='1'  OR cVar2S25S87P015nsss(0)='1'  )then
          oVar1S492(0) <='1';
          else
          oVar1S492(0) <='0';
          end if;
        if(cVar2S0S88P007P005P013nsss(0)='1'  OR cVar2S1S88N007P012nsss(0)='1'  OR cVar2S2S88N007P012P013nsss(0)='1'  OR cVar2S3S88P008P016P012nsss(0)='1'  )then
          oVar1S493(0) <='1';
          else
          oVar1S493(0) <='0';
          end if;
        if(cVar2S4S88P008N016P036nsss(0)='1'  OR cVar2S5S88P059P018nsss(0)='1'  OR cVar2S6S88N059P066P062nsss(0)='1'  OR cVar2S7S88P007nsss(0)='1'  )then
          oVar1S494(0) <='1';
          else
          oVar1S494(0) <='0';
          end if;
        if(cVar2S8S88P058P028P052nsss(0)='1'  OR cVar2S9S88P058P028P054nsss(0)='1'  OR cVar2S10S88P058P037P052nsss(0)='1'  OR cVar1S11S88P060N009P053P028nsss(0)='1'  )then
          oVar1S495(0) <='1';
          else
          oVar1S495(0) <='0';
          end if;
        if(cVar2S12S88P008P026nsss(0)='1'  OR cVar2S13S88N008P029nsss(0)='1'  OR cVar2S14S88N008N029P048nsss(0)='1'  OR cVar2S15S88P034nsss(0)='1'  )then
          oVar1S496(0) <='1';
          else
          oVar1S496(0) <='0';
          end if;
        if(cVar2S16S88N034P009P016nsss(0)='1'  OR cVar2S17S88P012nsss(0)='1'  OR cVar2S18S88N012P013nsss(0)='1'  OR cVar2S19S88P069P014nsss(0)='1'  )then
          oVar1S497(0) <='1';
          else
          oVar1S497(0) <='0';
          end if;
        if(cVar2S20S88N069P065P066nsss(0)='1'  )then
          oVar1S498(0) <='1';
          else
          oVar1S498(0) <='0';
          end if;
        if(cVar2S0S89P005P013nsss(0)='1'  OR cVar2S1S89P005P013P019nsss(0)='1'  OR cVar2S2S89P030P012nsss(0)='1'  OR cVar2S3S89P066P016nsss(0)='1'  )then
          oVar1S499(0) <='1';
          else
          oVar1S499(0) <='0';
          end if;
        if(cVar1S4S89P009P068P002P047nsss(0)='1'  OR cVar2S5S89P059P017nsss(0)='1'  OR cVar2S6S89N059P066P050nsss(0)='1'  OR cVar1S7S89N009P049P023P005nsss(0)='1'  )then
          oVar1S500(0) <='1';
          else
          oVar1S500(0) <='0';
          end if;
        if(cVar2S8S89P042nsss(0)='1'  OR cVar2S9S89N042P007nsss(0)='1'  OR cVar2S10S89N042N007P036nsss(0)='1'  OR cVar2S11S89P022P045P012nsss(0)='1'  )then
          oVar1S501(0) <='1';
          else
          oVar1S501(0) <='0';
          end if;
        if(cVar2S12S89P022P014P042nsss(0)='1'  OR cVar2S13S89P022nsss(0)='1'  OR cVar2S14S89N022P024P045nsss(0)='1'  OR cVar2S15S89N022N024P007nsss(0)='1'  )then
          oVar1S502(0) <='1';
          else
          oVar1S502(0) <='0';
          end if;
        if(cVar1S16S89N009P049P026P014nsss(0)='1'  OR cVar2S17S89P047nsss(0)='1'  OR cVar2S18S89P046nsss(0)='1'  OR cVar2S19S89N046P005nsss(0)='1'  )then
          oVar1S503(0) <='1';
          else
          oVar1S503(0) <='0';
          end if;
        if(cVar2S20S89N046N005P007nsss(0)='1'  )then
          oVar1S504(0) <='1';
          else
          oVar1S504(0) <='0';
          end if;
        if(cVar1S0S90P049P052P065P069nsss(0)='1'  OR cVar2S1S90P035nsss(0)='1'  OR cVar2S2S90P050P018P016nsss(0)='1'  OR cVar2S3S90P050P018P029nsss(0)='1'  )then
          oVar1S505(0) <='1';
          else
          oVar1S505(0) <='0';
          end if;
        if(cVar2S4S90N050P066nsss(0)='1'  OR cVar2S5S90N050N066P013nsss(0)='1'  OR cVar2S6S90P026P010P057nsss(0)='1'  OR cVar2S7S90P026N010P006nsss(0)='1'  )then
          oVar1S506(0) <='1';
          else
          oVar1S506(0) <='0';
          end if;
        if(cVar2S8S90P043P022P045nsss(0)='1'  OR cVar2S9S90P043P022P002nsss(0)='1'  OR cVar2S10S90P043P022nsss(0)='1'  OR cVar2S11S90P043N022P023nsss(0)='1'  )then
          oVar1S507(0) <='1';
          else
          oVar1S507(0) <='0';
          end if;
        if(cVar2S12S90P019nsss(0)='1'  OR cVar2S13S90P051nsss(0)='1'  OR cVar1S14S90P049P026P063nsss(0)='1'  OR cVar1S15S90P049N026P027P009nsss(0)='1'  )then
          oVar1S508(0) <='1';
          else
          oVar1S508(0) <='0';
          end if;
        if(cVar2S16S90P047nsss(0)='1'  OR cVar2S17S90P046nsss(0)='1'  OR cVar2S18S90N046P016P051nsss(0)='1'  OR cVar2S19S90N046N016P005nsss(0)='1'  )then
          oVar1S509(0) <='1';
          else
          oVar1S509(0) <='0';
          end if;
        if(cVar1S0S91P052P065P069nsss(0)='1'  OR cVar1S1S91P052N065P062P035nsss(0)='1'  OR cVar2S2S91P034P016nsss(0)='1'  OR cVar2S3S91P034P016P015nsss(0)='1'  )then
          oVar1S511(0) <='1';
          else
          oVar1S511(0) <='0';
          end if;
        if(cVar2S4S91P067nsss(0)='1'  OR cVar2S5S91N067P066nsss(0)='1'  OR cVar2S6S91N067N066P013nsss(0)='1'  OR cVar2S7S91P025nsss(0)='1'  )then
          oVar1S512(0) <='1';
          else
          oVar1S512(0) <='0';
          end if;
        if(cVar2S8S91N025P018nsss(0)='1'  OR cVar2S9S91P037P062nsss(0)='1'  OR cVar2S10S91P037N062P067nsss(0)='1'  OR cVar2S11S91P037P018P066nsss(0)='1'  )then
          oVar1S513(0) <='1';
          else
          oVar1S513(0) <='0';
          end if;
        if(cVar1S12S91N052P048P061P014nsss(0)='1'  OR cVar2S13S91P026P004nsss(0)='1'  OR cVar2S14S91P057P040P021nsss(0)='1'  OR cVar2S15S91P065P001P016nsss(0)='1'  )then
          oVar1S514(0) <='1';
          else
          oVar1S514(0) <='0';
          end if;
        if(cVar1S0S92P019P068P029P054nsss(0)='1'  OR cVar2S1S92P051nsss(0)='1'  OR cVar2S2S92N051P052nsss(0)='1'  OR cVar2S3S92N051N052P015nsss(0)='1'  )then
          oVar1S516(0) <='1';
          else
          oVar1S516(0) <='0';
          end if;
        if(cVar2S4S92P037P007P003nsss(0)='1'  OR cVar2S5S92P037P007P009nsss(0)='1'  OR cVar2S6S92N037P045nsss(0)='1'  OR cVar2S7S92N037N045P043nsss(0)='1'  )then
          oVar1S517(0) <='1';
          else
          oVar1S517(0) <='0';
          end if;
        if(cVar2S8S92P034nsss(0)='1'  OR cVar2S9S92N034P026P030nsss(0)='1'  OR cVar2S10S92P010nsss(0)='1'  OR cVar2S11S92P011P029P056nsss(0)='1'  )then
          oVar1S518(0) <='1';
          else
          oVar1S518(0) <='0';
          end if;
        if(cVar1S12S92P019P068P055P010nsss(0)='1'  OR cVar1S13S92P019P066P009P046nsss(0)='1'  OR cVar2S14S92P050P061P059nsss(0)='1'  OR cVar2S15S92P050N061P048nsss(0)='1'  )then
          oVar1S519(0) <='1';
          else
          oVar1S519(0) <='0';
          end if;
        if(cVar2S16S92P050P052nsss(0)='1'  OR cVar2S17S92P004P006nsss(0)='1'  OR cVar2S18S92P004N006P013nsss(0)='1'  OR cVar2S19S92P015P011nsss(0)='1'  )then
          oVar1S520(0) <='1';
          else
          oVar1S520(0) <='0';
          end if;
        if(cVar2S20S92N015P028P018nsss(0)='1'  OR cVar2S21S92N015N028P048nsss(0)='1'  OR cVar2S22S92P058P015nsss(0)='1'  OR cVar2S23S92N058P067P015nsss(0)='1'  )then
          oVar1S521(0) <='1';
          else
          oVar1S521(0) <='0';
          end if;
        if(cVar2S24S92P036P063nsss(0)='1'  OR cVar2S25S92P036N063P008nsss(0)='1'  OR cVar2S26S92P013P065P014nsss(0)='1'  )then
          oVar1S522(0) <='1';
          else
          oVar1S522(0) <='0';
          end if;
        if(cVar2S0S93P012P036nsss(0)='1'  OR cVar2S1S93P012N036P069nsss(0)='1'  OR cVar2S2S93P012P010nsss(0)='1'  OR cVar2S3S93P069P065P059nsss(0)='1'  )then
          oVar1S523(0) <='1';
          else
          oVar1S523(0) <='0';
          end if;
        if(cVar2S4S93P069N065P030nsss(0)='1'  OR cVar2S5S93N069P047nsss(0)='1'  OR cVar2S6S93N069N047P036nsss(0)='1'  OR cVar2S7S93P036P010nsss(0)='1'  )then
          oVar1S524(0) <='1';
          else
          oVar1S524(0) <='0';
          end if;
        if(cVar2S8S93P067P014nsss(0)='1'  OR cVar2S9S93P008P013nsss(0)='1'  OR cVar2S10S93N008P017P013nsss(0)='1'  OR cVar1S11S93N019P056P054P013nsss(0)='1'  )then
          oVar1S525(0) <='1';
          else
          oVar1S525(0) <='0';
          end if;
        if(cVar2S12S93P016nsss(0)='1'  OR cVar2S13S93P012nsss(0)='1'  OR cVar2S14S93N012P060nsss(0)='1'  OR cVar2S15S93P037P017P015nsss(0)='1'  )then
          oVar1S526(0) <='1';
          else
          oVar1S526(0) <='0';
          end if;
        if(cVar2S16S93P029P028nsss(0)='1'  OR cVar2S17S93P029N028P003nsss(0)='1'  OR cVar2S18S93P007P025nsss(0)='1'  OR cVar2S19S93P007N025P002nsss(0)='1'  )then
          oVar1S527(0) <='1';
          else
          oVar1S527(0) <='0';
          end if;
        if(cVar2S20S93N007P053P009nsss(0)='1'  OR cVar2S21S93P034nsss(0)='1'  OR cVar2S22S93N034P063P036nsss(0)='1'  )then
          oVar1S528(0) <='1';
          else
          oVar1S528(0) <='0';
          end if;
        if(cVar2S0S94P054nsss(0)='1'  OR cVar2S1S94N054P051nsss(0)='1'  OR cVar2S2S94N054N051P052nsss(0)='1'  OR cVar2S3S94P034nsss(0)='1'  )then
          oVar1S529(0) <='1';
          else
          oVar1S529(0) <='0';
          end if;
        if(cVar2S4S94N034P015nsss(0)='1'  OR cVar2S5S94N034N015P052nsss(0)='1'  OR cVar2S6S94P005nsss(0)='1'  OR cVar2S7S94N005P024nsss(0)='1'  )then
          oVar1S530(0) <='1';
          else
          oVar1S530(0) <='0';
          end if;
        if(cVar2S8S94N005N024P007nsss(0)='1'  OR cVar2S9S94P022P043nsss(0)='1'  OR cVar2S10S94P022P043P008nsss(0)='1'  OR cVar1S11S94P019P037P059P028nsss(0)='1'  )then
          oVar1S531(0) <='1';
          else
          oVar1S531(0) <='0';
          end if;
        if(cVar2S12S94P055P008P057nsss(0)='1'  OR cVar2S13S94P017nsss(0)='1'  OR cVar2S14S94N017P061nsss(0)='1'  OR cVar2S15S94P042nsss(0)='1'  )then
          oVar1S532(0) <='1';
          else
          oVar1S532(0) <='0';
          end if;
        if(cVar2S16S94N042P002nsss(0)='1'  OR cVar2S17S94P053nsss(0)='1'  OR cVar2S18S94P008P063P066nsss(0)='1'  OR cVar2S19S94P008N063P032nsss(0)='1'  )then
          oVar1S533(0) <='1';
          else
          oVar1S533(0) <='0';
          end if;
        if(cVar2S20S94N008P018P061nsss(0)='1'  OR cVar2S21S94P018P030nsss(0)='1'  OR cVar2S22S94P018N030P036nsss(0)='1'  OR cVar2S23S94P018P068P055nsss(0)='1'  )then
          oVar1S534(0) <='1';
          else
          oVar1S534(0) <='0';
          end if;
        if(cVar2S0S95P066P012nsss(0)='1'  OR cVar2S1S95P066P012P069nsss(0)='1'  OR cVar2S2S95P066P014nsss(0)='1'  OR cVar2S3S95P032P004P016nsss(0)='1'  )then
          oVar1S536(0) <='1';
          else
          oVar1S536(0) <='0';
          end if;
        if(cVar2S4S95P032P012P014nsss(0)='1'  OR cVar2S5S95P009P004P012nsss(0)='1'  OR cVar2S6S95P009N004P044nsss(0)='1'  OR cVar2S7S95P009P017P063nsss(0)='1'  )then
          oVar1S537(0) <='1';
          else
          oVar1S537(0) <='0';
          end if;
        if(cVar2S8S95P007nsss(0)='1'  OR cVar2S9S95N007P010P015nsss(0)='1'  OR cVar1S10S95P019P057P030P056nsss(0)='1'  OR cVar2S11S95P017P068nsss(0)='1'  )then
          oVar1S538(0) <='1';
          else
          oVar1S538(0) <='0';
          end if;
        if(cVar2S12S95P060P014P037nsss(0)='1'  OR cVar1S13S95N019P045P062P005nsss(0)='1'  OR cVar2S14S95P007nsss(0)='1'  OR cVar2S15S95N007P069P024nsss(0)='1'  )then
          oVar1S539(0) <='1';
          else
          oVar1S539(0) <='0';
          end if;
        if(cVar2S16S95P054nsss(0)='1'  OR cVar2S17S95N054P051nsss(0)='1'  OR cVar2S18S95N054N051P052nsss(0)='1'  OR cVar2S19S95P055P008nsss(0)='1'  )then
          oVar1S540(0) <='1';
          else
          oVar1S540(0) <='0';
          end if;
        if(cVar2S20S95P055N008P015nsss(0)='1'  OR cVar2S21S95P013P011nsss(0)='1'  OR cVar2S22S95N013P016P012nsss(0)='1'  OR cVar2S23S95N013P016P012nsss(0)='1'  )then
          oVar1S541(0) <='1';
          else
          oVar1S541(0) <='0';
          end if;
        if(cVar2S24S95P054P002P026nsss(0)='1'  OR cVar2S25S95P054N002P028nsss(0)='1'  OR cVar2S26S95P054P030nsss(0)='1'  )then
          oVar1S542(0) <='1';
          else
          oVar1S542(0) <='0';
          end if;
        if(cVar1S0S96P019P037P045P005nsss(0)='1'  OR cVar2S1S96P069P024nsss(0)='1'  OR cVar2S2S96P069N024P011nsss(0)='1'  OR cVar2S3S96P011nsss(0)='1'  )then
          oVar1S543(0) <='1';
          else
          oVar1S543(0) <='0';
          end if;
        if(cVar2S4S96N011P034nsss(0)='1'  OR cVar2S5S96N011N034P015nsss(0)='1'  OR cVar2S6S96P040P038nsss(0)='1'  OR cVar2S7S96P040N038P042nsss(0)='1'  )then
          oVar1S544(0) <='1';
          else
          oVar1S544(0) <='0';
          end if;
        if(cVar2S8S96N040P038P022nsss(0)='1'  OR cVar1S9S96P019P037P059P028nsss(0)='1'  OR cVar2S10S96P049P064P018nsss(0)='1'  OR cVar2S11S96P049N064P041nsss(0)='1'  )then
          oVar1S545(0) <='1';
          else
          oVar1S545(0) <='0';
          end if;
        if(cVar2S12S96P017nsss(0)='1'  OR cVar2S13S96N017P061nsss(0)='1'  OR cVar2S14S96P060P034P012nsss(0)='1'  OR cVar2S15S96P051P056nsss(0)='1'  )then
          oVar1S546(0) <='1';
          else
          oVar1S546(0) <='0';
          end if;
        if(cVar2S16S96P051N056P011nsss(0)='1'  OR cVar2S17S96P051P012P016nsss(0)='1'  OR cVar2S18S96P034P037nsss(0)='1'  OR cVar2S19S96P034N037P013nsss(0)='1'  )then
          oVar1S547(0) <='1';
          else
          oVar1S547(0) <='0';
          end if;
        if(cVar2S20S96P064P012nsss(0)='1'  OR cVar2S21S96P064N012P068nsss(0)='1'  OR cVar2S22S96N064P061P062nsss(0)='1'  OR cVar2S23S96P065P031P004nsss(0)='1'  )then
          oVar1S548(0) <='1';
          else
          oVar1S548(0) <='0';
          end if;
        if(cVar2S24S96P065P031P058nsss(0)='1'  OR cVar2S25S96P065P034P066nsss(0)='1'  OR cVar2S26S96P020P039nsss(0)='1'  )then
          oVar1S549(0) <='1';
          else
          oVar1S549(0) <='0';
          end if;
        if(cVar1S0S97P045P035P025nsss(0)='1'  OR cVar1S1S97P045P035N025P022nsss(0)='1'  OR cVar2S2S97P023nsss(0)='1'  OR cVar2S3S97N023P024nsss(0)='1'  )then
          oVar1S550(0) <='1';
          else
          oVar1S550(0) <='0';
          end if;
        if(cVar2S4S97P004P030P031nsss(0)='1'  OR cVar2S5S97P004N030P057nsss(0)='1'  OR cVar2S6S97P012P017nsss(0)='1'  OR cVar2S7S97P029P011nsss(0)='1'  )then
          oVar1S551(0) <='1';
          else
          oVar1S551(0) <='0';
          end if;
        if(cVar2S8S97P029N011P008nsss(0)='1'  OR cVar2S9S97N029P037P025nsss(0)='1'  OR cVar2S10S97N029N037P040nsss(0)='1'  OR cVar2S11S97P014P035P006nsss(0)='1'  )then
          oVar1S552(0) <='1';
          else
          oVar1S552(0) <='0';
          end if;
        if(cVar1S12S97N045P043P022nsss(0)='1'  OR cVar1S13S97N045P043N022P057nsss(0)='1'  OR cVar2S14S97P034P008P015nsss(0)='1'  )then
          oVar1S553(0) <='1';
          else
          oVar1S553(0) <='0';
          end if;
        if(cVar2S0S98P005nsss(0)='1'  OR cVar2S1S98N005P069nsss(0)='1'  OR cVar2S2S98P069nsss(0)='1'  OR cVar2S3S98N069P054nsss(0)='1'  )then
          oVar1S554(0) <='1';
          else
          oVar1S554(0) <='0';
          end if;
        if(cVar2S4S98P049P043P025nsss(0)='1'  OR cVar2S5S98P049P026nsss(0)='1'  OR cVar2S6S98P049N026P027nsss(0)='1'  OR cVar2S7S98P027P049P047nsss(0)='1'  )then
          oVar1S555(0) <='1';
          else
          oVar1S555(0) <='0';
          end if;
        if(cVar2S8S98P012nsss(0)='1'  OR cVar2S9S98N012P015nsss(0)='1'  OR cVar2S10S98P015nsss(0)='1'  OR cVar2S11S98P000P012P033nsss(0)='1'  )then
          oVar1S556(0) <='1';
          else
          oVar1S556(0) <='0';
          end if;
        if(cVar2S12S98P000P012P010nsss(0)='1'  OR cVar2S13S98N000P030P031nsss(0)='1'  OR cVar2S14S98N000N030P031nsss(0)='1'  OR cVar2S15S98P052nsss(0)='1'  )then
          oVar1S557(0) <='1';
          else
          oVar1S557(0) <='0';
          end if;
        if(cVar2S16S98P067P014nsss(0)='1'  OR cVar2S17S98P012nsss(0)='1'  OR cVar2S18S98P017P014P018nsss(0)='1'  )then
          oVar1S558(0) <='1';
          else
          oVar1S558(0) <='0';
          end if;
        if(cVar1S0S99P045P030P025nsss(0)='1'  OR cVar1S1S99P045P030N025P022nsss(0)='1'  OR cVar2S2S99P023nsss(0)='1'  OR cVar2S3S99N023P024nsss(0)='1'  )then
          oVar1S559(0) <='1';
          else
          oVar1S559(0) <='0';
          end if;
        if(cVar2S4S99P029P067P024nsss(0)='1'  OR cVar2S5S99P029N067P052nsss(0)='1'  OR cVar2S6S99P029P052nsss(0)='1'  OR cVar2S7S99P024P037P067nsss(0)='1'  )then
          oVar1S560(0) <='1';
          else
          oVar1S560(0) <='0';
          end if;
        if(cVar2S8S99P024N037P008nsss(0)='1'  OR cVar2S9S99P017nsss(0)='1'  OR cVar2S10S99N017P018nsss(0)='1'  OR cVar2S11S99P054nsss(0)='1'  )then
          oVar1S561(0) <='1';
          else
          oVar1S561(0) <='0';
          end if;
        if(cVar2S12S99N054P051nsss(0)='1'  OR cVar2S13S99N054N051P052nsss(0)='1'  OR cVar2S14S99P055P008nsss(0)='1'  OR cVar2S15S99P055N008P010nsss(0)='1'  )then
          oVar1S562(0) <='1';
          else
          oVar1S562(0) <='0';
          end if;
        if(cVar2S16S99P036P013P063nsss(0)='1'  OR cVar2S17S99P036N013P010nsss(0)='1'  OR cVar2S18S99P048P017P003nsss(0)='1'  OR cVar2S19S99N048P031P013nsss(0)='1'  )then
          oVar1S563(0) <='1';
          else
          oVar1S563(0) <='0';
          end if;
        if(cVar2S0S100P005nsss(0)='1'  OR cVar2S1S100N005P069nsss(0)='1'  OR cVar2S2S100P054nsss(0)='1'  OR cVar2S3S100N054P051nsss(0)='1'  )then
          oVar1S565(0) <='1';
          else
          oVar1S565(0) <='0';
          end if;
        if(cVar2S4S100N054N051P052nsss(0)='1'  OR cVar2S5S100P055P034nsss(0)='1'  OR cVar2S6S100P055N034P015nsss(0)='1'  OR cVar2S7S100P053P012nsss(0)='1'  )then
          oVar1S566(0) <='1';
          else
          oVar1S566(0) <='0';
          end if;
        if(cVar2S8S100P053N012P000nsss(0)='1'  OR cVar2S9S100P053P056P009nsss(0)='1'  OR cVar2S10S100P053P013nsss(0)='1'  OR cVar2S11S100N053P006P014nsss(0)='1'  )then
          oVar1S567(0) <='1';
          else
          oVar1S567(0) <='0';
          end if;
        if(cVar1S12S100P019P013P045P043nsss(0)='1'  OR cVar2S13S100P012nsss(0)='1'  OR cVar2S14S100N012P066P018nsss(0)='1'  OR cVar2S15S100P018P052nsss(0)='1'  )then
          oVar1S568(0) <='1';
          else
          oVar1S568(0) <='0';
          end if;
        if(cVar2S16S100P018N052P010nsss(0)='1'  OR cVar2S17S100P048P058P015nsss(0)='1'  OR cVar2S18S100P048P016P046nsss(0)='1'  OR cVar2S19S100P020P029P015nsss(0)='1'  )then
          oVar1S569(0) <='1';
          else
          oVar1S569(0) <='0';
          end if;
        if(cVar1S0S101P045P030P035P025nsss(0)='1'  OR cVar2S1S101P022nsss(0)='1'  OR cVar2S2S101N022P023nsss(0)='1'  OR cVar2S3S101N022N023P024nsss(0)='1'  )then
          oVar1S571(0) <='1';
          else
          oVar1S571(0) <='0';
          end if;
        if(cVar2S4S101P006P044P002nsss(0)='1'  OR cVar2S5S101P006P044P016nsss(0)='1'  OR cVar2S6S101P006P036P030nsss(0)='1'  OR cVar2S7S101P012P017nsss(0)='1'  )then
          oVar1S572(0) <='1';
          else
          oVar1S572(0) <='0';
          end if;
        if(cVar2S8S101P017nsss(0)='1'  OR cVar2S9S101N017P018nsss(0)='1'  OR cVar2S10S101P069nsss(0)='1'  OR cVar2S11S101N069P028P018nsss(0)='1'  )then
          oVar1S573(0) <='1';
          else
          oVar1S573(0) <='0';
          end if;
        if(cVar2S12S101P002nsss(0)='1'  OR cVar2S13S101N002P021nsss(0)='1'  )then
          oVar1S574(0) <='1';
          else
          oVar1S574(0) <='0';
          end if;
        if(cVar1S0S102P019P045P026P005nsss(0)='1'  OR cVar2S1S102P062nsss(0)='1'  OR cVar2S2S102P069nsss(0)='1'  OR cVar2S3S102N069P028P026nsss(0)='1'  )then
          oVar1S575(0) <='1';
          else
          oVar1S575(0) <='0';
          end if;
        if(cVar2S4S102P056P053nsss(0)='1'  OR cVar2S5S102P056N053P051nsss(0)='1'  OR cVar2S6S102P056P058P012nsss(0)='1'  OR cVar2S7S102P056N058P062nsss(0)='1'  )then
          oVar1S576(0) <='1';
          else
          oVar1S576(0) <='0';
          end if;
        if(cVar2S8S102P031P068nsss(0)='1'  OR cVar2S9S102P031N068P063nsss(0)='1'  OR cVar2S10S102N031P004P034nsss(0)='1'  OR cVar2S11S102P030P033P050nsss(0)='1'  )then
          oVar1S577(0) <='1';
          else
          oVar1S577(0) <='0';
          end if;
        if(cVar2S12S102P030P033P061nsss(0)='1'  OR cVar2S13S102P030P016P017nsss(0)='1'  OR cVar2S14S102P008P055P068nsss(0)='1'  OR cVar2S15S102P050P065P013nsss(0)='1'  )then
          oVar1S578(0) <='1';
          else
          oVar1S578(0) <='0';
          end if;
        if(cVar2S16S102N050P024P016nsss(0)='1'  OR cVar2S17S102N050N024P055nsss(0)='1'  OR cVar2S18S102P017P015nsss(0)='1'  OR cVar2S19S102P034P036P014nsss(0)='1'  )then
          oVar1S579(0) <='1';
          else
          oVar1S579(0) <='0';
          end if;
        if(cVar2S20S102P064P026nsss(0)='1'  )then
          oVar1S580(0) <='1';
          else
          oVar1S580(0) <='0';
          end if;
        if(cVar1S0S103P045P030P025nsss(0)='1'  OR cVar1S1S103P045P030N025P022nsss(0)='1'  OR cVar2S2S103P023nsss(0)='1'  OR cVar2S3S103N023P024nsss(0)='1'  )then
          oVar1S581(0) <='1';
          else
          oVar1S581(0) <='0';
          end if;
        if(cVar1S4S103N045P052P065nsss(0)='1'  OR cVar1S5S103N045P052N065P062nsss(0)='1'  OR cVar2S6S103P008P014nsss(0)='1'  OR cVar2S7S103N008P010nsss(0)='1'  )then
          oVar1S582(0) <='1';
          else
          oVar1S582(0) <='0';
          end if;
        if(cVar2S8S103P005P061P019nsss(0)='1'  OR cVar2S9S103P005P008P042nsss(0)='1'  OR cVar2S10S103P039P025P067nsss(0)='1'  OR cVar2S11S103P039P025P007nsss(0)='1'  )then
          oVar1S583(0) <='1';
          else
          oVar1S583(0) <='0';
          end if;
        if(cVar2S12S103P039P016P017nsss(0)='1'  OR cVar2S13S103P003nsss(0)='1'  OR cVar2S14S103N003P013P024nsss(0)='1'  )then
          oVar1S584(0) <='1';
          else
          oVar1S584(0) <='0';
          end if;
        if(cVar1S0S104P019P045P026P005nsss(0)='1'  OR cVar2S1S104P062P069nsss(0)='1'  OR cVar2S2S104P013nsss(0)='1'  OR cVar2S3S104P055P009nsss(0)='1'  )then
          oVar1S585(0) <='1';
          else
          oVar1S585(0) <='0';
          end if;
        if(cVar2S4S104P055N009P008nsss(0)='1'  OR cVar2S5S104P051P011P012nsss(0)='1'  OR cVar2S6S104P051N011P010nsss(0)='1'  OR cVar2S7S104N051P053nsss(0)='1'  )then
          oVar1S586(0) <='1';
          else
          oVar1S586(0) <='0';
          end if;
        if(cVar2S8S104P009P044nsss(0)='1'  OR cVar2S9S104P009P036P011nsss(0)='1'  OR cVar1S10S104P019P067P047P006nsss(0)='1'  OR cVar2S11S104P049nsss(0)='1'  )then
          oVar1S587(0) <='1';
          else
          oVar1S587(0) <='0';
          end if;
        if(cVar2S12S104P049P018nsss(0)='1'  OR cVar2S13S104P018P005P012nsss(0)='1'  OR cVar2S14S104N018P054P012nsss(0)='1'  OR cVar2S15S104P014P036nsss(0)='1'  )then
          oVar1S588(0) <='1';
          else
          oVar1S588(0) <='0';
          end if;
        if(cVar2S16S104P014N036P011nsss(0)='1'  OR cVar1S17S104P019P067P024P042nsss(0)='1'  OR cVar2S18S104P052nsss(0)='1'  OR cVar2S19S104P063P018nsss(0)='1'  )then
          oVar1S589(0) <='1';
          else
          oVar1S589(0) <='0';
          end if;
        if(cVar1S0S105P045P030P035P025nsss(0)='1'  OR cVar2S1S105P022nsss(0)='1'  OR cVar2S2S105N022P057nsss(0)='1'  OR cVar2S3S105P051nsss(0)='1'  )then
          oVar1S591(0) <='1';
          else
          oVar1S591(0) <='0';
          end if;
        if(cVar2S4S105N051P000P033nsss(0)='1'  OR cVar2S5S105P052P008nsss(0)='1'  OR cVar2S6S105N052P035P051nsss(0)='1'  OR cVar2S7S105P064P000P051nsss(0)='1'  )then
          oVar1S592(0) <='1';
          else
          oVar1S592(0) <='0';
          end if;
        if(cVar2S8S105P064N000P020nsss(0)='1'  OR cVar2S9S105P064P057nsss(0)='1'  OR cVar1S10S105N045N029P043P022nsss(0)='1'  OR cVar2S11S105P050P008P019nsss(0)='1'  )then
          oVar1S593(0) <='1';
          else
          oVar1S593(0) <='0';
          end if;
        if(cVar2S0S106P051P011P069nsss(0)='1'  OR cVar2S1S106P051N011P008nsss(0)='1'  OR cVar2S2S106N051P045nsss(0)='1'  OR cVar2S3S106N051N045P007nsss(0)='1'  )then
          oVar1S595(0) <='1';
          else
          oVar1S595(0) <='0';
          end if;
        if(cVar2S4S106P042nsss(0)='1'  OR cVar2S5S106N042P007P014nsss(0)='1'  OR cVar2S6S106N042N007P030nsss(0)='1'  OR cVar1S7S106P020P039P041P033nsss(0)='1'  )then
          oVar1S596(0) <='1';
          else
          oVar1S596(0) <='0';
          end if;
        if(cVar2S8S106P003nsss(0)='1'  OR cVar2S9S106N003P033nsss(0)='1'  OR cVar2S10S106N003N033P014nsss(0)='1'  OR cVar1S11S106P020P039P041nsss(0)='1'  )then
          oVar1S597(0) <='1';
          else
          oVar1S597(0) <='0';
          end if;
        if(cVar2S12S106P011P036nsss(0)='1'  OR cVar2S13S106P011N036P062nsss(0)='1'  OR cVar2S14S106P035P034nsss(0)='1'  )then
          oVar1S598(0) <='1';
          else
          oVar1S598(0) <='0';
          end if;
        if(cVar2S0S107P000nsss(0)='1'  OR cVar2S1S107P069P015nsss(0)='1'  OR cVar2S2S107P069P015P049nsss(0)='1'  OR cVar2S3S107P018P053nsss(0)='1'  )then
          oVar1S599(0) <='1';
          else
          oVar1S599(0) <='0';
          end if;
        if(cVar1S4S107N051P053P007P025nsss(0)='1'  OR cVar2S5S107P065P009P011nsss(0)='1'  OR cVar2S6S107P065N009P055nsss(0)='1'  OR cVar2S7S107P065P006P034nsss(0)='1'  )then
          oVar1S600(0) <='1';
          else
          oVar1S600(0) <='0';
          end if;
        if(cVar2S8S107P025P059P004nsss(0)='1'  OR cVar2S9S107P025P010P024nsss(0)='1'  OR cVar2S10S107P037P062nsss(0)='1'  OR cVar2S11S107P016P013P036nsss(0)='1'  )then
          oVar1S601(0) <='1';
          else
          oVar1S601(0) <='0';
          end if;
        if(cVar2S0S108P024nsss(0)='1'  OR cVar2S1S108P024P012P016nsss(0)='1'  OR cVar2S2S108P022nsss(0)='1'  OR cVar2S3S108N022P025nsss(0)='1'  )then
          oVar1S603(0) <='1';
          else
          oVar1S603(0) <='0';
          end if;
        if(cVar2S4S108N022N025P030nsss(0)='1'  OR cVar2S5S108P041P020nsss(0)='1'  OR cVar2S6S108P041N020P016nsss(0)='1'  OR cVar2S7S108N041P043nsss(0)='1'  )then
          oVar1S604(0) <='1';
          else
          oVar1S604(0) <='0';
          end if;
        if(cVar2S8S108N041P043P003nsss(0)='1'  OR cVar2S9S108P057P012nsss(0)='1'  OR cVar2S10S108P057N012P014nsss(0)='1'  OR cVar2S11S108N057P006nsss(0)='1'  )then
          oVar1S605(0) <='1';
          else
          oVar1S605(0) <='0';
          end if;
        if(cVar2S12S108P032nsss(0)='1'  OR cVar2S13S108P058nsss(0)='1'  OR cVar2S14S108P059P031nsss(0)='1'  OR cVar2S15S108N059P032nsss(0)='1'  )then
          oVar1S606(0) <='1';
          else
          oVar1S606(0) <='0';
          end if;
        if(cVar2S16S108N059N032P055nsss(0)='1'  )then
          oVar1S607(0) <='1';
          else
          oVar1S607(0) <='0';
          end if;
        if(cVar1S0S109P022P043nsss(0)='1'  OR cVar1S1S109P022N043P002nsss(0)='1'  OR cVar2S2S109P033nsss(0)='1'  OR cVar2S3S109P030nsss(0)='1'  )then
          oVar1S608(0) <='1';
          else
          oVar1S608(0) <='0';
          end if;
        if(cVar2S4S109N030P013P031nsss(0)='1'  OR cVar2S5S109P054P053P028nsss(0)='1'  OR cVar2S6S109P054P044nsss(0)='1'  OR cVar1S7S109N022P043P025nsss(0)='1'  )then
          oVar1S609(0) <='1';
          else
          oVar1S609(0) <='0';
          end if;
        if(cVar2S8S109P023nsss(0)='1'  OR cVar2S9S109N023P034P006nsss(0)='1'  )then
          oVar1S610(0) <='1';
          else
          oVar1S610(0) <='0';
          end if;
        if(cVar2S0S110P009P069nsss(0)='1'  OR cVar2S1S110N009P011P012nsss(0)='1'  OR cVar2S2S110N009N011P008nsss(0)='1'  OR cVar2S3S110P069P015nsss(0)='1'  )then
          oVar1S611(0) <='1';
          else
          oVar1S611(0) <='0';
          end if;
        if(cVar2S4S110P069P015P008nsss(0)='1'  OR cVar2S5S110P023nsss(0)='1'  OR cVar2S6S110N023P025nsss(0)='1'  OR cVar2S7S110P042P023nsss(0)='1'  )then
          oVar1S612(0) <='1';
          else
          oVar1S612(0) <='0';
          end if;
        if(cVar2S8S110P042P023P045nsss(0)='1'  OR cVar2S9S110P042P005nsss(0)='1'  OR cVar2S10S110P064P066nsss(0)='1'  OR cVar2S11S110P056P048nsss(0)='1'  )then
          oVar1S613(0) <='1';
          else
          oVar1S613(0) <='0';
          end if;
        if(cVar2S0S111P011P069nsss(0)='1'  OR cVar2S1S111N011P008nsss(0)='1'  OR cVar2S2S111N011N008P009nsss(0)='1'  OR cVar2S3S111P064nsss(0)='1'  )then
          oVar1S615(0) <='1';
          else
          oVar1S615(0) <='0';
          end if;
        if(cVar2S4S111N064P059P054nsss(0)='1'  OR cVar1S5S111N053P044P025nsss(0)='1'  OR cVar1S6S111N053P044N025P023nsss(0)='1'  OR cVar2S7S111P026P022nsss(0)='1'  )then
          oVar1S616(0) <='1';
          else
          oVar1S616(0) <='0';
          end if;
        if(cVar2S8S111P056P004P039nsss(0)='1'  OR cVar2S9S111N056P054P022nsss(0)='1'  OR cVar2S10S111P045nsss(0)='1'  OR cVar2S11S111N045P064nsss(0)='1'  )then
          oVar1S617(0) <='1';
          else
          oVar1S617(0) <='0';
          end if;
        if(cVar1S12S111N053N044P042P005nsss(0)='1'  OR cVar2S13S111P009P016P018nsss(0)='1'  )then
          oVar1S618(0) <='1';
          else
          oVar1S618(0) <='0';
          end if;
        if(cVar1S0S112P044P023nsss(0)='1'  OR cVar1S1S112P044N023P025nsss(0)='1'  OR cVar2S2S112P000P013P058nsss(0)='1'  OR cVar2S3S112P000P013P067nsss(0)='1'  )then
          oVar1S619(0) <='1';
          else
          oVar1S619(0) <='0';
          end if;
        if(cVar2S4S112P041P053P000nsss(0)='1'  OR cVar2S5S112P041N053P069nsss(0)='1'  OR cVar2S6S112P053P041P020nsss(0)='1'  OR cVar2S7S112P053N041P039nsss(0)='1'  )then
          oVar1S620(0) <='1';
          else
          oVar1S620(0) <='0';
          end if;
        if(cVar2S8S112P045nsss(0)='1'  OR cVar2S9S112N045P064nsss(0)='1'  OR cVar2S10S112P063nsss(0)='1'  OR cVar2S11S112N063P068nsss(0)='1'  )then
          oVar1S621(0) <='1';
          else
          oVar1S621(0) <='0';
          end if;
        if(cVar1S0S113P044P025nsss(0)='1'  OR cVar1S1S113P044N025P023nsss(0)='1'  OR cVar2S2S113P000P013nsss(0)='1'  OR cVar2S3S113P041P053P000nsss(0)='1'  )then
          oVar1S623(0) <='1';
          else
          oVar1S623(0) <='0';
          end if;
        if(cVar2S4S113P041N053P069nsss(0)='1'  OR cVar2S5S113P041P020nsss(0)='1'  OR cVar2S6S113P041N020P016nsss(0)='1'  OR cVar2S7S113N041P039P016nsss(0)='1'  )then
          oVar1S624(0) <='1';
          else
          oVar1S624(0) <='0';
          end if;
        if(cVar2S8S113P045nsss(0)='1'  OR cVar2S9S113N045P034P035nsss(0)='1'  OR cVar2S10S113P063nsss(0)='1'  OR cVar2S11S113N063P068nsss(0)='1'  )then
          oVar1S625(0) <='1';
          else
          oVar1S625(0) <='0';
          end if;
        if(cVar1S0S114P016P044P023nsss(0)='1'  OR cVar1S1S114P016P044N023P025nsss(0)='1'  OR cVar2S2S114P026P048P022nsss(0)='1'  OR cVar1S3S114P016N044P041P020nsss(0)='1'  )then
          oVar1S627(0) <='1';
          else
          oVar1S627(0) <='0';
          end if;
        if(cVar2S4S114P062P061nsss(0)='1'  OR cVar2S5S114P004P008P017nsss(0)='1'  OR cVar2S6S114P004N008P047nsss(0)='1'  OR cVar2S7S114P004P003P006nsss(0)='1'  )then
          oVar1S628(0) <='1';
          else
          oVar1S628(0) <='0';
          end if;
        if(cVar2S8S114P040nsss(0)='1'  OR cVar2S9S114N040P064P007nsss(0)='1'  OR cVar2S10S114P002P015P003nsss(0)='1'  OR cVar2S11S114P002P066P068nsss(0)='1'  )then
          oVar1S629(0) <='1';
          else
          oVar1S629(0) <='0';
          end if;
        if(cVar2S12S114P002N066P009nsss(0)='1'  OR cVar2S13S114P069P010P012nsss(0)='1'  OR cVar2S14S114P018nsss(0)='1'  OR cVar1S15S114P016P039P005nsss(0)='1'  )then
          oVar1S630(0) <='1';
          else
          oVar1S630(0) <='0';
          end if;
        if(cVar2S16S114P034nsss(0)='1'  )then
          oVar1S631(0) <='1';
          else
          oVar1S631(0) <='0';
          end if;
        if(cVar1S0S115P044P025nsss(0)='1'  OR cVar1S1S115P044N025P023nsss(0)='1'  OR cVar2S2S115P000P056P006nsss(0)='1'  OR cVar2S3S115P031P032nsss(0)='1'  )then
          oVar1S632(0) <='1';
          else
          oVar1S632(0) <='0';
          end if;
        if(cVar2S4S115P031P032P068nsss(0)='1'  OR cVar2S5S115P031P059nsss(0)='1'  OR cVar2S6S115P016P022nsss(0)='1'  OR cVar2S7S115P016P022P018nsss(0)='1'  )then
          oVar1S633(0) <='1';
          else
          oVar1S633(0) <='0';
          end if;
        if(cVar2S8S115N016P022P043nsss(0)='1'  OR cVar2S9S115P006nsss(0)='1'  OR cVar2S10S115N006P045nsss(0)='1'  OR cVar2S11S115N006N045P064nsss(0)='1'  )then
          oVar1S634(0) <='1';
          else
          oVar1S634(0) <='0';
          end if;
        if(cVar1S12S115N044P042P024P005nsss(0)='1'  OR cVar2S13S115P009P062P004nsss(0)='1'  )then
          oVar1S635(0) <='1';
          else
          oVar1S635(0) <='0';
          end if;
        if(cVar1S0S116P016P044P023nsss(0)='1'  OR cVar1S1S116P016P044N023P025nsss(0)='1'  OR cVar2S2S116P026P048nsss(0)='1'  OR cVar1S3S116P016N044P041P020nsss(0)='1'  )then
          oVar1S636(0) <='1';
          else
          oVar1S636(0) <='0';
          end if;
        if(cVar2S4S116P062P061nsss(0)='1'  OR cVar2S5S116P010P028P014nsss(0)='1'  OR cVar2S6S116P010N028P039nsss(0)='1'  OR cVar2S7S116N010P027P014nsss(0)='1'  )then
          oVar1S637(0) <='1';
          else
          oVar1S637(0) <='0';
          end if;
        if(cVar2S8S116N010N027P020nsss(0)='1'  OR cVar2S9S116P003P040nsss(0)='1'  OR cVar2S10S116P002P015P013nsss(0)='1'  OR cVar2S11S116P002P066P067nsss(0)='1'  )then
          oVar1S638(0) <='1';
          else
          oVar1S638(0) <='0';
          end if;
        if(cVar2S12S116P002N066P004nsss(0)='1'  OR cVar2S13S116P019P011nsss(0)='1'  OR cVar2S14S116P010P012nsss(0)='1'  OR cVar1S15S116P016P039P005nsss(0)='1'  )then
          oVar1S639(0) <='1';
          else
          oVar1S639(0) <='0';
          end if;
        if(cVar2S16S116P034nsss(0)='1'  )then
          oVar1S640(0) <='1';
          else
          oVar1S640(0) <='0';
          end if;
        if(cVar1S0S117P044P025nsss(0)='1'  OR cVar1S1S117P044N025P023nsss(0)='1'  OR cVar2S2S117P000P056P067nsss(0)='1'  OR cVar2S3S117P005P039P029nsss(0)='1'  )then
          oVar1S641(0) <='1';
          else
          oVar1S641(0) <='0';
          end if;
        if(cVar2S4S117P005P039P003nsss(0)='1'  OR cVar2S5S117P005P031P020nsss(0)='1'  OR cVar2S6S117P038nsss(0)='1'  OR cVar2S7S117N038P054P030nsss(0)='1'  )then
          oVar1S642(0) <='1';
          else
          oVar1S642(0) <='0';
          end if;
        if(cVar2S8S117P002nsss(0)='1'  OR cVar2S9S117N002P069nsss(0)='1'  OR cVar2S10S117N002N069P064nsss(0)='1'  OR cVar1S11S117N044P023P024P005nsss(0)='1'  )then
          oVar1S643(0) <='1';
          else
          oVar1S643(0) <='0';
          end if;
        if(cVar2S12S117P068nsss(0)='1'  )then
          oVar1S644(0) <='1';
          else
          oVar1S644(0) <='0';
          end if;
        if(cVar1S0S118P044P025nsss(0)='1'  OR cVar1S1S118P044N025P023nsss(0)='1'  OR cVar2S2S118P000P056nsss(0)='1'  OR cVar2S3S118P005P039nsss(0)='1'  )then
          oVar1S645(0) <='1';
          else
          oVar1S645(0) <='0';
          end if;
        if(cVar2S4S118P005P039P003nsss(0)='1'  OR cVar2S5S118P005P031P041nsss(0)='1'  OR cVar2S6S118P038nsss(0)='1'  OR cVar2S7S118P002nsss(0)='1'  )then
          oVar1S646(0) <='1';
          else
          oVar1S646(0) <='0';
          end if;
        if(cVar2S8S118N002P069nsss(0)='1'  OR cVar2S9S118N002N069P003nsss(0)='1'  OR cVar1S10S118N044P023P024P005nsss(0)='1'  OR cVar2S11S118P068nsss(0)='1'  )then
          oVar1S647(0) <='1';
          else
          oVar1S647(0) <='0';
          end if;
        if(cVar1S0S119P044P025nsss(0)='1'  OR cVar1S1S119P044N025P023nsss(0)='1'  OR cVar2S2S119P032P013P058nsss(0)='1'  OR cVar2S3S119P004P051nsss(0)='1'  )then
          oVar1S649(0) <='1';
          else
          oVar1S649(0) <='0';
          end if;
        if(cVar2S4S119P051P041P020nsss(0)='1'  OR cVar2S5S119P002nsss(0)='1'  OR cVar2S6S119N002P063nsss(0)='1'  OR cVar2S7S119N002N063P069nsss(0)='1'  )then
          oVar1S650(0) <='1';
          else
          oVar1S650(0) <='0';
          end if;
        if(cVar1S8S119N044P023P024P008nsss(0)='1'  OR cVar2S9S119P069P036nsss(0)='1'  OR cVar2S10S119P069N036P068nsss(0)='1'  )then
          oVar1S651(0) <='1';
          else
          oVar1S651(0) <='0';
          end if;
        if(cVar1S0S120P044P025nsss(0)='1'  OR cVar1S1S120P044N025P023nsss(0)='1'  OR cVar2S2S120P032P013nsss(0)='1'  OR cVar2S3S120P056P030P057nsss(0)='1'  )then
          oVar1S652(0) <='1';
          else
          oVar1S652(0) <='0';
          end if;
        if(cVar2S4S120P056P058nsss(0)='1'  OR cVar2S5S120P056P004nsss(0)='1'  OR cVar2S6S120P062P065nsss(0)='1'  OR cVar2S7S120P062N065P068nsss(0)='1'  )then
          oVar1S653(0) <='1';
          else
          oVar1S653(0) <='0';
          end if;
        if(cVar1S8S120N044P023P024P005nsss(0)='1'  OR cVar2S9S120P068nsss(0)='1'  )then
          oVar1S654(0) <='1';
          else
          oVar1S654(0) <='0';
          end if;
        if(cVar1S0S121P042P023nsss(0)='1'  OR cVar1S1S121P042N023P002nsss(0)='1'  OR cVar1S2S121P042N023N002P055nsss(0)='1'  OR cVar2S3S121P006P044nsss(0)='1'  )then
          oVar1S655(0) <='1';
          else
          oVar1S655(0) <='0';
          end if;
        if(cVar2S4S121N006P024P065nsss(0)='1'  OR cVar2S5S121P036nsss(0)='1'  OR cVar2S6S121P062nsss(0)='1'  OR cVar2S7S121N062P050P013nsss(0)='1'  )then
          oVar1S656(0) <='1';
          else
          oVar1S656(0) <='0';
          end if;
        if(cVar2S8S121N062N050P053nsss(0)='1'  OR cVar2S9S121P046P025nsss(0)='1'  OR cVar2S10S121N046P025P045nsss(0)='1'  OR cVar2S11S121P004P063P048nsss(0)='1'  )then
          oVar1S657(0) <='1';
          else
          oVar1S657(0) <='0';
          end if;
        if(cVar1S12S121N042P023P024P008nsss(0)='1'  OR cVar2S13S121P069P036nsss(0)='1'  OR cVar2S14S121P069N036P068nsss(0)='1'  )then
          oVar1S658(0) <='1';
          else
          oVar1S658(0) <='0';
          end if;
        if(cVar1S0S122P044P026P025nsss(0)='1'  OR cVar2S1S122P023nsss(0)='1'  OR cVar2S2S122N023P032P067nsss(0)='1'  OR cVar2S3S122P039nsss(0)='1'  )then
          oVar1S659(0) <='1';
          else
          oVar1S659(0) <='0';
          end if;
        if(cVar2S4S122N039P062P008nsss(0)='1'  OR cVar2S5S122N039P062P014nsss(0)='1'  OR cVar2S6S122P039P059P004nsss(0)='1'  OR cVar2S7S122P039N059P061nsss(0)='1'  )then
          oVar1S660(0) <='1';
          else
          oVar1S660(0) <='0';
          end if;
        if(cVar2S8S122P039P012P050nsss(0)='1'  OR cVar2S9S122P062P063nsss(0)='1'  OR cVar2S10S122P062N063P003nsss(0)='1'  OR cVar1S11S122N044P023P024P006nsss(0)='1'  )then
          oVar1S661(0) <='1';
          else
          oVar1S661(0) <='0';
          end if;
        if(cVar2S12S122P045nsss(0)='1'  OR cVar2S13S122N045P069P014nsss(0)='1'  )then
          oVar1S662(0) <='1';
          else
          oVar1S662(0) <='0';
          end if;
        if(cVar1S0S123P042P023nsss(0)='1'  OR cVar1S1S123P042N023P002nsss(0)='1'  OR cVar1S2S123P042N023N002P055nsss(0)='1'  OR cVar2S3S123P006P044nsss(0)='1'  )then
          oVar1S663(0) <='1';
          else
          oVar1S663(0) <='0';
          end if;
        if(cVar2S4S123N006P024P065nsss(0)='1'  OR cVar2S5S123P067P069nsss(0)='1'  OR cVar2S6S123P067P069P014nsss(0)='1'  OR cVar2S7S123P067P024P055nsss(0)='1'  )then
          oVar1S664(0) <='1';
          else
          oVar1S664(0) <='0';
          end if;
        if(cVar2S8S123P046nsss(0)='1'  OR cVar2S9S123P045P029nsss(0)='1'  OR cVar2S10S123P045N029P009nsss(0)='1'  OR cVar2S11S123P051P011nsss(0)='1'  )then
          oVar1S665(0) <='1';
          else
          oVar1S665(0) <='0';
          end if;
        if(cVar2S12S123P051N011P010nsss(0)='1'  OR cVar2S13S123N051P038P040nsss(0)='1'  OR cVar1S14S123N042P023P024P007nsss(0)='1'  OR cVar2S15S123P005nsss(0)='1'  )then
          oVar1S666(0) <='1';
          else
          oVar1S666(0) <='0';
          end if;
        if(cVar2S0S124P003nsss(0)='1'  OR cVar2S1S124N003P020nsss(0)='1'  OR cVar2S2S124N003N020P013nsss(0)='1'  OR cVar2S3S124P063P058nsss(0)='1'  )then
          oVar1S668(0) <='1';
          else
          oVar1S668(0) <='0';
          end if;
        if(cVar2S4S124P063N058P001nsss(0)='1'  OR cVar2S5S124N063P065nsss(0)='1'  OR cVar2S6S124P006P021P044nsss(0)='1'  OR cVar2S7S124P006P012P014nsss(0)='1'  )then
          oVar1S669(0) <='1';
          else
          oVar1S669(0) <='0';
          end if;
        if(cVar2S8S124P007P015nsss(0)='1'  OR cVar2S9S124P007P015P014nsss(0)='1'  OR cVar2S10S124P006P066nsss(0)='1'  OR cVar2S11S124N006P009P065nsss(0)='1'  )then
          oVar1S670(0) <='1';
          else
          oVar1S670(0) <='0';
          end if;
        if(cVar2S12S124P016nsss(0)='1'  OR cVar1S13S124P019P051P042P067nsss(0)='1'  OR cVar2S14S124P037nsss(0)='1'  OR cVar2S15S124N037P015nsss(0)='1'  )then
          oVar1S671(0) <='1';
          else
          oVar1S671(0) <='0';
          end if;
        if(cVar2S16S124P013P048P005nsss(0)='1'  OR cVar2S17S124P013P048P016nsss(0)='1'  OR cVar2S18S124P010nsss(0)='1'  OR cVar2S19S124N010P067P013nsss(0)='1'  )then
          oVar1S672(0) <='1';
          else
          oVar1S672(0) <='0';
          end if;
        if(cVar2S20S124P061nsss(0)='1'  OR cVar2S21S124N061P017P014nsss(0)='1'  OR cVar2S22S124P026nsss(0)='1'  OR cVar2S23S124N026P017P014nsss(0)='1'  )then
          oVar1S673(0) <='1';
          else
          oVar1S673(0) <='0';
          end if;
        if(cVar2S0S125P061P033nsss(0)='1'  OR cVar2S1S125P061N033P064nsss(0)='1'  OR cVar2S2S125N061P059nsss(0)='1'  OR cVar2S3S125P013P014nsss(0)='1'  )then
          oVar1S675(0) <='1';
          else
          oVar1S675(0) <='0';
          end if;
        if(cVar2S4S125P013P014P016nsss(0)='1'  OR cVar2S5S125P016nsss(0)='1'  OR cVar2S6S125P013nsss(0)='1'  OR cVar2S7S125P056P034nsss(0)='1'  )then
          oVar1S676(0) <='1';
          else
          oVar1S676(0) <='0';
          end if;
        if(cVar2S8S125P056N034P016nsss(0)='1'  OR cVar2S9S125P016P010nsss(0)='1'  OR cVar2S10S125P020nsss(0)='1'  OR cVar2S11S125N020P012nsss(0)='1'  )then
          oVar1S677(0) <='1';
          else
          oVar1S677(0) <='0';
          end if;
        if(cVar2S12S125P032nsss(0)='1'  OR cVar2S13S125N032P034nsss(0)='1'  OR cVar2S14S125N032N034P016nsss(0)='1'  OR cVar2S15S125P044P054P031nsss(0)='1'  )then
          oVar1S678(0) <='1';
          else
          oVar1S678(0) <='0';
          end if;
        if(cVar2S16S125P044P054P065nsss(0)='1'  OR cVar2S17S125P062nsss(0)='1'  OR cVar2S18S125P042P030P012nsss(0)='1'  OR cVar2S19S125P042N030P028nsss(0)='1'  )then
          oVar1S679(0) <='1';
          else
          oVar1S679(0) <='0';
          end if;
        if(cVar2S20S125P042P040nsss(0)='1'  )then
          oVar1S680(0) <='1';
          else
          oVar1S680(0) <='0';
          end if;
        if(cVar2S0S126P042nsss(0)='1'  OR cVar2S1S126N042P013P011nsss(0)='1'  OR cVar2S2S126N042N013P015nsss(0)='1'  OR cVar2S3S126P030P059nsss(0)='1'  )then
          oVar1S681(0) <='1';
          else
          oVar1S681(0) <='0';
          end if;
        if(cVar2S4S126P030N059P031nsss(0)='1'  OR cVar2S5S126N030P055P017nsss(0)='1'  OR cVar2S6S126N030P055P063nsss(0)='1'  OR cVar2S7S126P006P062P064nsss(0)='1'  )then
          oVar1S682(0) <='1';
          else
          oVar1S682(0) <='0';
          end if;
        if(cVar2S8S126P006N062psss(0)='1'  OR cVar2S9S126P036P006P019nsss(0)='1'  OR cVar2S10S126P036N006P055nsss(0)='1'  OR cVar1S11S126P018P014P060P032nsss(0)='1'  )then
          oVar1S683(0) <='1';
          else
          oVar1S683(0) <='0';
          end if;
        if(cVar2S12S126P034nsss(0)='1'  OR cVar2S13S126N034P016P067nsss(0)='1'  OR cVar2S14S126N034P016P017nsss(0)='1'  OR cVar2S15S126P046P027P017nsss(0)='1'  )then
          oVar1S684(0) <='1';
          else
          oVar1S684(0) <='0';
          end if;
        if(cVar1S16S126P018P061P033nsss(0)='1'  OR cVar2S17S126P011P067nsss(0)='1'  OR cVar2S18S126N011P035P062nsss(0)='1'  OR cVar2S19S126N011N035P036nsss(0)='1'  )then
          oVar1S685(0) <='1';
          else
          oVar1S685(0) <='0';
          end if;
        if(cVar1S20S126P018N061P042P063nsss(0)='1'  OR cVar2S21S126P010P016P014nsss(0)='1'  OR cVar2S22S126P010P016P015nsss(0)='1'  OR cVar2S23S126P001P009nsss(0)='1'  )then
          oVar1S686(0) <='1';
          else
          oVar1S686(0) <='0';
          end if;
        if(cVar2S24S126N001P023P003nsss(0)='1'  OR cVar2S25S126P000P049nsss(0)='1'  )then
          oVar1S687(0) <='1';
          else
          oVar1S687(0) <='0';
          end if;
        if(cVar2S0S127P036nsss(0)='1'  OR cVar2S1S127N036P028nsss(0)='1'  OR cVar2S2S127N036N028P035nsss(0)='1'  OR cVar2S3S127P032P019nsss(0)='1'  )then
          oVar1S688(0) <='1';
          else
          oVar1S688(0) <='0';
          end if;
        if(cVar2S4S127P032P019P016nsss(0)='1'  OR cVar2S5S127N032P023nsss(0)='1'  OR cVar2S6S127P010P032P056nsss(0)='1'  OR cVar2S7S127P010P032P059nsss(0)='1'  )then
          oVar1S689(0) <='1';
          else
          oVar1S689(0) <='0';
          end if;
        if(cVar2S8S127P010P006P019nsss(0)='1'  OR cVar2S9S127P068P013P018nsss(0)='1'  OR cVar2S10S127P068N013P012nsss(0)='1'  OR cVar2S11S127P028P016nsss(0)='1'  )then
          oVar1S690(0) <='1';
          else
          oVar1S690(0) <='0';
          end if;
        if(cVar2S12S127P028P016P040nsss(0)='1'  OR cVar2S13S127P061P020nsss(0)='1'  OR cVar2S14S127P061P013P016nsss(0)='1'  OR cVar2S15S127P063nsss(0)='1'  )then
          oVar1S691(0) <='1';
          else
          oVar1S691(0) <='0';
          end if;
        if(cVar2S16S127N063P010P016nsss(0)='1'  OR cVar1S17S127N017P018P027P014nsss(0)='1'  OR cVar2S18S127P004nsss(0)='1'  OR cVar2S19S127N004P016P014nsss(0)='1'  )then
          oVar1S692(0) <='1';
          else
          oVar1S692(0) <='0';
          end if;
        if(cVar2S20S127P050P044nsss(0)='1'  OR cVar2S21S127P050N044P025nsss(0)='1'  OR cVar2S22S127P050P029nsss(0)='1'  OR cVar2S23S127P036P035P039nsss(0)='1'  )then
          oVar1S693(0) <='1';
          else
          oVar1S693(0) <='0';
          end if;
        if(cVar2S24S127P036P035P014nsss(0)='1'  OR cVar2S25S127P036P016P011nsss(0)='1'  OR cVar2S26S127P011P055nsss(0)='1'  OR cVar2S27S127P011N055P000nsss(0)='1'  )then
          oVar1S694(0) <='1';
          else
          oVar1S694(0) <='0';
          end if;
        if(cVar2S28S127N011P036P026nsss(0)='1'  OR cVar2S29S127P027nsss(0)='1'  OR cVar2S30S127N027P007P011nsss(0)='1'  OR cVar2S31S127N027N007P065nsss(0)='1'  )then
          oVar1S695(0) <='1';
          else
          oVar1S695(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV4 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar1S0(0)='1'  OR oVar1S1(0)='1'  OR oVar1S2(0)='1'  OR oVar1S3(0)='1'  )then
          oVar2S0(0) <='1';
          else
          oVar2S0(0) <='0';
          end if;
        if(oVar1S4(0)='1'  )then
          oVar2S1(0) <='1';
          else
          oVar2S1(0) <='0';
          end if;
        if(oVar1S5(0)='1'  OR oVar1S6(0)='1'  OR oVar1S7(0)='1'  OR oVar1S8(0)='1'  )then
          oVar2S2(0) <='1';
          else
          oVar2S2(0) <='0';
          end if;
        if(oVar1S9(0)='1'  OR oVar1S10(0)='1'  OR oVar1S11(0)='1'  )then
          oVar2S3(0) <='1';
          else
          oVar2S3(0) <='0';
          end if;
        if(oVar1S12(0)='1'  OR oVar1S13(0)='1'  OR oVar1S14(0)='1'  OR oVar1S15(0)='1'  )then
          oVar2S4(0) <='1';
          else
          oVar2S4(0) <='0';
          end if;
        if(oVar1S16(0)='1'  OR oVar1S17(0)='1'  OR oVar1S18(0)='1'  )then
          oVar2S5(0) <='1';
          else
          oVar2S5(0) <='0';
          end if;
        if(oVar1S19(0)='1'  OR oVar1S20(0)='1'  OR oVar1S21(0)='1'  OR oVar1S22(0)='1'  )then
          oVar2S6(0) <='1';
          else
          oVar2S6(0) <='0';
          end if;
        if(oVar1S23(0)='1'  )then
          oVar2S7(0) <='1';
          else
          oVar2S7(0) <='0';
          end if;
        if(oVar1S24(0)='1'  OR oVar1S25(0)='1'  OR oVar1S26(0)='1'  OR oVar1S27(0)='1'  )then
          oVar2S8(0) <='1';
          else
          oVar2S8(0) <='0';
          end if;
        if(oVar1S28(0)='1'  OR oVar1S29(0)='1'  OR oVar1S30(0)='1'  )then
          oVar2S9(0) <='1';
          else
          oVar2S9(0) <='0';
          end if;
        if(oVar1S31(0)='1'  OR oVar1S32(0)='1'  OR oVar1S33(0)='1'  OR oVar1S34(0)='1'  )then
          oVar2S10(0) <='1';
          else
          oVar2S10(0) <='0';
          end if;
        if(oVar1S35(0)='1'  OR oVar1S36(0)='1'  )then
          oVar2S11(0) <='1';
          else
          oVar2S11(0) <='0';
          end if;
        if(oVar1S37(0)='1'  OR oVar1S38(0)='1'  OR oVar1S39(0)='1'  OR oVar1S40(0)='1'  )then
          oVar2S12(0) <='1';
          else
          oVar2S12(0) <='0';
          end if;
        if(oVar1S41(0)='1'  OR oVar1S42(0)='1'  OR oVar1S43(0)='1'  OR oVar1S44(0)='1'  )then
          oVar2S14(0) <='1';
          else
          oVar2S14(0) <='0';
          end if;
        if(oVar1S45(0)='1'  )then
          oVar2S15(0) <='1';
          else
          oVar2S15(0) <='0';
          end if;
        if(oVar1S47(0)='1'  OR oVar1S48(0)='1'  OR oVar1S49(0)='1'  OR oVar1S50(0)='1'  )then
          oVar2S16(0) <='1';
          else
          oVar2S16(0) <='0';
          end if;
        if(oVar1S51(0)='1'  OR oVar1S52(0)='1'  )then
          oVar2S17(0) <='1';
          else
          oVar2S17(0) <='0';
          end if;
        if(oVar1S53(0)='1'  OR oVar1S54(0)='1'  OR oVar1S55(0)='1'  OR oVar1S56(0)='1'  )then
          oVar2S18(0) <='1';
          else
          oVar2S18(0) <='0';
          end if;
        if(oVar1S57(0)='1'  )then
          oVar2S19(0) <='1';
          else
          oVar2S19(0) <='0';
          end if;
        if(oVar1S58(0)='1'  OR oVar1S59(0)='1'  OR oVar1S60(0)='1'  OR oVar1S61(0)='1'  )then
          oVar2S20(0) <='1';
          else
          oVar2S20(0) <='0';
          end if;
        if(oVar1S62(0)='1'  OR oVar1S63(0)='1'  )then
          oVar2S21(0) <='1';
          else
          oVar2S21(0) <='0';
          end if;
        if(oVar1S65(0)='1'  OR oVar1S66(0)='1'  OR oVar1S67(0)='1'  OR oVar1S68(0)='1'  )then
          oVar2S22(0) <='1';
          else
          oVar2S22(0) <='0';
          end if;
        if(oVar1S69(0)='1'  )then
          oVar2S23(0) <='1';
          else
          oVar2S23(0) <='0';
          end if;
        if(oVar1S70(0)='1'  OR oVar1S71(0)='1'  OR oVar1S72(0)='1'  OR oVar1S73(0)='1'  )then
          oVar2S24(0) <='1';
          else
          oVar2S24(0) <='0';
          end if;
        if(oVar1S74(0)='1'  OR oVar1S75(0)='1'  )then
          oVar2S25(0) <='1';
          else
          oVar2S25(0) <='0';
          end if;
        if(oVar1S77(0)='1'  OR oVar1S78(0)='1'  OR oVar1S79(0)='1'  OR oVar1S80(0)='1'  )then
          oVar2S26(0) <='1';
          else
          oVar2S26(0) <='0';
          end if;
        if(oVar1S81(0)='1'  )then
          oVar2S27(0) <='1';
          else
          oVar2S27(0) <='0';
          end if;
        if(oVar1S83(0)='1'  OR oVar1S84(0)='1'  OR oVar1S85(0)='1'  OR oVar1S86(0)='1'  )then
          oVar2S28(0) <='1';
          else
          oVar2S28(0) <='0';
          end if;
        if(oVar1S87(0)='1'  OR oVar1S88(0)='1'  OR oVar1S89(0)='1'  )then
          oVar2S29(0) <='1';
          else
          oVar2S29(0) <='0';
          end if;
        if(oVar1S90(0)='1'  OR oVar1S91(0)='1'  OR oVar1S92(0)='1'  OR oVar1S93(0)='1'  )then
          oVar2S30(0) <='1';
          else
          oVar2S30(0) <='0';
          end if;
        if(oVar1S94(0)='1'  )then
          oVar2S31(0) <='1';
          else
          oVar2S31(0) <='0';
          end if;
        if(oVar1S96(0)='1'  OR oVar1S97(0)='1'  OR oVar1S98(0)='1'  OR oVar1S99(0)='1'  )then
          oVar2S32(0) <='1';
          else
          oVar2S32(0) <='0';
          end if;
        if(oVar1S100(0)='1'  )then
          oVar2S33(0) <='1';
          else
          oVar2S33(0) <='0';
          end if;
        if(oVar1S101(0)='1'  OR oVar1S102(0)='1'  OR oVar1S103(0)='1'  OR oVar1S104(0)='1'  )then
          oVar2S34(0) <='1';
          else
          oVar2S34(0) <='0';
          end if;
        if(oVar1S106(0)='1'  OR oVar1S107(0)='1'  OR oVar1S108(0)='1'  OR oVar1S109(0)='1'  )then
          oVar2S36(0) <='1';
          else
          oVar2S36(0) <='0';
          end if;
        if(oVar1S110(0)='1'  )then
          oVar2S37(0) <='1';
          else
          oVar2S37(0) <='0';
          end if;
        if(oVar1S112(0)='1'  OR oVar1S113(0)='1'  OR oVar1S114(0)='1'  )then
          oVar2S38(0) <='1';
          else
          oVar2S38(0) <='0';
          end if;
        if(oVar1S115(0)='1'  OR oVar1S116(0)='1'  OR oVar1S117(0)='1'  OR oVar1S118(0)='1'  )then
          oVar2S39(0) <='1';
          else
          oVar2S39(0) <='0';
          end if;
        if(oVar1S120(0)='1'  OR oVar1S121(0)='1'  OR oVar1S122(0)='1'  )then
          oVar2S41(0) <='1';
          else
          oVar2S41(0) <='0';
          end if;
        if(oVar1S123(0)='1'  OR oVar1S124(0)='1'  OR oVar1S125(0)='1'  OR oVar1S126(0)='1'  )then
          oVar2S42(0) <='1';
          else
          oVar2S42(0) <='0';
          end if;
        if(oVar1S127(0)='1'  OR oVar1S128(0)='1'  OR oVar1S129(0)='1'  OR oVar1S130(0)='1'  )then
          oVar2S44(0) <='1';
          else
          oVar2S44(0) <='0';
          end if;
        if(oVar1S131(0)='1'  OR oVar1S132(0)='1'  OR oVar1S133(0)='1'  OR oVar1S134(0)='1'  )then
          oVar2S46(0) <='1';
          else
          oVar2S46(0) <='0';
          end if;
        if(oVar1S135(0)='1'  )then
          oVar2S47(0) <='1';
          else
          oVar2S47(0) <='0';
          end if;
        if(oVar1S136(0)='1'  OR oVar1S137(0)='1'  OR oVar1S138(0)='1'  OR oVar1S139(0)='1'  )then
          oVar2S48(0) <='1';
          else
          oVar2S48(0) <='0';
          end if;
        if(oVar1S140(0)='1'  OR oVar1S141(0)='1'  OR oVar1S142(0)='1'  OR oVar1S143(0)='1'  )then
          oVar2S50(0) <='1';
          else
          oVar2S50(0) <='0';
          end if;
        if(oVar1S144(0)='1'  OR oVar1S145(0)='1'  OR oVar1S146(0)='1'  OR oVar1S147(0)='1'  )then
          oVar2S51(0) <='1';
          else
          oVar2S51(0) <='0';
          end if;
        if(oVar1S149(0)='1'  OR oVar1S150(0)='1'  OR oVar1S151(0)='1'  OR oVar1S152(0)='1'  )then
          oVar2S53(0) <='1';
          else
          oVar2S53(0) <='0';
          end if;
        if(oVar1S153(0)='1'  OR oVar1S154(0)='1'  )then
          oVar2S54(0) <='1';
          else
          oVar2S54(0) <='0';
          end if;
        if(oVar1S155(0)='1'  OR oVar1S156(0)='1'  OR oVar1S157(0)='1'  OR oVar1S158(0)='1'  )then
          oVar2S55(0) <='1';
          else
          oVar2S55(0) <='0';
          end if;
        if(oVar1S159(0)='1'  OR oVar1S160(0)='1'  OR oVar1S161(0)='1'  )then
          oVar2S56(0) <='1';
          else
          oVar2S56(0) <='0';
          end if;
        if(oVar1S163(0)='1'  OR oVar1S164(0)='1'  OR oVar1S165(0)='1'  OR oVar1S166(0)='1'  )then
          oVar2S58(0) <='1';
          else
          oVar2S58(0) <='0';
          end if;
        if(oVar1S167(0)='1'  )then
          oVar2S59(0) <='1';
          else
          oVar2S59(0) <='0';
          end if;
        if(oVar1S169(0)='1'  OR oVar1S170(0)='1'  OR oVar1S171(0)='1'  OR oVar1S172(0)='1'  )then
          oVar2S60(0) <='1';
          else
          oVar2S60(0) <='0';
          end if;
        if(oVar1S173(0)='1'  )then
          oVar2S61(0) <='1';
          else
          oVar2S61(0) <='0';
          end if;
        if(oVar1S175(0)='1'  OR oVar1S176(0)='1'  OR oVar1S177(0)='1'  OR oVar1S178(0)='1'  )then
          oVar2S62(0) <='1';
          else
          oVar2S62(0) <='0';
          end if;
        if(oVar1S179(0)='1'  )then
          oVar2S63(0) <='1';
          else
          oVar2S63(0) <='0';
          end if;
        if(oVar1S180(0)='1'  OR oVar1S181(0)='1'  OR oVar1S182(0)='1'  OR oVar1S183(0)='1'  )then
          oVar2S64(0) <='1';
          else
          oVar2S64(0) <='0';
          end if;
        if(oVar1S184(0)='1'  OR oVar1S185(0)='1'  )then
          oVar2S65(0) <='1';
          else
          oVar2S65(0) <='0';
          end if;
        if(oVar1S186(0)='1'  OR oVar1S187(0)='1'  OR oVar1S188(0)='1'  OR oVar1S189(0)='1'  )then
          oVar2S66(0) <='1';
          else
          oVar2S66(0) <='0';
          end if;
        if(oVar1S190(0)='1'  )then
          oVar2S67(0) <='1';
          else
          oVar2S67(0) <='0';
          end if;
        if(oVar1S191(0)='1'  OR oVar1S192(0)='1'  OR oVar1S193(0)='1'  OR oVar1S194(0)='1'  )then
          oVar2S68(0) <='1';
          else
          oVar2S68(0) <='0';
          end if;
        if(oVar1S195(0)='1'  )then
          oVar2S69(0) <='1';
          else
          oVar2S69(0) <='0';
          end if;
        if(oVar1S196(0)='1'  OR oVar1S197(0)='1'  OR oVar1S198(0)='1'  OR oVar1S199(0)='1'  )then
          oVar2S70(0) <='1';
          else
          oVar2S70(0) <='0';
          end if;
        if(oVar1S200(0)='1'  OR oVar1S201(0)='1'  )then
          oVar2S71(0) <='1';
          else
          oVar2S71(0) <='0';
          end if;
        if(oVar1S202(0)='1'  OR oVar1S203(0)='1'  OR oVar1S204(0)='1'  OR oVar1S205(0)='1'  )then
          oVar2S72(0) <='1';
          else
          oVar2S72(0) <='0';
          end if;
        if(oVar1S206(0)='1'  OR oVar1S207(0)='1'  )then
          oVar2S73(0) <='1';
          else
          oVar2S73(0) <='0';
          end if;
        if(oVar1S208(0)='1'  OR oVar1S209(0)='1'  OR oVar1S210(0)='1'  OR oVar1S211(0)='1'  )then
          oVar2S74(0) <='1';
          else
          oVar2S74(0) <='0';
          end if;
        if(oVar1S212(0)='1'  )then
          oVar2S75(0) <='1';
          else
          oVar2S75(0) <='0';
          end if;
        if(oVar1S213(0)='1'  OR oVar1S214(0)='1'  OR oVar1S215(0)='1'  OR oVar1S216(0)='1'  )then
          oVar2S76(0) <='1';
          else
          oVar2S76(0) <='0';
          end if;
        if(oVar1S217(0)='1'  )then
          oVar2S77(0) <='1';
          else
          oVar2S77(0) <='0';
          end if;
        if(oVar1S218(0)='1'  OR oVar1S219(0)='1'  OR oVar1S220(0)='1'  OR oVar1S221(0)='1'  )then
          oVar2S78(0) <='1';
          else
          oVar2S78(0) <='0';
          end if;
        if(oVar1S222(0)='1'  )then
          oVar2S79(0) <='1';
          else
          oVar2S79(0) <='0';
          end if;
        if(oVar1S223(0)='1'  OR oVar1S224(0)='1'  OR oVar1S225(0)='1'  OR oVar1S226(0)='1'  )then
          oVar2S80(0) <='1';
          else
          oVar2S80(0) <='0';
          end if;
        if(oVar1S227(0)='1'  OR oVar1S228(0)='1'  )then
          oVar2S81(0) <='1';
          else
          oVar2S81(0) <='0';
          end if;
        if(oVar1S229(0)='1'  OR oVar1S230(0)='1'  OR oVar1S231(0)='1'  OR oVar1S232(0)='1'  )then
          oVar2S82(0) <='1';
          else
          oVar2S82(0) <='0';
          end if;
        if(oVar1S233(0)='1'  )then
          oVar2S83(0) <='1';
          else
          oVar2S83(0) <='0';
          end if;
        if(oVar1S235(0)='1'  OR oVar1S236(0)='1'  OR oVar1S237(0)='1'  OR oVar1S238(0)='1'  )then
          oVar2S84(0) <='1';
          else
          oVar2S84(0) <='0';
          end if;
        if(oVar1S239(0)='1'  OR oVar1S240(0)='1'  )then
          oVar2S85(0) <='1';
          else
          oVar2S85(0) <='0';
          end if;
        if(oVar1S241(0)='1'  OR oVar1S242(0)='1'  OR oVar1S243(0)='1'  OR oVar1S244(0)='1'  )then
          oVar2S86(0) <='1';
          else
          oVar2S86(0) <='0';
          end if;
        if(oVar1S245(0)='1'  )then
          oVar2S87(0) <='1';
          else
          oVar2S87(0) <='0';
          end if;
        if(oVar1S246(0)='1'  OR oVar1S247(0)='1'  OR oVar1S248(0)='1'  OR oVar1S249(0)='1'  )then
          oVar2S88(0) <='1';
          else
          oVar2S88(0) <='0';
          end if;
        if(oVar1S250(0)='1'  OR oVar1S251(0)='1'  )then
          oVar2S89(0) <='1';
          else
          oVar2S89(0) <='0';
          end if;
        if(oVar1S252(0)='1'  OR oVar1S253(0)='1'  OR oVar1S254(0)='1'  OR oVar1S255(0)='1'  )then
          oVar2S90(0) <='1';
          else
          oVar2S90(0) <='0';
          end if;
        if(oVar1S256(0)='1'  OR oVar1S257(0)='1'  )then
          oVar2S91(0) <='1';
          else
          oVar2S91(0) <='0';
          end if;
        if(oVar1S258(0)='1'  OR oVar1S259(0)='1'  OR oVar1S260(0)='1'  OR oVar1S261(0)='1'  )then
          oVar2S92(0) <='1';
          else
          oVar2S92(0) <='0';
          end if;
        if(oVar1S262(0)='1'  OR oVar1S263(0)='1'  )then
          oVar2S93(0) <='1';
          else
          oVar2S93(0) <='0';
          end if;
        if(oVar1S264(0)='1'  OR oVar1S265(0)='1'  OR oVar1S266(0)='1'  OR oVar1S267(0)='1'  )then
          oVar2S94(0) <='1';
          else
          oVar2S94(0) <='0';
          end if;
        if(oVar1S268(0)='1'  OR oVar1S269(0)='1'  )then
          oVar2S95(0) <='1';
          else
          oVar2S95(0) <='0';
          end if;
        if(oVar1S270(0)='1'  OR oVar1S271(0)='1'  OR oVar1S272(0)='1'  OR oVar1S273(0)='1'  )then
          oVar2S96(0) <='1';
          else
          oVar2S96(0) <='0';
          end if;
        if(oVar1S274(0)='1'  )then
          oVar2S97(0) <='1';
          else
          oVar2S97(0) <='0';
          end if;
        if(oVar1S275(0)='1'  OR oVar1S276(0)='1'  OR oVar1S277(0)='1'  OR oVar1S278(0)='1'  )then
          oVar2S98(0) <='1';
          else
          oVar2S98(0) <='0';
          end if;
        if(oVar1S279(0)='1'  OR oVar1S280(0)='1'  )then
          oVar2S99(0) <='1';
          else
          oVar2S99(0) <='0';
          end if;
        if(oVar1S281(0)='1'  OR oVar1S282(0)='1'  OR oVar1S283(0)='1'  OR oVar1S284(0)='1'  )then
          oVar2S100(0) <='1';
          else
          oVar2S100(0) <='0';
          end if;
        if(oVar1S285(0)='1'  )then
          oVar2S101(0) <='1';
          else
          oVar2S101(0) <='0';
          end if;
        if(oVar1S286(0)='1'  OR oVar1S287(0)='1'  OR oVar1S288(0)='1'  OR oVar1S289(0)='1'  )then
          oVar2S102(0) <='1';
          else
          oVar2S102(0) <='0';
          end if;
        if(oVar1S290(0)='1'  OR oVar1S291(0)='1'  )then
          oVar2S103(0) <='1';
          else
          oVar2S103(0) <='0';
          end if;
        if(oVar1S292(0)='1'  OR oVar1S293(0)='1'  OR oVar1S294(0)='1'  OR oVar1S295(0)='1'  )then
          oVar2S104(0) <='1';
          else
          oVar2S104(0) <='0';
          end if;
        if(oVar1S296(0)='1'  OR oVar1S297(0)='1'  )then
          oVar2S105(0) <='1';
          else
          oVar2S105(0) <='0';
          end if;
        if(oVar1S298(0)='1'  OR oVar1S299(0)='1'  OR oVar1S300(0)='1'  OR oVar1S301(0)='1'  )then
          oVar2S106(0) <='1';
          else
          oVar2S106(0) <='0';
          end if;
        if(oVar1S302(0)='1'  )then
          oVar2S107(0) <='1';
          else
          oVar2S107(0) <='0';
          end if;
        if(oVar1S303(0)='1'  OR oVar1S304(0)='1'  OR oVar1S305(0)='1'  OR oVar1S306(0)='1'  )then
          oVar2S108(0) <='1';
          else
          oVar2S108(0) <='0';
          end if;
        if(oVar1S307(0)='1'  OR oVar1S308(0)='1'  OR oVar1S309(0)='1'  )then
          oVar2S109(0) <='1';
          else
          oVar2S109(0) <='0';
          end if;
        if(oVar1S310(0)='1'  OR oVar1S311(0)='1'  OR oVar1S312(0)='1'  OR oVar1S313(0)='1'  )then
          oVar2S110(0) <='1';
          else
          oVar2S110(0) <='0';
          end if;
        if(oVar1S314(0)='1'  OR oVar1S315(0)='1'  OR oVar1S316(0)='1'  )then
          oVar2S111(0) <='1';
          else
          oVar2S111(0) <='0';
          end if;
        if(oVar1S317(0)='1'  OR oVar1S318(0)='1'  OR oVar1S319(0)='1'  OR oVar1S320(0)='1'  )then
          oVar2S112(0) <='1';
          else
          oVar2S112(0) <='0';
          end if;
        if(oVar1S321(0)='1'  OR oVar1S322(0)='1'  )then
          oVar2S113(0) <='1';
          else
          oVar2S113(0) <='0';
          end if;
        if(oVar1S323(0)='1'  OR oVar1S324(0)='1'  OR oVar1S325(0)='1'  OR oVar1S326(0)='1'  )then
          oVar2S114(0) <='1';
          else
          oVar2S114(0) <='0';
          end if;
        if(oVar1S327(0)='1'  OR oVar1S328(0)='1'  )then
          oVar2S115(0) <='1';
          else
          oVar2S115(0) <='0';
          end if;
        if(oVar1S329(0)='1'  OR oVar1S330(0)='1'  OR oVar1S331(0)='1'  OR oVar1S332(0)='1'  )then
          oVar2S116(0) <='1';
          else
          oVar2S116(0) <='0';
          end if;
        if(oVar1S333(0)='1'  OR oVar1S334(0)='1'  )then
          oVar2S117(0) <='1';
          else
          oVar2S117(0) <='0';
          end if;
        if(oVar1S335(0)='1'  OR oVar1S336(0)='1'  OR oVar1S337(0)='1'  OR oVar1S338(0)='1'  )then
          oVar2S118(0) <='1';
          else
          oVar2S118(0) <='0';
          end if;
        if(oVar1S339(0)='1'  OR oVar1S340(0)='1'  )then
          oVar2S119(0) <='1';
          else
          oVar2S119(0) <='0';
          end if;
        if(oVar1S341(0)='1'  OR oVar1S342(0)='1'  OR oVar1S343(0)='1'  OR oVar1S344(0)='1'  )then
          oVar2S120(0) <='1';
          else
          oVar2S120(0) <='0';
          end if;
        if(oVar1S345(0)='1'  OR oVar1S346(0)='1'  )then
          oVar2S121(0) <='1';
          else
          oVar2S121(0) <='0';
          end if;
        if(oVar1S347(0)='1'  OR oVar1S348(0)='1'  OR oVar1S349(0)='1'  OR oVar1S350(0)='1'  )then
          oVar2S122(0) <='1';
          else
          oVar2S122(0) <='0';
          end if;
        if(oVar1S351(0)='1'  OR oVar1S352(0)='1'  )then
          oVar2S123(0) <='1';
          else
          oVar2S123(0) <='0';
          end if;
        if(oVar1S353(0)='1'  OR oVar1S354(0)='1'  OR oVar1S355(0)='1'  OR oVar1S356(0)='1'  )then
          oVar2S124(0) <='1';
          else
          oVar2S124(0) <='0';
          end if;
        if(oVar1S357(0)='1'  OR oVar1S358(0)='1'  OR oVar1S359(0)='1'  OR oVar1S360(0)='1'  )then
          oVar2S126(0) <='1';
          else
          oVar2S126(0) <='0';
          end if;
        if(oVar1S361(0)='1'  )then
          oVar2S127(0) <='1';
          else
          oVar2S127(0) <='0';
          end if;
        if(oVar1S362(0)='1'  OR oVar1S363(0)='1'  OR oVar1S364(0)='1'  OR oVar1S365(0)='1'  )then
          oVar2S128(0) <='1';
          else
          oVar2S128(0) <='0';
          end if;
        if(oVar1S366(0)='1'  OR oVar1S367(0)='1'  )then
          oVar2S129(0) <='1';
          else
          oVar2S129(0) <='0';
          end if;
        if(oVar1S368(0)='1'  OR oVar1S369(0)='1'  OR oVar1S370(0)='1'  OR oVar1S371(0)='1'  )then
          oVar2S130(0) <='1';
          else
          oVar2S130(0) <='0';
          end if;
        if(oVar1S372(0)='1'  OR oVar1S373(0)='1'  )then
          oVar2S131(0) <='1';
          else
          oVar2S131(0) <='0';
          end if;
        if(oVar1S374(0)='1'  OR oVar1S375(0)='1'  OR oVar1S376(0)='1'  OR oVar1S377(0)='1'  )then
          oVar2S132(0) <='1';
          else
          oVar2S132(0) <='0';
          end if;
        if(oVar1S378(0)='1'  OR oVar1S379(0)='1'  OR oVar1S380(0)='1'  OR oVar1S381(0)='1'  )then
          oVar2S134(0) <='1';
          else
          oVar2S134(0) <='0';
          end if;
        if(oVar1S383(0)='1'  OR oVar1S384(0)='1'  OR oVar1S385(0)='1'  OR oVar1S386(0)='1'  )then
          oVar2S136(0) <='1';
          else
          oVar2S136(0) <='0';
          end if;
        if(oVar1S387(0)='1'  )then
          oVar2S137(0) <='1';
          else
          oVar2S137(0) <='0';
          end if;
        if(oVar1S388(0)='1'  OR oVar1S389(0)='1'  OR oVar1S390(0)='1'  OR oVar1S391(0)='1'  )then
          oVar2S138(0) <='1';
          else
          oVar2S138(0) <='0';
          end if;
        if(oVar1S392(0)='1'  OR oVar1S393(0)='1'  OR oVar1S394(0)='1'  OR oVar1S395(0)='1'  )then
          oVar2S140(0) <='1';
          else
          oVar2S140(0) <='0';
          end if;
        if(oVar1S397(0)='1'  OR oVar1S398(0)='1'  OR oVar1S399(0)='1'  OR oVar1S400(0)='1'  )then
          oVar2S142(0) <='1';
          else
          oVar2S142(0) <='0';
          end if;
        if(oVar1S401(0)='1'  OR oVar1S402(0)='1'  OR oVar1S403(0)='1'  OR oVar1S404(0)='1'  )then
          oVar2S144(0) <='1';
          else
          oVar2S144(0) <='0';
          end if;
        if(oVar1S405(0)='1'  OR oVar1S406(0)='1'  OR oVar1S407(0)='1'  OR oVar1S408(0)='1'  )then
          oVar2S146(0) <='1';
          else
          oVar2S146(0) <='0';
          end if;
        if(oVar1S409(0)='1'  OR oVar1S410(0)='1'  OR oVar1S411(0)='1'  OR oVar1S412(0)='1'  )then
          oVar2S148(0) <='1';
          else
          oVar2S148(0) <='0';
          end if;
        if(oVar1S413(0)='1'  OR oVar1S414(0)='1'  )then
          oVar2S149(0) <='1';
          else
          oVar2S149(0) <='0';
          end if;
        if(oVar1S415(0)='1'  OR oVar1S416(0)='1'  OR oVar1S417(0)='1'  OR oVar1S418(0)='1'  )then
          oVar2S150(0) <='1';
          else
          oVar2S150(0) <='0';
          end if;
        if(oVar1S419(0)='1'  OR oVar1S420(0)='1'  )then
          oVar2S151(0) <='1';
          else
          oVar2S151(0) <='0';
          end if;
        if(oVar1S421(0)='1'  OR oVar1S422(0)='1'  OR oVar1S423(0)='1'  OR oVar1S424(0)='1'  )then
          oVar2S152(0) <='1';
          else
          oVar2S152(0) <='0';
          end if;
        if(oVar1S425(0)='1'  )then
          oVar2S153(0) <='1';
          else
          oVar2S153(0) <='0';
          end if;
        if(oVar1S427(0)='1'  OR oVar1S428(0)='1'  OR oVar1S429(0)='1'  OR oVar1S430(0)='1'  )then
          oVar2S154(0) <='1';
          else
          oVar2S154(0) <='0';
          end if;
        if(oVar1S431(0)='1'  )then
          oVar2S155(0) <='1';
          else
          oVar2S155(0) <='0';
          end if;
        if(oVar1S433(0)='1'  OR oVar1S434(0)='1'  OR oVar1S435(0)='1'  )then
          oVar2S156(0) <='1';
          else
          oVar2S156(0) <='0';
          end if;
        if(oVar1S436(0)='1'  OR oVar1S437(0)='1'  OR oVar1S438(0)='1'  OR oVar1S439(0)='1'  )then
          oVar2S157(0) <='1';
          else
          oVar2S157(0) <='0';
          end if;
        if(oVar1S440(0)='1'  OR oVar1S441(0)='1'  OR oVar1S442(0)='1'  OR oVar1S443(0)='1'  )then
          oVar2S159(0) <='1';
          else
          oVar2S159(0) <='0';
          end if;
        if(oVar1S444(0)='1'  OR oVar1S445(0)='1'  OR oVar1S446(0)='1'  )then
          oVar2S160(0) <='1';
          else
          oVar2S160(0) <='0';
          end if;
        if(oVar1S447(0)='1'  OR oVar1S448(0)='1'  OR oVar1S449(0)='1'  OR oVar1S450(0)='1'  )then
          oVar2S161(0) <='1';
          else
          oVar2S161(0) <='0';
          end if;
        if(oVar1S451(0)='1'  OR oVar1S452(0)='1'  OR oVar1S453(0)='1'  OR oVar1S454(0)='1'  )then
          oVar2S162(0) <='1';
          else
          oVar2S162(0) <='0';
          end if;
        if(oVar1S455(0)='1'  OR oVar1S456(0)='1'  OR oVar1S457(0)='1'  OR oVar1S458(0)='1'  )then
          oVar2S164(0) <='1';
          else
          oVar2S164(0) <='0';
          end if;
        if(oVar1S459(0)='1'  )then
          oVar2S165(0) <='1';
          else
          oVar2S165(0) <='0';
          end if;
        if(oVar1S461(0)='1'  OR oVar1S462(0)='1'  OR oVar1S463(0)='1'  OR oVar1S464(0)='1'  )then
          oVar2S166(0) <='1';
          else
          oVar2S166(0) <='0';
          end if;
        if(oVar1S465(0)='1'  OR oVar1S466(0)='1'  )then
          oVar2S167(0) <='1';
          else
          oVar2S167(0) <='0';
          end if;
        if(oVar1S467(0)='1'  OR oVar1S468(0)='1'  OR oVar1S469(0)='1'  OR oVar1S470(0)='1'  )then
          oVar2S168(0) <='1';
          else
          oVar2S168(0) <='0';
          end if;
        if(oVar1S471(0)='1'  OR oVar1S472(0)='1'  )then
          oVar2S169(0) <='1';
          else
          oVar2S169(0) <='0';
          end if;
        if(oVar1S473(0)='1'  OR oVar1S474(0)='1'  OR oVar1S475(0)='1'  OR oVar1S476(0)='1'  )then
          oVar2S170(0) <='1';
          else
          oVar2S170(0) <='0';
          end if;
        if(oVar1S477(0)='1'  OR oVar1S478(0)='1'  OR oVar1S479(0)='1'  )then
          oVar2S171(0) <='1';
          else
          oVar2S171(0) <='0';
          end if;
        if(oVar1S480(0)='1'  OR oVar1S481(0)='1'  OR oVar1S482(0)='1'  OR oVar1S483(0)='1'  )then
          oVar2S172(0) <='1';
          else
          oVar2S172(0) <='0';
          end if;
        if(oVar1S484(0)='1'  )then
          oVar2S173(0) <='1';
          else
          oVar2S173(0) <='0';
          end if;
        if(oVar1S486(0)='1'  OR oVar1S487(0)='1'  OR oVar1S488(0)='1'  OR oVar1S489(0)='1'  )then
          oVar2S174(0) <='1';
          else
          oVar2S174(0) <='0';
          end if;
        if(oVar1S490(0)='1'  OR oVar1S491(0)='1'  OR oVar1S492(0)='1'  )then
          oVar2S175(0) <='1';
          else
          oVar2S175(0) <='0';
          end if;
        if(oVar1S493(0)='1'  OR oVar1S494(0)='1'  OR oVar1S495(0)='1'  OR oVar1S496(0)='1'  )then
          oVar2S176(0) <='1';
          else
          oVar2S176(0) <='0';
          end if;
        if(oVar1S497(0)='1'  OR oVar1S498(0)='1'  )then
          oVar2S177(0) <='1';
          else
          oVar2S177(0) <='0';
          end if;
        if(oVar1S499(0)='1'  OR oVar1S500(0)='1'  OR oVar1S501(0)='1'  OR oVar1S502(0)='1'  )then
          oVar2S178(0) <='1';
          else
          oVar2S178(0) <='0';
          end if;
        if(oVar1S503(0)='1'  OR oVar1S504(0)='1'  )then
          oVar2S179(0) <='1';
          else
          oVar2S179(0) <='0';
          end if;
        if(oVar1S505(0)='1'  OR oVar1S506(0)='1'  OR oVar1S507(0)='1'  OR oVar1S508(0)='1'  )then
          oVar2S180(0) <='1';
          else
          oVar2S180(0) <='0';
          end if;
        if(oVar1S509(0)='1'  )then
          oVar2S181(0) <='1';
          else
          oVar2S181(0) <='0';
          end if;
        if(oVar1S511(0)='1'  OR oVar1S512(0)='1'  OR oVar1S513(0)='1'  OR oVar1S514(0)='1'  )then
          oVar2S182(0) <='1';
          else
          oVar2S182(0) <='0';
          end if;
        if(oVar1S516(0)='1'  OR oVar1S517(0)='1'  OR oVar1S518(0)='1'  OR oVar1S519(0)='1'  )then
          oVar2S184(0) <='1';
          else
          oVar2S184(0) <='0';
          end if;
        if(oVar1S520(0)='1'  OR oVar1S521(0)='1'  OR oVar1S522(0)='1'  )then
          oVar2S185(0) <='1';
          else
          oVar2S185(0) <='0';
          end if;
        if(oVar1S523(0)='1'  OR oVar1S524(0)='1'  OR oVar1S525(0)='1'  OR oVar1S526(0)='1'  )then
          oVar2S186(0) <='1';
          else
          oVar2S186(0) <='0';
          end if;
        if(oVar1S527(0)='1'  OR oVar1S528(0)='1'  )then
          oVar2S187(0) <='1';
          else
          oVar2S187(0) <='0';
          end if;
        if(oVar1S529(0)='1'  OR oVar1S530(0)='1'  OR oVar1S531(0)='1'  OR oVar1S532(0)='1'  )then
          oVar2S188(0) <='1';
          else
          oVar2S188(0) <='0';
          end if;
        if(oVar1S533(0)='1'  OR oVar1S534(0)='1'  )then
          oVar2S189(0) <='1';
          else
          oVar2S189(0) <='0';
          end if;
        if(oVar1S536(0)='1'  OR oVar1S537(0)='1'  OR oVar1S538(0)='1'  OR oVar1S539(0)='1'  )then
          oVar2S190(0) <='1';
          else
          oVar2S190(0) <='0';
          end if;
        if(oVar1S540(0)='1'  OR oVar1S541(0)='1'  OR oVar1S542(0)='1'  )then
          oVar2S191(0) <='1';
          else
          oVar2S191(0) <='0';
          end if;
        if(oVar1S543(0)='1'  OR oVar1S544(0)='1'  OR oVar1S545(0)='1'  OR oVar1S546(0)='1'  )then
          oVar2S192(0) <='1';
          else
          oVar2S192(0) <='0';
          end if;
        if(oVar1S547(0)='1'  OR oVar1S548(0)='1'  OR oVar1S549(0)='1'  )then
          oVar2S193(0) <='1';
          else
          oVar2S193(0) <='0';
          end if;
        if(oVar1S550(0)='1'  OR oVar1S551(0)='1'  OR oVar1S552(0)='1'  OR oVar1S553(0)='1'  )then
          oVar2S194(0) <='1';
          else
          oVar2S194(0) <='0';
          end if;
        if(oVar1S554(0)='1'  OR oVar1S555(0)='1'  OR oVar1S556(0)='1'  OR oVar1S557(0)='1'  )then
          oVar2S196(0) <='1';
          else
          oVar2S196(0) <='0';
          end if;
        if(oVar1S558(0)='1'  )then
          oVar2S197(0) <='1';
          else
          oVar2S197(0) <='0';
          end if;
        if(oVar1S559(0)='1'  OR oVar1S560(0)='1'  OR oVar1S561(0)='1'  OR oVar1S562(0)='1'  )then
          oVar2S198(0) <='1';
          else
          oVar2S198(0) <='0';
          end if;
        if(oVar1S563(0)='1'  )then
          oVar2S199(0) <='1';
          else
          oVar2S199(0) <='0';
          end if;
        if(oVar1S565(0)='1'  OR oVar1S566(0)='1'  OR oVar1S567(0)='1'  OR oVar1S568(0)='1'  )then
          oVar2S200(0) <='1';
          else
          oVar2S200(0) <='0';
          end if;
        if(oVar1S569(0)='1'  )then
          oVar2S201(0) <='1';
          else
          oVar2S201(0) <='0';
          end if;
        if(oVar1S571(0)='1'  OR oVar1S572(0)='1'  OR oVar1S573(0)='1'  OR oVar1S574(0)='1'  )then
          oVar2S202(0) <='1';
          else
          oVar2S202(0) <='0';
          end if;
        if(oVar1S575(0)='1'  OR oVar1S576(0)='1'  OR oVar1S577(0)='1'  OR oVar1S578(0)='1'  )then
          oVar2S204(0) <='1';
          else
          oVar2S204(0) <='0';
          end if;
        if(oVar1S579(0)='1'  OR oVar1S580(0)='1'  )then
          oVar2S205(0) <='1';
          else
          oVar2S205(0) <='0';
          end if;
        if(oVar1S581(0)='1'  OR oVar1S582(0)='1'  OR oVar1S583(0)='1'  OR oVar1S584(0)='1'  )then
          oVar2S206(0) <='1';
          else
          oVar2S206(0) <='0';
          end if;
        if(oVar1S585(0)='1'  OR oVar1S586(0)='1'  OR oVar1S587(0)='1'  OR oVar1S588(0)='1'  )then
          oVar2S208(0) <='1';
          else
          oVar2S208(0) <='0';
          end if;
        if(oVar1S589(0)='1'  )then
          oVar2S209(0) <='1';
          else
          oVar2S209(0) <='0';
          end if;
        if(oVar1S591(0)='1'  OR oVar1S592(0)='1'  OR oVar1S593(0)='1'  )then
          oVar2S210(0) <='1';
          else
          oVar2S210(0) <='0';
          end if;
        if(oVar1S595(0)='1'  OR oVar1S596(0)='1'  OR oVar1S597(0)='1'  OR oVar1S598(0)='1'  )then
          oVar2S212(0) <='1';
          else
          oVar2S212(0) <='0';
          end if;
        if(oVar1S599(0)='1'  OR oVar1S600(0)='1'  OR oVar1S601(0)='1'  )then
          oVar2S214(0) <='1';
          else
          oVar2S214(0) <='0';
          end if;
        if(oVar1S603(0)='1'  OR oVar1S604(0)='1'  OR oVar1S605(0)='1'  OR oVar1S606(0)='1'  )then
          oVar2S216(0) <='1';
          else
          oVar2S216(0) <='0';
          end if;
        if(oVar1S607(0)='1'  )then
          oVar2S217(0) <='1';
          else
          oVar2S217(0) <='0';
          end if;
        if(oVar1S608(0)='1'  OR oVar1S609(0)='1'  OR oVar1S610(0)='1'  )then
          oVar2S218(0) <='1';
          else
          oVar2S218(0) <='0';
          end if;
        if(oVar1S611(0)='1'  OR oVar1S612(0)='1'  OR oVar1S613(0)='1'  )then
          oVar2S219(0) <='1';
          else
          oVar2S219(0) <='0';
          end if;
        if(oVar1S615(0)='1'  OR oVar1S616(0)='1'  OR oVar1S617(0)='1'  OR oVar1S618(0)='1'  )then
          oVar2S221(0) <='1';
          else
          oVar2S221(0) <='0';
          end if;
        if(oVar1S619(0)='1'  OR oVar1S620(0)='1'  OR oVar1S621(0)='1'  )then
          oVar2S223(0) <='1';
          else
          oVar2S223(0) <='0';
          end if;
        if(oVar1S623(0)='1'  OR oVar1S624(0)='1'  OR oVar1S625(0)='1'  )then
          oVar2S225(0) <='1';
          else
          oVar2S225(0) <='0';
          end if;
        if(oVar1S627(0)='1'  OR oVar1S628(0)='1'  OR oVar1S629(0)='1'  OR oVar1S630(0)='1'  )then
          oVar2S227(0) <='1';
          else
          oVar2S227(0) <='0';
          end if;
        if(oVar1S631(0)='1'  )then
          oVar2S228(0) <='1';
          else
          oVar2S228(0) <='0';
          end if;
        if(oVar1S632(0)='1'  OR oVar1S633(0)='1'  OR oVar1S634(0)='1'  OR oVar1S635(0)='1'  )then
          oVar2S229(0) <='1';
          else
          oVar2S229(0) <='0';
          end if;
        if(oVar1S636(0)='1'  OR oVar1S637(0)='1'  OR oVar1S638(0)='1'  OR oVar1S639(0)='1'  )then
          oVar2S231(0) <='1';
          else
          oVar2S231(0) <='0';
          end if;
        if(oVar1S640(0)='1'  )then
          oVar2S232(0) <='1';
          else
          oVar2S232(0) <='0';
          end if;
        if(oVar1S641(0)='1'  OR oVar1S642(0)='1'  OR oVar1S643(0)='1'  OR oVar1S644(0)='1'  )then
          oVar2S233(0) <='1';
          else
          oVar2S233(0) <='0';
          end if;
        if(oVar1S645(0)='1'  OR oVar1S646(0)='1'  OR oVar1S647(0)='1'  )then
          oVar2S235(0) <='1';
          else
          oVar2S235(0) <='0';
          end if;
        if(oVar1S649(0)='1'  OR oVar1S650(0)='1'  OR oVar1S651(0)='1'  )then
          oVar2S237(0) <='1';
          else
          oVar2S237(0) <='0';
          end if;
        if(oVar1S652(0)='1'  OR oVar1S653(0)='1'  OR oVar1S654(0)='1'  )then
          oVar2S238(0) <='1';
          else
          oVar2S238(0) <='0';
          end if;
        if(oVar1S655(0)='1'  OR oVar1S656(0)='1'  OR oVar1S657(0)='1'  OR oVar1S658(0)='1'  )then
          oVar2S239(0) <='1';
          else
          oVar2S239(0) <='0';
          end if;
        if(oVar1S659(0)='1'  OR oVar1S660(0)='1'  OR oVar1S661(0)='1'  OR oVar1S662(0)='1'  )then
          oVar2S241(0) <='1';
          else
          oVar2S241(0) <='0';
          end if;
        if(oVar1S663(0)='1'  OR oVar1S664(0)='1'  OR oVar1S665(0)='1'  OR oVar1S666(0)='1'  )then
          oVar2S243(0) <='1';
          else
          oVar2S243(0) <='0';
          end if;
        if(oVar1S668(0)='1'  OR oVar1S669(0)='1'  OR oVar1S670(0)='1'  OR oVar1S671(0)='1'  )then
          oVar2S245(0) <='1';
          else
          oVar2S245(0) <='0';
          end if;
        if(oVar1S672(0)='1'  OR oVar1S673(0)='1'  )then
          oVar2S246(0) <='1';
          else
          oVar2S246(0) <='0';
          end if;
        if(oVar1S675(0)='1'  OR oVar1S676(0)='1'  OR oVar1S677(0)='1'  OR oVar1S678(0)='1'  )then
          oVar2S247(0) <='1';
          else
          oVar2S247(0) <='0';
          end if;
        if(oVar1S679(0)='1'  OR oVar1S680(0)='1'  )then
          oVar2S248(0) <='1';
          else
          oVar2S248(0) <='0';
          end if;
        if(oVar1S681(0)='1'  OR oVar1S682(0)='1'  OR oVar1S683(0)='1'  OR oVar1S684(0)='1'  )then
          oVar2S249(0) <='1';
          else
          oVar2S249(0) <='0';
          end if;
        if(oVar1S685(0)='1'  OR oVar1S686(0)='1'  OR oVar1S687(0)='1'  )then
          oVar2S250(0) <='1';
          else
          oVar2S250(0) <='0';
          end if;
        if(oVar1S688(0)='1'  OR oVar1S689(0)='1'  OR oVar1S690(0)='1'  OR oVar1S691(0)='1'  )then
          oVar2S251(0) <='1';
          else
          oVar2S251(0) <='0';
          end if;
        if(oVar1S692(0)='1'  OR oVar1S693(0)='1'  OR oVar1S694(0)='1'  OR oVar1S695(0)='1'  )then
          oVar2S252(0) <='1';
          else
          oVar2S252(0) <='0';
          end if;
 end if;
end process;
lookuptable_LV5 : process(c1)
begin
 if c1'event and c1='1' then
        if(oVar2S106(0)='1' OR oVar2S107(0)='1' )then
          ADDM4K3S8(7)<='1';
          else
          ADDM4K3S8(7)<='0';
          end if;
        if(oVar2S128(0)='1' OR oVar2S129(0)='1' )then
          ADDM4K3S8(6)<='1';
          else
          ADDM4K3S8(6)<='0';
          end if;
        if(oVar2S122(0)='1' OR oVar2S123(0)='1' )then
          ADDM4K3S8(5)<='1';
          else
          ADDM4K3S8(5)<='0';
          end if;
        if(oVar2S116(0)='1' OR oVar2S117(0)='1' )then
          ADDM4K3S8(4)<='1';
          else
          ADDM4K3S8(4)<='0';
          end if;
        if(oVar2S86(0)='1' OR oVar2S87(0)='1' )then
          ADDM4K3S8(3)<='1';
          else
          ADDM4K3S8(3)<='0';
          end if;
        if(oVar2S104(0)='1' OR oVar2S105(0)='1' )then
          ADDM4K3S8(2)<='1';
          else
          ADDM4K3S8(2)<='0';
          end if;
        if(oVar2S170(0)='1' OR oVar2S171(0)='1' )then
          ADDM4K3S8(1)<='1';
          else
          ADDM4K3S8(1)<='0';
          end if;
        if(oVar2S251(0)='1' OR oVar2S252(0)='1' )then
          ADDM4K3S8(0)<='1';
          else
          ADDM4K3S8(0)<='0';
          end if;
        if(oVar2S118(0)='1' OR oVar2S119(0)='1' )then
          ADDM4K3S9(7)<='1';
          else
          ADDM4K3S9(7)<='0';
          end if;
        if(oVar2S94(0)='1' OR oVar2S95(0)='1' )then
          ADDM4K3S9(6)<='1';
          else
          ADDM4K3S9(6)<='0';
          end if;
        if(oVar1S112(0)='1' OR oVar1S113(0)='1' OR oVar1S114(0)='1' )then
          ADDM4K3S9(5)<='1';
          else
          ADDM4K3S9(5)<='0';
          end if;
        if(oVar2S102(0)='1' OR oVar2S103(0)='1' )then
          ADDM4K3S9(4)<='1';
          else
          ADDM4K3S9(4)<='0';
          end if;
        if(oVar2S114(0)='1' OR oVar2S115(0)='1' )then
          ADDM4K3S9(3)<='1';
          else
          ADDM4K3S9(3)<='0';
          end if;
        if(oVar2S168(0)='1' OR oVar2S169(0)='1' )then
          ADDM4K3S9(2)<='1';
          else
          ADDM4K3S9(2)<='0';
          end if;
        if(oVar2S48(0)='1' )then
          ADDM4K3S9(1)<='1';
          else
          ADDM4K3S9(1)<='0';
          end if;
        if(oVar2S76(0)='1' OR oVar2S77(0)='1' )then
          ADDM4K3S9(0)<='1';
          else
          ADDM4K3S9(0)<='0';
          end if;
        if(oVar2S90(0)='1' OR oVar2S91(0)='1' )then
          ADDM4K3S12(7)<='1';
          else
          ADDM4K3S12(7)<='0';
          end if;
        if(oVar2S60(0)='1' OR oVar2S61(0)='1' )then
          ADDM4K3S12(6)<='1';
          else
          ADDM4K3S12(6)<='0';
          end if;
        if(oVar2S68(0)='1' OR oVar2S69(0)='1' )then
          ADDM4K3S12(5)<='1';
          else
          ADDM4K3S12(5)<='0';
          end if;
        if(oVar2S44(0)='1' )then
          ADDM4K3S12(4)<='1';
          else
          ADDM4K3S12(4)<='0';
          end if;
        if(oVar2S88(0)='1' OR oVar2S89(0)='1' )then
          ADDM4K3S12(3)<='1';
          else
          ADDM4K3S12(3)<='0';
          end if;
        if(oVar2S62(0)='1' OR oVar2S63(0)='1' )then
          ADDM4K3S12(2)<='1';
          else
          ADDM4K3S12(2)<='0';
          end if;
        if(oVar2S72(0)='1' OR oVar2S73(0)='1' )then
          ADDM4K3S12(1)<='1';
          else
          ADDM4K3S12(1)<='0';
          end if;
        if(oVar2S66(0)='1' OR oVar2S67(0)='1' )then
          ADDM4K3S12(0)<='1';
          else
          ADDM4K3S12(0)<='0';
          end if;
        if(oVar2S34(0)='1' )then
          ADDM4K3S13(7)<='1';
          else
          ADDM4K3S13(7)<='0';
          end if;
        if(oVar2S70(0)='1' OR oVar2S71(0)='1' )then
          ADDM4K3S13(6)<='1';
          else
          ADDM4K3S13(6)<='0';
          end if;
        if(oVar2S28(0)='1' OR oVar2S29(0)='1' )then
          ADDM4K3S13(5)<='1';
          else
          ADDM4K3S13(5)<='0';
          end if;
        if(oVar2S64(0)='1' OR oVar2S65(0)='1' )then
          ADDM4K3S13(4)<='1';
          else
          ADDM4K3S13(4)<='0';
          end if;
        if(oVar2S58(0)='1' OR oVar2S59(0)='1' )then
          ADDM4K3S13(3)<='1';
          else
          ADDM4K3S13(3)<='0';
          end if;
        if(oVar2S32(0)='1' OR oVar2S33(0)='1' )then
          ADDM4K3S13(2)<='1';
          else
          ADDM4K3S13(2)<='0';
          end if;
        if(oVar2S55(0)='1' OR oVar2S56(0)='1' )then
          ADDM4K3S13(1)<='1';
          else
          ADDM4K3S13(1)<='0';
          end if;
        if(oVar2S50(0)='1' OR oVar2S51(0)='1' )then
          ADDM4K3S13(0)<='1';
          else
          ADDM4K3S13(0)<='0';
          end if;
        if(oVar2S96(0)='1' OR oVar2S97(0)='1' )then
          ADDM4K3S10(7)<='1';
          else
          ADDM4K3S10(7)<='0';
          end if;
        if(oVar2S98(0)='1' OR oVar2S99(0)='1' )then
          ADDM4K3S10(6)<='1';
          else
          ADDM4K3S10(6)<='0';
          end if;
        if(oVar1S120(0)='1' OR oVar1S121(0)='1' OR oVar1S122(0)='1' )then
          ADDM4K3S10(5)<='1';
          else
          ADDM4K3S10(5)<='0';
          end if;
        if(oVar2S161(0)='1' OR oVar2S162(0)='1' )then
          ADDM4K3S10(4)<='1';
          else
          ADDM4K3S10(4)<='0';
          end if;
        if(oVar2S82(0)='1' OR oVar2S83(0)='1' )then
          ADDM4K3S10(3)<='1';
          else
          ADDM4K3S10(3)<='0';
          end if;
        if(oVar2S110(0)='1' OR oVar2S111(0)='1' )then
          ADDM4K3S10(2)<='1';
          else
          ADDM4K3S10(2)<='0';
          end if;
        if(oVar2S120(0)='1' OR oVar2S121(0)='1' )then
          ADDM4K3S10(1)<='1';
          else
          ADDM4K3S10(1)<='0';
          end if;
        if(oVar2S42(0)='1' )then
          ADDM4K3S10(0)<='1';
          else
          ADDM4K3S10(0)<='0';
          end if;
        if(oVar2S78(0)='1' OR oVar2S79(0)='1' )then
          ADDM4K3S11(7)<='1';
          else
          ADDM4K3S11(7)<='0';
          end if;
        if(oVar2S39(0)='1' )then
          ADDM4K3S11(6)<='1';
          else
          ADDM4K3S11(6)<='0';
          end if;
        if(oVar2S84(0)='1' OR oVar2S85(0)='1' )then
          ADDM4K3S11(5)<='1';
          else
          ADDM4K3S11(5)<='0';
          end if;
        if(oVar2S74(0)='1' OR oVar2S75(0)='1' )then
          ADDM4K3S11(4)<='1';
          else
          ADDM4K3S11(4)<='0';
          end if;
        if(oVar2S108(0)='1' OR oVar2S109(0)='1' )then
          ADDM4K3S11(3)<='1';
          else
          ADDM4K3S11(3)<='0';
          end if;
        if(oVar2S100(0)='1' OR oVar2S101(0)='1' )then
          ADDM4K3S11(2)<='1';
          else
          ADDM4K3S11(2)<='0';
          end if;
        if(oVar2S46(0)='1' OR oVar2S47(0)='1' )then
          ADDM4K3S11(1)<='1';
          else
          ADDM4K3S11(1)<='0';
          end if;
        if(oVar2S36(0)='1' OR oVar2S37(0)='1' )then
          ADDM4K3S11(0)<='1';
          else
          ADDM4K3S11(0)<='0';
          end if;
        if(oVar2S53(0)='1' OR oVar2S54(0)='1' )then
          ADDM4K3S14(7)<='1';
          else
          ADDM4K3S14(7)<='0';
          end if;
        if(oVar2S20(0)='1' OR oVar2S21(0)='1' )then
          ADDM4K3S14(6)<='1';
          else
          ADDM4K3S14(6)<='0';
          end if;
        if(oVar2S30(0)='1' OR oVar2S31(0)='1' )then
          ADDM4K3S14(5)<='1';
          else
          ADDM4K3S14(5)<='0';
          end if;
        if(oVar2S26(0)='1' OR oVar2S27(0)='1' )then
          ADDM4K3S14(4)<='1';
          else
          ADDM4K3S14(4)<='0';
          end if;
        if(oVar2S18(0)='1' OR oVar2S19(0)='1' )then
          ADDM4K3S14(3)<='1';
          else
          ADDM4K3S14(3)<='0';
          end if;
        if(oVar2S22(0)='1' OR oVar2S23(0)='1' )then
          ADDM4K3S14(2)<='1';
          else
          ADDM4K3S14(2)<='0';
          end if;
        if(oVar2S12(0)='1' )then
          ADDM4K3S14(1)<='1';
          else
          ADDM4K3S14(1)<='0';
          end if;
        if(oVar2S16(0)='1' OR oVar2S17(0)='1' )then
          ADDM4K3S14(0)<='1';
          else
          ADDM4K3S14(0)<='0';
          end if;
        if(oVar2S14(0)='1' OR oVar2S15(0)='1' )then
          ADDM4K3S15(7)<='1';
          else
          ADDM4K3S15(7)<='0';
          end if;
        if(oVar2S24(0)='1' OR oVar2S25(0)='1' )then
          ADDM4K3S15(6)<='1';
          else
          ADDM4K3S15(6)<='0';
          end if;
        if(oVar2S6(0)='1' OR oVar2S7(0)='1' )then
          ADDM4K3S15(5)<='1';
          else
          ADDM4K3S15(5)<='0';
          end if;
        if(oVar2S8(0)='1' OR oVar2S9(0)='1' )then
          ADDM4K3S15(4)<='1';
          else
          ADDM4K3S15(4)<='0';
          end if;
        if(oVar2S10(0)='1' OR oVar2S11(0)='1' )then
          ADDM4K3S15(3)<='1';
          else
          ADDM4K3S15(3)<='0';
          end if;
        if(oVar2S4(0)='1' OR oVar2S5(0)='1' )then
          ADDM4K3S15(2)<='1';
          else
          ADDM4K3S15(2)<='0';
          end if;
        if(oVar2S2(0)='1' OR oVar2S3(0)='1' )then
          ADDM4K3S15(1)<='1';
          else
          ADDM4K3S15(1)<='0';
          end if;
        if(oVar2S0(0)='1' OR oVar2S1(0)='1' )then
          ADDM4K3S15(0)<='1';
          else
          ADDM4K3S15(0)<='0';
          end if;
        if(oVar2S208(0)='1' OR oVar2S209(0)='1' )then
          ADDM4K3S2(7)<='1';
          else
          ADDM4K3S2(7)<='0';
          end if;
        if(oVar2S154(0)='1' OR oVar2S155(0)='1' )then
          ADDM4K3S2(6)<='1';
          else
          ADDM4K3S2(6)<='0';
          end if;
        if(oVar2S202(0)='1' )then
          ADDM4K3S2(5)<='1';
          else
          ADDM4K3S2(5)<='0';
          end if;
        if(oVar2S214(0)='1' )then
          ADDM4K3S2(4)<='1';
          else
          ADDM4K3S2(4)<='0';
          end if;
        if(oVar2S157(0)='1' )then
          ADDM4K3S2(3)<='1';
          else
          ADDM4K3S2(3)<='0';
          end if;
        if(oVar2S146(0)='1' )then
          ADDM4K3S2(2)<='1';
          else
          ADDM4K3S2(2)<='0';
          end if;
        if(oVar2S210(0)='1' )then
          ADDM4K3S2(1)<='1';
          else
          ADDM4K3S2(1)<='0';
          end if;
        if(oVar2S212(0)='1' )then
          ADDM4K3S2(0)<='1';
          else
          ADDM4K3S2(0)<='0';
          end if;
        if(oVar2S144(0)='1' )then
          ADDM4K3S3(7)<='1';
          else
          ADDM4K3S3(7)<='0';
          end if;
        if(oVar2S245(0)='1' OR oVar2S246(0)='1' )then
          ADDM4K3S3(6)<='1';
          else
          ADDM4K3S3(6)<='0';
          end if;
        if(oVar2S204(0)='1' OR oVar2S205(0)='1' )then
          ADDM4K3S3(5)<='1';
          else
          ADDM4K3S3(5)<='0';
          end if;
        if(oVar1S433(0)='1' OR oVar1S434(0)='1' OR oVar1S435(0)='1' )then
          ADDM4K3S3(4)<='1';
          else
          ADDM4K3S3(4)<='0';
          end if;
        if(oVar2S196(0)='1' OR oVar2S197(0)='1' )then
          ADDM4K3S3(3)<='1';
          else
          ADDM4K3S3(3)<='0';
          end if;
        if(oVar2S206(0)='1' )then
          ADDM4K3S3(2)<='1';
          else
          ADDM4K3S3(2)<='0';
          end if;
        if(oVar2S194(0)='1' )then
          ADDM4K3S3(1)<='1';
          else
          ADDM4K3S3(1)<='0';
          end if;
        if(oVar2S138(0)='1' )then
          ADDM4K3S3(0)<='1';
          else
          ADDM4K3S3(0)<='0';
          end if;
        if(oVar2S142(0)='1' )then
          ADDM4K3S4(7)<='1';
          else
          ADDM4K3S4(7)<='0';
          end if;
        if(oVar2S247(0)='1' OR oVar2S248(0)='1' )then
          ADDM4K3S4(6)<='1';
          else
          ADDM4K3S4(6)<='0';
          end if;
        if(oVar2S148(0)='1' OR oVar2S149(0)='1' )then
          ADDM4K3S4(5)<='1';
          else
          ADDM4K3S4(5)<='0';
          end if;
        if(oVar2S198(0)='1' OR oVar2S199(0)='1' )then
          ADDM4K3S4(4)<='1';
          else
          ADDM4K3S4(4)<='0';
          end if;
        if(oVar2S182(0)='1' )then
          ADDM4K3S4(3)<='1';
          else
          ADDM4K3S4(3)<='0';
          end if;
        if(oVar2S152(0)='1' OR oVar2S153(0)='1' )then
          ADDM4K3S4(2)<='1';
          else
          ADDM4K3S4(2)<='0';
          end if;
        if(oVar2S140(0)='1' )then
          ADDM4K3S4(1)<='1';
          else
          ADDM4K3S4(1)<='0';
          end if;
        if(oVar2S200(0)='1' OR oVar2S201(0)='1' )then
          ADDM4K3S4(0)<='1';
          else
          ADDM4K3S4(0)<='0';
          end if;
        if(oVar2S188(0)='1' OR oVar2S189(0)='1' )then
          ADDM4K3S5(7)<='1';
          else
          ADDM4K3S5(7)<='0';
          end if;
        if(oVar2S134(0)='1' )then
          ADDM4K3S5(6)<='1';
          else
          ADDM4K3S5(6)<='0';
          end if;
        if(oVar2S92(0)='1' OR oVar2S93(0)='1' )then
          ADDM4K3S5(5)<='1';
          else
          ADDM4K3S5(5)<='0';
          end if;
        if(oVar2S180(0)='1' OR oVar2S181(0)='1' )then
          ADDM4K3S5(4)<='1';
          else
          ADDM4K3S5(4)<='0';
          end if;
        if(oVar2S124(0)='1' )then
          ADDM4K3S5(3)<='1';
          else
          ADDM4K3S5(3)<='0';
          end if;
        if(oVar2S126(0)='1' OR oVar2S127(0)='1' )then
          ADDM4K3S5(2)<='1';
          else
          ADDM4K3S5(2)<='0';
          end if;
        if(oVar2S132(0)='1' )then
          ADDM4K3S5(1)<='1';
          else
          ADDM4K3S5(1)<='0';
          end if;
        if(oVar2S249(0)='1' OR oVar2S250(0)='1' )then
          ADDM4K3S5(0)<='1';
          else
          ADDM4K3S5(0)<='0';
          end if;
        if(oVar2S186(0)='1' OR oVar2S187(0)='1' )then
          ADDM4K3S6(7)<='1';
          else
          ADDM4K3S6(7)<='0';
          end if;
        if(oVar2S176(0)='1' OR oVar2S177(0)='1' )then
          ADDM4K3S6(6)<='1';
          else
          ADDM4K3S6(6)<='0';
          end if;
        if(oVar2S164(0)='1' OR oVar2S165(0)='1' )then
          ADDM4K3S6(5)<='1';
          else
          ADDM4K3S6(5)<='0';
          end if;
        if(oVar2S172(0)='1' OR oVar2S173(0)='1' )then
          ADDM4K3S6(4)<='1';
          else
          ADDM4K3S6(4)<='0';
          end if;
        if(oVar2S174(0)='1' OR oVar2S175(0)='1' )then
          ADDM4K3S6(3)<='1';
          else
          ADDM4K3S6(3)<='0';
          end if;
        if(oVar2S166(0)='1' OR oVar2S167(0)='1' )then
          ADDM4K3S6(2)<='1';
          else
          ADDM4K3S6(2)<='0';
          end if;
        if(oVar2S150(0)='1' OR oVar2S151(0)='1' )then
          ADDM4K3S6(1)<='1';
          else
          ADDM4K3S6(1)<='0';
          end if;
        if(oVar2S159(0)='1' OR oVar2S160(0)='1' )then
          ADDM4K3S6(0)<='1';
          else
          ADDM4K3S6(0)<='0';
          end if;
        if(oVar2S178(0)='1' OR oVar2S179(0)='1' )then
          ADDM4K3S7(7)<='1';
          else
          ADDM4K3S7(7)<='0';
          end if;
        if(oVar2S192(0)='1' OR oVar2S193(0)='1' )then
          ADDM4K3S7(6)<='1';
          else
          ADDM4K3S7(6)<='0';
          end if;
        if(oVar2S184(0)='1' OR oVar2S185(0)='1' )then
          ADDM4K3S7(5)<='1';
          else
          ADDM4K3S7(5)<='0';
          end if;
        if(oVar2S136(0)='1' OR oVar2S137(0)='1' )then
          ADDM4K3S7(4)<='1';
          else
          ADDM4K3S7(4)<='0';
          end if;
        if(oVar2S112(0)='1' OR oVar2S113(0)='1' )then
          ADDM4K3S7(3)<='1';
          else
          ADDM4K3S7(3)<='0';
          end if;
        if(oVar2S190(0)='1' OR oVar2S191(0)='1' )then
          ADDM4K3S7(2)<='1';
          else
          ADDM4K3S7(2)<='0';
          end if;
        if(oVar2S130(0)='1' OR oVar2S131(0)='1' )then
          ADDM4K3S7(1)<='1';
          else
          ADDM4K3S7(1)<='0';
          end if;
        if(oVar2S80(0)='1' OR oVar2S81(0)='1' )then
          ADDM4K3S7(0)<='1';
          else
          ADDM4K3S7(0)<='0';
          end if;
        if(oVar1S649(0)='1' OR oVar1S650(0)='1' OR oVar1S651(0)='1' )then
          ADDM4K3S0(7)<='1';
          else
          ADDM4K3S0(7)<='0';
          end if;
        if(oVar2S235(0)='1' )then
          ADDM4K3S0(6)<='1';
          else
          ADDM4K3S0(6)<='0';
          end if;
        if(oVar2S233(0)='1' )then
          ADDM4K3S0(5)<='1';
          else
          ADDM4K3S0(5)<='0';
          end if;
        if(oVar2S241(0)='1' )then
          ADDM4K3S0(4)<='1';
          else
          ADDM4K3S0(4)<='0';
          end if;
        if(oVar1S652(0)='1' OR oVar1S653(0)='1' OR oVar1S654(0)='1' )then
          ADDM4K3S0(3)<='1';
          else
          ADDM4K3S0(3)<='0';
          end if;
        if(oVar2S225(0)='1' )then
          ADDM4K3S0(2)<='1';
          else
          ADDM4K3S0(2)<='0';
          end if;
        if(oVar2S231(0)='1' OR oVar2S232(0)='1' )then
          ADDM4K3S0(1)<='1';
          else
          ADDM4K3S0(1)<='0';
          end if;
        if(oVar2S223(0)='1' )then
          ADDM4K3S0(0)<='1';
          else
          ADDM4K3S0(0)<='0';
          end if;
        if(oVar2S229(0)='1' )then
          ADDM4K3S1(7)<='1';
          else
          ADDM4K3S1(7)<='0';
          end if;
        if(oVar2S227(0)='1' OR oVar2S228(0)='1' )then
          ADDM4K3S1(6)<='1';
          else
          ADDM4K3S1(6)<='0';
          end if;
        if(oVar2S239(0)='1' )then
          ADDM4K3S1(5)<='1';
          else
          ADDM4K3S1(5)<='0';
          end if;
        if(oVar1S608(0)='1' OR oVar1S609(0)='1' OR oVar1S610(0)='1' )then
          ADDM4K3S1(4)<='1';
          else
          ADDM4K3S1(4)<='0';
          end if;
        if(oVar2S219(0)='1' )then
          ADDM4K3S1(3)<='1';
          else
          ADDM4K3S1(3)<='0';
          end if;
        if(oVar2S243(0)='1' )then
          ADDM4K3S1(2)<='1';
          else
          ADDM4K3S1(2)<='0';
          end if;
        if(oVar2S216(0)='1' OR oVar2S217(0)='1' )then
          ADDM4K3S1(1)<='1';
          else
          ADDM4K3S1(1)<='0';
          end if;
        if(oVar2S221(0)='1' )then
          ADDM4K3S1(0)<='1';
          else
          ADDM4K3S1(0)<='0';
          end if;
 end if;
end process;
ADDM4K3S8c : ADDM4K3S8RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S8,
                q    => aVar3S8
    );
ADDM4K3S9c : ADDM4K3S9RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S9,
                q    => aVar3S9
    );
ADDM4K3S12c : ADDM4K3S12RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S12,
                q    => aVar3S12
    );
ADDM4K3S13c : ADDM4K3S13RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S13,
                q    => aVar3S13
    );
ADDM4K3S10c : ADDM4K3S10RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S10,
                q    => aVar3S10
    );
ADDM4K3S11c : ADDM4K3S11RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S11,
                q    => aVar3S11
    );
ADDM4K3S14c : ADDM4K3S14RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S14,
                q    => aVar3S14
    );
ADDM4K3S15c : ADDM4K3S15RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S15,
                q    => aVar3S15
    );
ADDM4K3S2c : ADDM4K3S2RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S2,
                q    => aVar3S2
    );
ADDM4K3S3c : ADDM4K3S3RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S3,
                q    => aVar3S3
    );
ADDM4K3S4c : ADDM4K3S4RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S4,
                q    => aVar3S4
    );
ADDM4K3S5c : ADDM4K3S5RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S5,
                q    => aVar3S5
    );
ADDM4K3S6c : ADDM4K3S6RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S6,
                q    => aVar3S6
    );
ADDM4K3S7c : ADDM4K3S7RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S7,
                q    => aVar3S7
    );
ADDM4K3S0c : ADDM4K3S0RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S0,
                q    => aVar3S0
    );
ADDM4K3S1c : ADDM4K3S1RAM PORT MAP (
                clock    => c1,
                address    => ADDM4K3S1,
                q    => aVar3S1
    );
Adder_1: Adder_type
port map(
dataa => aVar3S0, 
datab => aVar3S1, 
result => aVar4S0
);

Adder_2: Adder_type
port map(
dataa => aVar3S2, 
datab => aVar3S3, 
result => aVar4S1
);

Adder_3: Adder_type
port map(
dataa => aVar3S4, 
datab => aVar3S5, 
result => aVar4S2
);

Adder_4: Adder_type
port map(
dataa => aVar3S6, 
datab => aVar3S7, 
result => aVar4S3
);

Adder_5: Adder_type
port map(
dataa => aVar3S8, 
datab => aVar3S9, 
result => aVar4S4
);

Adder_6: Adder_type
port map(
dataa => aVar3S10, 
datab => aVar3S11, 
result => aVar4S5
);

Adder_7: Adder_type
port map(
dataa => aVar3S12, 
datab => aVar3S13, 
result => aVar4S6
);

Adder_8: Adder_type
port map(
dataa => aVar3S14, 
datab => aVar3S15, 
result => aVar4S7
);

Adder_9: Adder_type
port map(
dataa => aVar4S0, 
datab => aVar4S1, 
result => aVar5S0
);

Adder_10: Adder_type
port map(
dataa => aVar4S2, 
datab => aVar4S3, 
result => aVar5S1
);

Adder_11: Adder_type
port map(
dataa => aVar4S4, 
datab => aVar4S5, 
result => aVar5S2
);

Adder_12: Adder_type
port map(
dataa => aVar4S6, 
datab => aVar4S7, 
result => aVar5S3
);

Adder_13: Adder_type
port map(
dataa => aVar5S0, 
datab => aVar5S1, 
result => aVar6S0
);

Adder_14: Adder_type
port map(
dataa => aVar5S2, 
datab => aVar5S3, 
result => aVar6S1
);

Adder_15: Adder_type
port map(
dataa => aVar6S0, 
datab => aVar6S1, 
result => aVar7S0
);

end rtl;
